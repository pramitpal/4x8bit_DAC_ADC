* SPICE3 file created from dac_top.ext - technology: sky130A

.subckt dac_top VDDA VSSA VCCD VSSD VREFH Din0[0] Din0[1] Din0[2] Din0[3] Din0[4]
+ Din0[5] Din0[6] Din0[7] VOUT0 Din1[0] Din1[1] Din1[2] Din1[3] Din1[4] Din1[5] Din1[6]
+ Din1[7] VOUT1 Din2[0] Din2[1] Din2[2] Din2[3] Din2[4] Din2[5] Din2[6] Din2[7] VOUT2
+ Din3[0] Din3[1] Din3[2] Din3[3] Din3[4] Din3[5] Din3[6] Din3[7] VOUT3
X0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D5_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D5_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D5_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D5_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X8 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D1_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X10 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D1_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X11 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D1_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X12 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X13 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X14 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D1_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X15 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X16 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X17 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D0_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X18 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X19 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D0_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X20 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D0_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X21 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X22 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X23 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X24 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X25 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D0_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X26 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X27 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X28 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D0_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X29 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D0_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X30 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X31 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X32 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X33 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=506 ps=4.43k w=1 l=0.5
X34 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X35 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X36 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=250 ps=2.63k w=0.5 l=0.5
X37 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X38 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X39 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X40 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X41 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X42 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X43 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X44 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X45 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X46 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X47 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X48 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X49 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X50 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X51 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X52 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X53 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X54 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X55 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X56 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D2_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X57 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X58 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D2_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X59 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D2_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X60 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X61 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X62 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D2_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X63 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X64 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X65 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X66 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X67 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X68 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X69 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X70 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X71 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X72 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X73 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X74 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X75 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X76 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X77 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X78 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X79 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X80 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X81 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X82 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X83 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X84 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X85 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X86 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X87 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X88 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X89 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X90 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X91 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X92 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X93 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X94 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X95 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X96 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X97 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X98 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X99 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X100 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X101 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X102 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X103 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X104 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X105 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X106 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X107 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X108 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X109 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X110 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X111 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X112 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X113 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X114 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X115 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X116 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X117 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X118 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X119 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X120 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D3_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X121 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X122 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D3_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X123 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D3_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X124 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X125 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X126 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D3_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X127 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X128 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X129 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X130 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X131 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X132 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X133 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X134 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X135 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X136 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X137 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X138 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X139 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X140 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X141 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X142 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X143 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X144 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X145 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X146 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X147 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X148 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X149 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X150 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X151 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X152 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X153 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X154 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X155 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X156 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X157 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X158 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X159 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X160 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X161 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X162 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X163 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X164 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X165 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X166 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X167 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X168 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X169 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X170 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X171 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X172 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X173 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X174 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X175 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X176 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X177 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X178 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X179 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X180 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X181 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X182 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X183 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X184 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X185 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X186 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X187 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X188 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X189 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X190 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X191 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X192 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X193 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X194 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X195 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X196 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X197 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X198 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X199 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X200 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X201 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X202 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X203 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X204 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X205 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X206 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X207 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X208 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X209 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X210 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X211 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X212 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X213 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X214 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X215 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X216 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X217 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X218 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X219 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X220 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X221 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X222 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X223 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X224 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X225 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X226 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X227 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X228 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X229 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X230 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X231 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X232 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X233 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X234 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X235 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X236 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X237 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X238 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X239 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X240 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X241 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X242 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X243 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X244 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X245 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X246 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X247 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X248 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D4_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X249 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X250 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D4_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X251 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D4_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X252 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X253 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X254 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D4_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X255 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X256 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X257 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X258 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X259 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X260 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X261 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X262 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X263 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X264 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X265 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X266 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X267 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X268 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X269 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X270 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X271 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X272 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X273 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X274 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X275 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X276 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X277 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X278 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X279 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X280 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X281 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X282 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X283 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X284 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X285 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X286 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X287 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X288 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X289 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X290 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X291 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X292 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X293 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X294 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X295 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X296 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X297 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X298 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X299 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X300 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X301 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X302 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X303 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X304 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X305 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X306 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X307 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X308 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X309 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X310 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X311 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X312 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X313 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X314 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X315 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X316 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X317 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X318 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X319 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X320 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X321 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X322 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X323 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X324 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X325 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X326 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X327 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X328 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X329 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X330 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X331 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X332 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X333 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X334 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X335 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X336 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X337 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X338 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X339 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X340 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X341 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X342 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X343 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X344 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X345 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X346 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X347 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X348 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X349 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X350 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X351 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X352 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X353 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X354 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X355 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X356 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X357 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X358 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X359 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X360 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X361 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X362 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X363 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X364 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X365 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X366 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X367 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X368 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X369 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X370 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X371 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X372 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X373 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X374 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X375 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X376 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X377 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X378 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X379 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X380 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X381 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X382 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X383 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X384 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X385 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X386 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X387 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X388 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X389 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X390 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X391 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X392 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X393 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X394 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X395 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X396 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X397 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X398 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X399 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X400 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X401 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X402 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X403 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X404 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X405 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X406 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X407 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X408 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X409 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X410 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X411 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X412 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X413 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X414 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X415 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X416 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X417 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X418 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X419 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X420 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X421 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X422 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X423 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X424 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X425 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X426 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X427 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X428 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X429 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X430 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X431 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X432 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X433 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X434 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X435 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X436 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X437 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X438 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X439 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X440 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X441 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X442 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X443 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X444 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X445 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X446 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X447 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X448 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X449 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X450 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X451 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X452 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X453 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X454 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X455 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X456 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X457 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X458 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X459 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X460 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X461 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X462 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X463 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X464 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X465 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X466 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X467 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X468 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X469 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X470 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X471 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X472 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X473 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X474 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X475 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X476 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X477 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X478 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X479 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X480 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X481 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X482 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X483 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X484 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X485 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X486 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X487 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X488 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X489 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X490 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X491 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X492 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X493 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X494 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X495 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X496 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X497 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X498 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X499 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X500 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X501 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X502 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X503 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X504 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X505 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X506 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X507 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X508 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X509 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X510 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X511 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X512 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X513 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X514 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X515 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X516 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X517 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X518 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X519 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X520 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X521 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X522 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X523 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X524 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X525 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X526 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X527 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X528 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X529 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X530 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X531 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X532 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X533 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X534 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X535 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X536 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X537 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X538 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X539 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X540 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X541 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X542 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X543 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X544 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X545 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X546 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X547 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X548 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X549 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X550 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X551 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X552 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X553 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X554 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X555 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X556 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X557 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X558 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X559 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X560 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X561 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X562 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X563 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X564 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X565 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X566 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X567 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X568 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X569 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X570 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X571 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X572 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X573 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X574 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X575 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X576 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X577 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X578 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X579 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X580 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X581 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X582 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X583 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X584 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X585 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X586 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X587 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X588 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X589 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X590 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X591 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X592 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X593 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X594 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X595 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X596 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X597 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X598 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X599 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X600 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X601 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X602 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X603 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X604 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X605 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X606 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X607 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X608 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X609 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X610 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X611 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X612 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X613 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X614 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X615 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X616 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X617 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X618 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X619 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X620 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X621 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X622 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X623 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X624 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X625 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X626 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X627 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X628 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X629 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X630 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X631 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X632 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X633 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X634 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X635 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X636 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X637 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X638 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X639 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X640 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X641 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X642 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X643 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X644 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X645 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X646 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X647 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X648 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X649 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X650 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X651 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X652 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X653 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X654 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X655 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X656 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X657 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X658 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X659 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X660 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X661 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X662 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X663 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X664 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X665 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X666 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X667 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X668 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X669 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X670 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X671 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X672 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X673 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X674 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X675 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X676 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X677 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X678 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X679 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X680 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X681 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X682 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X683 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X684 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X685 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X686 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X687 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X688 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X689 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X690 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X691 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X692 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X693 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X694 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X695 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X696 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X697 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X698 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X699 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X700 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X701 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X702 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X703 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X704 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X705 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X706 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X707 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X708 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X709 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X710 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X711 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X712 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X713 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X714 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X715 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X716 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X717 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X718 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X719 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X720 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X721 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X722 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X723 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X724 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X725 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X726 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X727 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X728 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X729 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X730 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X731 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X732 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X733 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X734 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X735 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X736 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X737 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X738 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X739 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X740 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X741 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X742 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X743 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X744 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X745 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X746 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X747 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X748 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X749 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X750 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X751 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X752 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X753 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X754 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X755 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X756 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X757 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X758 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X759 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X760 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X761 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X762 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X763 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X764 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X765 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X766 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X767 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X768 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X769 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X770 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X771 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X772 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X773 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X774 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X775 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X776 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X777 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X778 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X779 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X780 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X781 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X782 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X783 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X784 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X785 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X786 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X787 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X788 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X789 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X790 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X791 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X792 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X793 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X794 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X795 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X796 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X797 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X798 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X799 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X800 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X801 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X802 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X803 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X804 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X805 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X806 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X807 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X808 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X809 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X810 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X811 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X812 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X813 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X814 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X815 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X816 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X817 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X818 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X819 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X820 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X821 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X822 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X823 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X824 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X825 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X826 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X827 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X828 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X829 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X830 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X831 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X832 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X833 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X834 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X835 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X836 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X837 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X838 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X839 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X840 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X841 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X842 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X843 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X844 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X845 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X846 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X847 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X848 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X849 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X850 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X851 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X852 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X853 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X854 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X855 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X856 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X857 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X858 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X859 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X860 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X861 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X862 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X863 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X864 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X865 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X866 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X867 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X868 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X869 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X870 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X871 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X872 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X873 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X874 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X875 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X876 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X877 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X878 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X879 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X880 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X881 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X882 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X883 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X884 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X885 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X886 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X887 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X888 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X889 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X890 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X891 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X892 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X893 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X894 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X895 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X896 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X897 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X898 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X899 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X900 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X901 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X902 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X903 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X904 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X905 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X906 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X907 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X908 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X909 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X910 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X911 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X912 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X913 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X914 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X915 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X916 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X917 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X918 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X919 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X920 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X921 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X922 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X923 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X924 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X925 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X926 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X927 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X928 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X929 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X930 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X931 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X932 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X933 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X934 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X935 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X936 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X937 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X938 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X939 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X940 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X941 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X942 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X943 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X944 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X945 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X946 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X947 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X948 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X949 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X950 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X951 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X952 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X953 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X954 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X955 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X956 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X957 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X958 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X959 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X960 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X961 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X962 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X963 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X964 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X965 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X966 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X967 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X968 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X969 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X970 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X971 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X972 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X973 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X974 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X975 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X976 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X977 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X978 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X979 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X980 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X981 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X982 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X983 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X984 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X985 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X986 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X987 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X988 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X989 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X990 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X991 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X992 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X993 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X994 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X995 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X996 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X997 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X998 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X999 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1000 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1001 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1002 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1003 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1004 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1005 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1006 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1007 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1008 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D6_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1009 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/D6 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1010 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D6_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1011 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D6_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1012 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/D6 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1013 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1014 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D6_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1015 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1016 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1017 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1018 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1019 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1020 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1021 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1022 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1023 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1024 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1025 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1026 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1027 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1028 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1029 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1030 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1031 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1032 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1033 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1034 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1035 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1036 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1037 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1038 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1039 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1040 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1041 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1042 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1043 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1044 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1045 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1046 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1047 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1048 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1049 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1050 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1051 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1052 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1053 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1054 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1055 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1056 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1057 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1058 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1059 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1060 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1061 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1062 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1063 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1064 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1065 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1066 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1067 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1068 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1069 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1070 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1071 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1072 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1073 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1074 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1075 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1076 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1077 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1078 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1079 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1080 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1081 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1082 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1083 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1084 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1085 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1086 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1087 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1088 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1089 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1090 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1091 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1092 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1093 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1094 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1095 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1096 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1097 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1098 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1099 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1100 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1101 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1102 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1103 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1104 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1105 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1106 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1107 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1108 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1109 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1110 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1111 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1112 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1113 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1114 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1115 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1116 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1117 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1118 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1119 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1120 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1121 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1122 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1123 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1124 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1125 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1126 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1127 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1128 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1129 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1130 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1131 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1132 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1133 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1134 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1135 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1136 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1137 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1138 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1139 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1140 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1141 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1142 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1143 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1144 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1145 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1146 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1147 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1148 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1149 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1150 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1151 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1152 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1153 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1154 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1155 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1156 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1157 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1158 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1159 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1160 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1161 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1162 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1163 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1164 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1165 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1166 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1167 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1168 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1169 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1170 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1171 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1172 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1173 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1174 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1175 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1176 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1177 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1178 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1179 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1180 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1181 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1182 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1183 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1184 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1185 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1186 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1187 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1188 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1189 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1190 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1191 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1192 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1193 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1194 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1195 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1196 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1197 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1198 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1199 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1200 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1201 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1202 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1203 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1204 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1205 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1206 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1207 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1208 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1209 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1210 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1211 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1212 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1213 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1214 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1215 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1216 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1217 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1218 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1219 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1220 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1221 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1222 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1223 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1224 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1225 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1226 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1227 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1228 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1229 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1230 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1231 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1232 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1233 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1234 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1235 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1236 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1237 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1238 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1239 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1240 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1241 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1242 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1243 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1244 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1245 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1246 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1247 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1248 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1249 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1250 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1251 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1252 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1253 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1254 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1255 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1256 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1257 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1258 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1259 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1260 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1261 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1262 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1263 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1264 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1265 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1266 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1267 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1268 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1269 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1270 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1271 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1272 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1273 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1274 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1275 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1276 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1277 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1278 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1279 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1280 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1281 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1282 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1283 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1284 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1285 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1286 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1287 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1288 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1289 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1290 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1291 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1292 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1293 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1294 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1295 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1296 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1297 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1298 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1299 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1300 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1301 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1302 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1303 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1304 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1305 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1306 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1307 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1308 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1309 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1310 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1311 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1312 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1313 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1314 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1315 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1316 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1317 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1318 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1319 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1320 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1321 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1322 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1323 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1324 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1325 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1326 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1327 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1328 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1329 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1330 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1331 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1332 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1333 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1334 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1335 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1336 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1337 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1338 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1339 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1340 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1341 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1342 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1343 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1344 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1345 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1346 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1347 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1348 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1349 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1350 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1351 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1352 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1353 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1354 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1355 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1356 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1357 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1358 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1359 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1360 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1361 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1362 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1363 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1364 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1365 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1366 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1367 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1368 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1369 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1370 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1371 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1372 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1373 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1374 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1375 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1376 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1377 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1378 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1379 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1380 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1381 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1382 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1383 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1384 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1385 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1386 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1387 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1388 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1389 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1390 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1391 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1392 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1393 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1394 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1395 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1396 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1397 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1398 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1399 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1400 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1401 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1402 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1403 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1404 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1405 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1406 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1407 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1408 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1409 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1410 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1411 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1412 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1413 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1414 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1415 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1416 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1417 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1418 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1419 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1420 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1421 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1422 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1423 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1424 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1425 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1426 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1427 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1428 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1429 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1430 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1431 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1432 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1433 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1434 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1435 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1436 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1437 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1438 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1439 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1440 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1441 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1442 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1443 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1444 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1445 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1446 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1447 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1448 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1449 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1450 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1451 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1452 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1453 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1454 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1455 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1456 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1457 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1458 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1459 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1460 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1461 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1462 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1463 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1464 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1465 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1466 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1467 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1468 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1469 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1470 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1471 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1472 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1473 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1474 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1475 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1476 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1477 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1478 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1479 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1480 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1481 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1482 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1483 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1484 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1485 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1486 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1487 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1488 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1489 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1490 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1491 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1492 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1493 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1494 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1495 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1496 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1497 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1498 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1499 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1500 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1501 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1502 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1503 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1504 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1505 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1506 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1507 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1508 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1509 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1510 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1511 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1512 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1513 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1514 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1515 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1516 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1517 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1518 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1519 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1520 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1521 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1522 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1523 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1524 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1525 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1526 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1527 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1528 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1529 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1530 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1531 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1532 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1533 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1534 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1535 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1536 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1537 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1538 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1539 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1540 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1541 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1542 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1543 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1544 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1545 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1546 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1547 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1548 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1549 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1550 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1551 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1552 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1553 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1554 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1555 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1556 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1557 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1558 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1559 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1560 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1561 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1562 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1563 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1564 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1565 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1566 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1567 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1568 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1569 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1570 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1571 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1572 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1573 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1574 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1575 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1576 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1577 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1578 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1579 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1580 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1581 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1582 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1583 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1584 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1585 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1586 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1587 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1588 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1589 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1590 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1591 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1592 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1593 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1594 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1595 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1596 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1597 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1598 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1599 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1600 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1601 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1602 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1603 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1604 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1605 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1606 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1607 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1608 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1609 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1610 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1611 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1612 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1613 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1614 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1615 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1616 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1617 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1618 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1619 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1620 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1621 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1622 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1623 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1624 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1625 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1626 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1627 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1628 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1629 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1630 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1631 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1632 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1633 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1634 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1635 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1636 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1637 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1638 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1639 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1640 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1641 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1642 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1643 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1644 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1645 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1646 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1647 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1648 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1649 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1650 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1651 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1652 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1653 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1654 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1655 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1656 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1657 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1658 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1659 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1660 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1661 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1662 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1663 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1664 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1665 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1666 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1667 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1668 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1669 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1670 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1671 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1672 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1673 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1674 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1675 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1676 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1677 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1678 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1679 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1680 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1681 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1682 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1683 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1684 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1685 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1686 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1687 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1688 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1689 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1690 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1691 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1692 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1693 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1694 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1695 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1696 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1697 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1698 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1699 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1700 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1701 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1702 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1703 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1704 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1705 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1706 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1707 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1708 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1709 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1710 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1711 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1712 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1713 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1714 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1715 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1716 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1717 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1718 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1719 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1720 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1721 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1722 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1723 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1724 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1725 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1726 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1727 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1728 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1729 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1730 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1731 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1732 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1733 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1734 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1735 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1736 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1737 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1738 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1739 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1740 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1741 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1742 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1743 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1744 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1745 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1746 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1747 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1748 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1749 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1750 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1751 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1752 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1753 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1754 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1755 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1756 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1757 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1758 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1759 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1760 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1761 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1762 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1763 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1764 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1765 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1766 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1767 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1768 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1769 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1770 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1771 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1772 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1773 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1774 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1775 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1776 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1777 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1778 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1779 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1780 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1781 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1782 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1783 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1784 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1785 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1786 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1787 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1788 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1789 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1790 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1791 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1792 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1793 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1794 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1795 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1796 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1797 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1798 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1799 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1800 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1801 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1802 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1803 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1804 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1805 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1806 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1807 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1808 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1809 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1810 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1811 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1812 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1813 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1814 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1815 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1816 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1817 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1818 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1819 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1820 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1821 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1822 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1823 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1824 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1825 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1826 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1827 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1828 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1829 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1830 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1831 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1832 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1833 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1834 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1835 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1836 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1837 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1838 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1839 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1840 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1841 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1842 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1843 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1844 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1845 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1846 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1847 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1848 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1849 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1850 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1851 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1852 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1853 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1854 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1855 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1856 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1857 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1858 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1859 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1860 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1861 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1862 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1863 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1864 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1865 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1866 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1867 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1868 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1869 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1870 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1871 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1872 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1873 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1874 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1875 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1876 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1877 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1878 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1879 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1880 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1881 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1882 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1883 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1884 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1885 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1886 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1887 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1888 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1889 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1890 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1891 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1892 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1893 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1894 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1895 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1896 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1897 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1898 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1899 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1900 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1901 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1902 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1903 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1904 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1905 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1906 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1907 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1908 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1909 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1910 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1911 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1912 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1913 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1914 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1915 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1916 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1917 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1918 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1919 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1920 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1921 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1922 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1923 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1924 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1925 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1926 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1927 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1928 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1929 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1930 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1931 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1932 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1933 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1934 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1935 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1936 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1937 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1938 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1939 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1940 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1941 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1942 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1943 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1944 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1945 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1946 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1947 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1948 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1949 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1950 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1951 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1952 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1953 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1954 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1955 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1956 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1957 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1958 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1959 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1960 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1961 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1962 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1963 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1964 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1965 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1966 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1967 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1968 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1969 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1970 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1971 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1972 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1973 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1974 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1975 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1976 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1977 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1978 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1979 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1980 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1981 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1982 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1983 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1984 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1985 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1986 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1987 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1988 VSSA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=95.1 pd=148 as=0 ps=0 w=1 l=0.5
X1989 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1990 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1991 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1992 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1993 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1994 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1995 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1996 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1997 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1998 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1999 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2000 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2001 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2002 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2003 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2004 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2005 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2006 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2007 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2008 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2009 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2010 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2011 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2012 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2013 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2014 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2015 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2016 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2017 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2018 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2019 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2020 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2021 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2022 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2023 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2024 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/D6 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2025 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D6 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2026 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/D6 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2027 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/D6 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2028 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D6 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2029 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2030 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/D6 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2031 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2032 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D7_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=3.16 as=0 ps=0 w=0.5 l=0.5
X2033 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D7 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2034 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D7_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2035 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D7_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.5
X2036 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D7 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2037 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2038 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D7_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2039 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/7_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2040 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1423_1248# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2041 VSSD Din0[0] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.2
X2042 VSSD Din0[0] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X2043 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2044 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1353_675# Din0[0] VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.2
X2045 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X2046 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1423_1248# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2047 VSSD Din0[1] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=3.9 pd=45.4 as=0.122 ps=1.42 w=0.42 l=0.2
X2048 VSSD Din0[1] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=9.28 pd=82.6 as=0.29 ps=2.58 w=1 l=0.5
X2049 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2050 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1353_675# Din0[1] VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=4.64 ps=50.6 w=0.5 l=0.2
X2051 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2052 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1423_1248# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2053 VSSD Din0[2] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X2054 VSSD Din0[2] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2055 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2056 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1353_675# Din0[2] VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X2057 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2058 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1423_1248# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2059 VSSD Din0[3] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X2060 VSSD Din0[3] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2061 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2062 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1353_675# Din0[3] VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X2063 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2064 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1423_1248# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2065 VSSD Din0[4] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X2066 VSSD Din0[4] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2067 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2068 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1353_675# Din0[4] VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X2069 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2070 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1423_1248# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2071 VSSD Din0[5] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X2072 VSSD Din0[5] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2073 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2074 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1353_675# Din0[5] VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X2075 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2076 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1423_1248# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D6 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2077 VSSD Din0[6] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X2078 VSSD Din0[6] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2079 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D6 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2080 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1353_675# Din0[6] VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X2081 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D6 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2082 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1423_1248# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D7 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2083 VSSD Din0[7] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X2084 VSSD Din0[7] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2085 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D7 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2086 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1353_675# Din0[7] VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X2087 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/8_bit_dac_0/D7 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2088 VSSA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_3246_n774# VOUT0 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=1
X2089 VOUT0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_3246_n774# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X2090 VDDA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_1618_n334# VOUT0 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X2091 VDDA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_394_n920# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_1704_376# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X2092 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_1704_376# VOUT0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_1446_376# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=1
X2093 VDDA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_1618_n334# VOUT0 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.6 as=1.16 ps=8.29 w=8 l=1
X2094 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_408_552# VSSA VSSA sky130_fd_pr__res_generic_nd__hv w=0.48 l=4.46
X2095 VSSA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_1022_n914# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_2158_n774# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X2096 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_2158_n774# VOUT0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_1900_n774# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X2097 VSSA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_2894_292# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_2894_292# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X2098 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_1022_n914# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_394_n920# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.6 as=1.16 ps=8.29 w=8 l=1
X2099 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_1776_n834# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_408_552# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_1618_n334# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X2100 VSSA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_1022_n914# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_1446_376# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X2101 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_2894_292# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_408_552# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_1900_n774# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X2102 VDDA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_408_552# VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=8.32
X2103 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_2416_n774# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_394_n920# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=1
X2104 VDDA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_394_n920# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_394_n920# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.29 as=2.32 ps=16.6 w=8 l=1
X2105 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_1446_376# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_408_552# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_1300_n354# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X2106 VOUT0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_3246_n774# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=1
X2107 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_2416_n774# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_2158_n774# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X2108 VOUT0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_1618_n334# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.29 as=2.32 ps=16.6 w=8 l=1
X2109 VOUT0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_1618_n334# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X2110 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_1776_n834# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_1704_376# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=1
X2111 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_1618_n334# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_1300_n354# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.6 as=1.16 ps=8.29 w=8 l=1
X2112 VSSA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_3246_n774# VOUT0 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X2113 VSSA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_1022_n914# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_1022_n914# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
X2114 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_1776_n834# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_1022_n914# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X2115 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_3246_n774# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_2894_292# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X2116 VSSA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_394_n920# VSSA sky130_fd_pr__res_generic_nd__hv w=0.41 l=15.7
X2117 VDDA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_394_n920# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_1900_n774# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=1
X2118 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_3246_n774# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_408_552# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_2416_n774# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X2119 VDDA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_1300_n354# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[0]/opamp_0/a_1300_n354# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.29 as=2.32 ps=16.6 w=8 l=1
X2120 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D5_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2121 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2122 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D5_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2123 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D5_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2124 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2125 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2126 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D5_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2127 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2128 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D1_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2129 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2130 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D1_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2131 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D1_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2132 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2133 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2134 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D1_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2135 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2136 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2137 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D0_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2138 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2139 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D0_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2140 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D0_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2141 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2142 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2143 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2144 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2145 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D0_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2146 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2147 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2148 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D0_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2149 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D0_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2150 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2151 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2152 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2153 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2154 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2155 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2156 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2157 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2158 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2159 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2160 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2161 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2162 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2163 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2164 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2165 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2166 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2167 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2168 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2169 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2170 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2171 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2172 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2173 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2174 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2175 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2176 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D2_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2177 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2178 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D2_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2179 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D2_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2180 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2181 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2182 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D2_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2183 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2184 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2185 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2186 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2187 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2188 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2189 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2190 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2191 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2192 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2193 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2194 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2195 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2196 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2197 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2198 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2199 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2200 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2201 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2202 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2203 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2204 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2205 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2206 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2207 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2208 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2209 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2210 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2211 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2212 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2213 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2214 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2215 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2216 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2217 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2218 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2219 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2220 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2221 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2222 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2223 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2224 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2225 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2226 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2227 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2228 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2229 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2230 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2231 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2232 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2233 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2234 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2235 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2236 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2237 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2238 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2239 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2240 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D3_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2241 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2242 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D3_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2243 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D3_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2244 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2245 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2246 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D3_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2247 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2248 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2249 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2250 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2251 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2252 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2253 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2254 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2255 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2256 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2257 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2258 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2259 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2260 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2261 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2262 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2263 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2264 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2265 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2266 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2267 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2268 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2269 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2270 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2271 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2272 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2273 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2274 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2275 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2276 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2277 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2278 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2279 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2280 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2281 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2282 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2283 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2284 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2285 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2286 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2287 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2288 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2289 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2290 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2291 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2292 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2293 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2294 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2295 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2296 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2297 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2298 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2299 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2300 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2301 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2302 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2303 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2304 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2305 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2306 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2307 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2308 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2309 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2310 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2311 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2312 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2313 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2314 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2315 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2316 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2317 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2318 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2319 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2320 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2321 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2322 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2323 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2324 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2325 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2326 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2327 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2328 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2329 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2330 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2331 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2332 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2333 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2334 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2335 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2336 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2337 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2338 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2339 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2340 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2341 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2342 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2343 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2344 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2345 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2346 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2347 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2348 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2349 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2350 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2351 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2352 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2353 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2354 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2355 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2356 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2357 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2358 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2359 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2360 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2361 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2362 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2363 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2364 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2365 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2366 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2367 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2368 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D4_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2369 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2370 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D4_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2371 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D4_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2372 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2373 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2374 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D4_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2375 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2376 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2377 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2378 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2379 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2380 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2381 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2382 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2383 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2384 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2385 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2386 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2387 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2388 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2389 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2390 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2391 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2392 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2393 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2394 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2395 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2396 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2397 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2398 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2399 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2400 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2401 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2402 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2403 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2404 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2405 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2406 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2407 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2408 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2409 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2410 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2411 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2412 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2413 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2414 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2415 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2416 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2417 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2418 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2419 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2420 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2421 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2422 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2423 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2424 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2425 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2426 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2427 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2428 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2429 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2430 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2431 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2432 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2433 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2434 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2435 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2436 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2437 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2438 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2439 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2440 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2441 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2442 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2443 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2444 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2445 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2446 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2447 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2448 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2449 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2450 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2451 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2452 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2453 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2454 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2455 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2456 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2457 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2458 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2459 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2460 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2461 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2462 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2463 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2464 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2465 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2466 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2467 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2468 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2469 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2470 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2471 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2472 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2473 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2474 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2475 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2476 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2477 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2478 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2479 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2480 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2481 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2482 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2483 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2484 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2485 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2486 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2487 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2488 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2489 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2490 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2491 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2492 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2493 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2494 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2495 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2496 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2497 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2498 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2499 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2500 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2501 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2502 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2503 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2504 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2505 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2506 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2507 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2508 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2509 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2510 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2511 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2512 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2513 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2514 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2515 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2516 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2517 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2518 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2519 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2520 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2521 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2522 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2523 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2524 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2525 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2526 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2527 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2528 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2529 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2530 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2531 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2532 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2533 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2534 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2535 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2536 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2537 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2538 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2539 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2540 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2541 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2542 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2543 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2544 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2545 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2546 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2547 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2548 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2549 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2550 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2551 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2552 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2553 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2554 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2555 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2556 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2557 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2558 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2559 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2560 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2561 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2562 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2563 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2564 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2565 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2566 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2567 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2568 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2569 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2570 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2571 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2572 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2573 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2574 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2575 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2576 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2577 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2578 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2579 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2580 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2581 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2582 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2583 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2584 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2585 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2586 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2587 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2588 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2589 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2590 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2591 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2592 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2593 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2594 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2595 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2596 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2597 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2598 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2599 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2600 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2601 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2602 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2603 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2604 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2605 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2606 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2607 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2608 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2609 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2610 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2611 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2612 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2613 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2614 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2615 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2616 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2617 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2618 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2619 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2620 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2621 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2622 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2623 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2624 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2625 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2626 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2627 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2628 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2629 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2630 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2631 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2632 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2633 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2634 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2635 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2636 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2637 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2638 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2639 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2640 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2641 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2642 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2643 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2644 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2645 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2646 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2647 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2648 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2649 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2650 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2651 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2652 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2653 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2654 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2655 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2656 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2657 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2658 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2659 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2660 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2661 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2662 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2663 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2664 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2665 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2666 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2667 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2668 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2669 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2670 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2671 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2672 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2673 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2674 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2675 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2676 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2677 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2678 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2679 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2680 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2681 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2682 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2683 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2684 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2685 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2686 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2687 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2688 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2689 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2690 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2691 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2692 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2693 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2694 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2695 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2696 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2697 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2698 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2699 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2700 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2701 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2702 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2703 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2704 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2705 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2706 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2707 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2708 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2709 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2710 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2711 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2712 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2713 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2714 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2715 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2716 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2717 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2718 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2719 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2720 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2721 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2722 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2723 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2724 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2725 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2726 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2727 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2728 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2729 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2730 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2731 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2732 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2733 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2734 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2735 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2736 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2737 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2738 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2739 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2740 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2741 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2742 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2743 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2744 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2745 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2746 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2747 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2748 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2749 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2750 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2751 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2752 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2753 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2754 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2755 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2756 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2757 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2758 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2759 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2760 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2761 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2762 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2763 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2764 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2765 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2766 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2767 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2768 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2769 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2770 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2771 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2772 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2773 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2774 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2775 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2776 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2777 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2778 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2779 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2780 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2781 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2782 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2783 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2784 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2785 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2786 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2787 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2788 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2789 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2790 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2791 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2792 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2793 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2794 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2795 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2796 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2797 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2798 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2799 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2800 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2801 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2802 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2803 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2804 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2805 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2806 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2807 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2808 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2809 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2810 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2811 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2812 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2813 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2814 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2815 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2816 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2817 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2818 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2819 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2820 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2821 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2822 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2823 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2824 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2825 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2826 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2827 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2828 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2829 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2830 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2831 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2832 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2833 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2834 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2835 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2836 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2837 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2838 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2839 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2840 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2841 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2842 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2843 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2844 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2845 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2846 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2847 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2848 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2849 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2850 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2851 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2852 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2853 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2854 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2855 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2856 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2857 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2858 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2859 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2860 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2861 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2862 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2863 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2864 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2865 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2866 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2867 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2868 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2869 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2870 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2871 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2872 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2873 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2874 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2875 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2876 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2877 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2878 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2879 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2880 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2881 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2882 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2883 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2884 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2885 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2886 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2887 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2888 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2889 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2890 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2891 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2892 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2893 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2894 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2895 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2896 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2897 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2898 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2899 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2900 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2901 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2902 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2903 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2904 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2905 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2906 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2907 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2908 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2909 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2910 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2911 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2912 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2913 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2914 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2915 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2916 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2917 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2918 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2919 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2920 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2921 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2922 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2923 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2924 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2925 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2926 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2927 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2928 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2929 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2930 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2931 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2932 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2933 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2934 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2935 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2936 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2937 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2938 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2939 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2940 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2941 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2942 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2943 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2944 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2945 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2946 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2947 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2948 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2949 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2950 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2951 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2952 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2953 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2954 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2955 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2956 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2957 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2958 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2959 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2960 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X2961 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2962 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2963 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X2964 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2965 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2966 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2967 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2968 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2969 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2970 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2971 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2972 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2973 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2974 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2975 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2976 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X2977 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2978 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2979 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2980 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X2981 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2982 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2983 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2984 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2985 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2986 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2987 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2988 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2989 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2990 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2991 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2992 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2993 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2994 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2995 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2996 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2997 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2998 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2999 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3000 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3001 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3002 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3003 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3004 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3005 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3006 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3007 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3008 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3009 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3010 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3011 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3012 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3013 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3014 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3015 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3016 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3017 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3018 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3019 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3020 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3021 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3022 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3023 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3024 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3025 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3026 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3027 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3028 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3029 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3030 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3031 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3032 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3033 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3034 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3035 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3036 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3037 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3038 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3039 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3040 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3041 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3042 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3043 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3044 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3045 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3046 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3047 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3048 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3049 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3050 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3051 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3052 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3053 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3054 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3055 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3056 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3057 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3058 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3059 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3060 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3061 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3062 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3063 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3064 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3065 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3066 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3067 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3068 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3069 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3070 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3071 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3072 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3073 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3074 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3075 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3076 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3077 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3078 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3079 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3080 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3081 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3082 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3083 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3084 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3085 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3086 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3087 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3088 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3089 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3090 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3091 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3092 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3093 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3094 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3095 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3096 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3097 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3098 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3099 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3100 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3101 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3102 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3103 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3104 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3105 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3106 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3107 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3108 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3109 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3110 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3111 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3112 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3113 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3114 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3115 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3116 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3117 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3118 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3119 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3120 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3121 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3122 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3123 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3124 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3125 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3126 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3127 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3128 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D6_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3129 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/D6 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3130 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D6_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3131 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D6_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3132 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/D6 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3133 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3134 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D6_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3135 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3136 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3137 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3138 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3139 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3140 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3141 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3142 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3143 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3144 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3145 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3146 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3147 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3148 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3149 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3150 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3151 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3152 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3153 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3154 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3155 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3156 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3157 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3158 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3159 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3160 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3161 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3162 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3163 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3164 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3165 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3166 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3167 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3168 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3169 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3170 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3171 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3172 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3173 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3174 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3175 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3176 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3177 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3178 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3179 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3180 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3181 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3182 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3183 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3184 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3185 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3186 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3187 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3188 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3189 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3190 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3191 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3192 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3193 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3194 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3195 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3196 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3197 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3198 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3199 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3200 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3201 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3202 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3203 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3204 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3205 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3206 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3207 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3208 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3209 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3210 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3211 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3212 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3213 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3214 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3215 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3216 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3217 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3218 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3219 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3220 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3221 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3222 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3223 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3224 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3225 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3226 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3227 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3228 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3229 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3230 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3231 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3232 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3233 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3234 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3235 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3236 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3237 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3238 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3239 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3240 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3241 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3242 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3243 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3244 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3245 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3246 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3247 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3248 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3249 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3250 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3251 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3252 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3253 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3254 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3255 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3256 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3257 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3258 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3259 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3260 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3261 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3262 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3263 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3264 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3265 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3266 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3267 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3268 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3269 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3270 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3271 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3272 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3273 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3274 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3275 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3276 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3277 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3278 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3279 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3280 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3281 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3282 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3283 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3284 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3285 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3286 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3287 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3288 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3289 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3290 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3291 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3292 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3293 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3294 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3295 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3296 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3297 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3298 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3299 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3300 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3301 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3302 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3303 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3304 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3305 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3306 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3307 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3308 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3309 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3310 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3311 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3312 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3313 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3314 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3315 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3316 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3317 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3318 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3319 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3320 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3321 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3322 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3323 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3324 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3325 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3326 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3327 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3328 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3329 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3330 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3331 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3332 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3333 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3334 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3335 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3336 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3337 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3338 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3339 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3340 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3341 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3342 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3343 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3344 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3345 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3346 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3347 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3348 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3349 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3350 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3351 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3352 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3353 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3354 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3355 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3356 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3357 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3358 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3359 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3360 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3361 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3362 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3363 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3364 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3365 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3366 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3367 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3368 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3369 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3370 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3371 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3372 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3373 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3374 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3375 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3376 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3377 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3378 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3379 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3380 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3381 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3382 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3383 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3384 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3385 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3386 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3387 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3388 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3389 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3390 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3391 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3392 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3393 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3394 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3395 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3396 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3397 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3398 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3399 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3400 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3401 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3402 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3403 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3404 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3405 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3406 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3407 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3408 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3409 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3410 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3411 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3412 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3413 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3414 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3415 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3416 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3417 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3418 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3419 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3420 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3421 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3422 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3423 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3424 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3425 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3426 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3427 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3428 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3429 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3430 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3431 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3432 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3433 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3434 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3435 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3436 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3437 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3438 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3439 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3440 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3441 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3442 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3443 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3444 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3445 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3446 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3447 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3448 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3449 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3450 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3451 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3452 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3453 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3454 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3455 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3456 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3457 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3458 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3459 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3460 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3461 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3462 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3463 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3464 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3465 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3466 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3467 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3468 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3469 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3470 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3471 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3472 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3473 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3474 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3475 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3476 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3477 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3478 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3479 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3480 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3481 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3482 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3483 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3484 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3485 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3486 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3487 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3488 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3489 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3490 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3491 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3492 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3493 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3494 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3495 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3496 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3497 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3498 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3499 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3500 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3501 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3502 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3503 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3504 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3505 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3506 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3507 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3508 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3509 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3510 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3511 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3512 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3513 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3514 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3515 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3516 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3517 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3518 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3519 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3520 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3521 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3522 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3523 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3524 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3525 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3526 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3527 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3528 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3529 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3530 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3531 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3532 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3533 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3534 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3535 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3536 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3537 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3538 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3539 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3540 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3541 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3542 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3543 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3544 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3545 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3546 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3547 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3548 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3549 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3550 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3551 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3552 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3553 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3554 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3555 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3556 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3557 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3558 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3559 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3560 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3561 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3562 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3563 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3564 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3565 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3566 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3567 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3568 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3569 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3570 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3571 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3572 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3573 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3574 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3575 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3576 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3577 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3578 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3579 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3580 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3581 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3582 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3583 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3584 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3585 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3586 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3587 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3588 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3589 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3590 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3591 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3592 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3593 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3594 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3595 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3596 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3597 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3598 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3599 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3600 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3601 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3602 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3603 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3604 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3605 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3606 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3607 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3608 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3609 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3610 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3611 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3612 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3613 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3614 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3615 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3616 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3617 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3618 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3619 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3620 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3621 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3622 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3623 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3624 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3625 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3626 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3627 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3628 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3629 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3630 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3631 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3632 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3633 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3634 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3635 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3636 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3637 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3638 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3639 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3640 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3641 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3642 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3643 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3644 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3645 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3646 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3647 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3648 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3649 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3650 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3651 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3652 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3653 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3654 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3655 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3656 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3657 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3658 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3659 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3660 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3661 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3662 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3663 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3664 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3665 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3666 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3667 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3668 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3669 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3670 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3671 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3672 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3673 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3674 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3675 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3676 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3677 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3678 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3679 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3680 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3681 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3682 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3683 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3684 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3685 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3686 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3687 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3688 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3689 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3690 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3691 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3692 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3693 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3694 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3695 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3696 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3697 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3698 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3699 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3700 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3701 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3702 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3703 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3704 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3705 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3706 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3707 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3708 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3709 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3710 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3711 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3712 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3713 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3714 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3715 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3716 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3717 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3718 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3719 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3720 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3721 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3722 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3723 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3724 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3725 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3726 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3727 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3728 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3729 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3730 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3731 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3732 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3733 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3734 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3735 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3736 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3737 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3738 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3739 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3740 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3741 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3742 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3743 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3744 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3745 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3746 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3747 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3748 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3749 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3750 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3751 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3752 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3753 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3754 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3755 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3756 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3757 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3758 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3759 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3760 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3761 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3762 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3763 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3764 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3765 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3766 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3767 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3768 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3769 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3770 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3771 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3772 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3773 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3774 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3775 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3776 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3777 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3778 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3779 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3780 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3781 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3782 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3783 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3784 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3785 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3786 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3787 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3788 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3789 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3790 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3791 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3792 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3793 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3794 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3795 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3796 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3797 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3798 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3799 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3800 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3801 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3802 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3803 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3804 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3805 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3806 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3807 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3808 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3809 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3810 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3811 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3812 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3813 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3814 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3815 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3816 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3817 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3818 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3819 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3820 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3821 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3822 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3823 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3824 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3825 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3826 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3827 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3828 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3829 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3830 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3831 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3832 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3833 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3834 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3835 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3836 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3837 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3838 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3839 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3840 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3841 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3842 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3843 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3844 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3845 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3846 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3847 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3848 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3849 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3850 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3851 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3852 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3853 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3854 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3855 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3856 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3857 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3858 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3859 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3860 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3861 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3862 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3863 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3864 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3865 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3866 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3867 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3868 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3869 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3870 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3871 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3872 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3873 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3874 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3875 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3876 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3877 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3878 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3879 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3880 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3881 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3882 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3883 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3884 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3885 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3886 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3887 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3888 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3889 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3890 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3891 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3892 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3893 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3894 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3895 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3896 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3897 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3898 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3899 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3900 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3901 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3902 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3903 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3904 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3905 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3906 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3907 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3908 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3909 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3910 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3911 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3912 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3913 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3914 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3915 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3916 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3917 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3918 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3919 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3920 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3921 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3922 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3923 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3924 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3925 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3926 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3927 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3928 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3929 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3930 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3931 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3932 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3933 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3934 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3935 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3936 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3937 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3938 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3939 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3940 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3941 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3942 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3943 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3944 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3945 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3946 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3947 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3948 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3949 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X3950 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3951 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X3952 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3953 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3954 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3955 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3956 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3957 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3958 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3959 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3960 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3961 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3962 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3963 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3964 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3965 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3966 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3967 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3968 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3969 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3970 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3971 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3972 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3973 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3974 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3975 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3976 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X3977 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3978 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3979 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X3980 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3981 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X3982 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3983 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X3984 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X3985 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3986 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3987 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3988 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3989 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3990 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X3991 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3992 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X3993 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3994 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3995 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3996 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X3997 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3998 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X3999 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4000 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4001 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4002 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4003 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4004 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4005 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4006 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4007 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4008 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4009 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4010 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4011 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4012 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4013 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4014 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4015 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4016 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4017 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4018 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4019 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4020 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4021 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4022 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4023 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4024 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4025 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4026 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4027 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4028 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4029 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4030 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4031 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4032 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4033 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4034 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4035 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4036 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4037 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4038 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4039 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4040 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4041 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4042 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4043 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4044 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4045 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4046 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4047 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4048 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4049 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4050 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4051 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4052 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4053 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4054 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4055 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4056 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4057 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4058 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4059 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4060 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4061 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4062 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4063 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4064 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4065 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4066 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4067 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4068 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4069 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4070 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4071 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4072 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4073 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4074 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4075 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4076 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4077 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4078 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4079 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4080 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4081 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4082 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4083 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4084 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4085 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4086 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4087 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4088 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4089 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4090 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4091 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4092 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4093 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4094 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4095 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4096 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4097 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4098 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4099 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4100 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4101 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4102 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4103 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4104 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4105 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4106 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4107 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4108 VSSA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4109 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4110 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4111 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4112 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4113 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4114 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4115 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4116 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4117 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4118 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4119 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4120 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4121 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4122 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4123 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4124 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4125 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4126 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4127 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4128 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4129 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4130 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4131 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4132 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4133 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4134 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4135 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4136 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4137 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4138 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4139 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4140 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4141 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4142 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4143 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4144 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/D6 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4145 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D6 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4146 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/D6 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4147 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/D6 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4148 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D6 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4149 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4150 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/D6 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4151 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4152 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D7_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=3.16 as=0 ps=0 w=0.5 l=0.5
X4153 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D7 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4154 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D7_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4155 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D7_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.5
X4156 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D7 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4157 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4158 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D7_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4159 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/7_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4160 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1423_1248# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4161 VSSD Din1[0] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X4162 VSSD Din1[0] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4163 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4164 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1353_675# Din1[0] VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X4165 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4166 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1423_1248# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4167 VSSD Din1[1] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X4168 VSSD Din1[1] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4169 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4170 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1353_675# Din1[1] VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X4171 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4172 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1423_1248# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4173 VSSD Din1[2] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X4174 VSSD Din1[2] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4175 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4176 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1353_675# Din1[2] VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X4177 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4178 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1423_1248# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4179 VSSD Din1[3] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X4180 VSSD Din1[3] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4181 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4182 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1353_675# Din1[3] VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X4183 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4184 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1423_1248# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4185 VSSD Din1[4] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X4186 VSSD Din1[4] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4187 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4188 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1353_675# Din1[4] VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X4189 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4190 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1423_1248# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4191 VSSD Din1[5] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X4192 VSSD Din1[5] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4193 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4194 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1353_675# Din1[5] VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X4195 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4196 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1423_1248# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D6 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4197 VSSD Din1[6] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X4198 VSSD Din1[6] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4199 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D6 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4200 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1353_675# Din1[6] VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X4201 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D6 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4202 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1423_1248# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D7 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4203 VSSD Din1[7] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X4204 VSSD Din1[7] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4205 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D7 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4206 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1353_675# Din1[7] VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X4207 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/8_bit_dac_0/D7 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4208 VSSA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_3246_n774# VOUT1 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=2.32 ps=17.2 w=4 l=1
X4209 VOUT1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_3246_n774# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4 l=1
X4210 VDDA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_1618_n334# VOUT1 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=4.64 ps=33.2 w=8 l=1
X4211 VDDA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_394_n920# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_1704_376# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=1.74 ps=13.2 w=2 l=1
X4212 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_1704_376# VOUT1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_1446_376# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=1
X4213 VDDA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_1618_n334# VOUT1 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=8 l=1
X4214 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_408_552# VSSA VSSA sky130_fd_pr__res_generic_nd__hv w=0.48 l=4.46
X4215 VSSA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_1022_n914# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_2158_n774# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.74 ps=13.2 w=4 l=1
X4216 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_2158_n774# VOUT1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_1900_n774# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.58 ps=4.58 w=2 l=1
X4217 VSSA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_2894_292# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_2894_292# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.58 ps=4.58 w=2 l=0.5
X4218 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_1022_n914# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_394_n920# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.6 as=0 ps=0 w=8 l=1
X4219 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_1776_n834# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_408_552# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_1618_n334# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=9.16 as=0.58 ps=4.58 w=2 l=0.5
X4220 VSSA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_1022_n914# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_1446_376# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=9.16 w=2 l=0.5
X4221 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_2894_292# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_408_552# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_1900_n774# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=1.74 ps=13.2 w=2 l=0.5
X4222 VDDA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_408_552# VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=8.32
X4223 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_2416_n774# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_394_n920# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=13.2 as=0 ps=0 w=4 l=1
X4224 VDDA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_394_n920# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_394_n920# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=2.32 ps=16.6 w=8 l=1
X4225 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_1446_376# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_408_552# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_1300_n354# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.58 ps=4.58 w=2 l=0.5
X4226 VOUT1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_3246_n774# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4 l=1
X4227 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_2416_n774# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_2158_n774# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=1
X4228 VOUT1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_1618_n334# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=8 l=1
X4229 VOUT1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_1618_n334# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=8 l=1
X4230 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_1776_n834# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_1704_376# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=1
X4231 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_1618_n334# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_1300_n354# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.6 as=0 ps=0 w=8 l=1
X4232 VSSA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_3246_n774# VOUT1 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4 l=1
X4233 VSSA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_1022_n914# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_1022_n914# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X4234 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_1776_n834# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_1022_n914# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=2 l=0.5
X4235 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_3246_n774# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_2894_292# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X4236 VSSA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_394_n920# VSSA sky130_fd_pr__res_generic_nd__hv w=0.41 l=15.7
X4237 VDDA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_394_n920# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_1900_n774# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4 l=1
X4238 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_3246_n774# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_408_552# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_2416_n774# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X4239 VDDA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_1300_n354# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[1]/opamp_0/a_1300_n354# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=2.32 ps=16.6 w=8 l=1
X4240 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D5_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4241 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4242 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D5_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4243 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D5_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4244 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4245 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4246 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D5_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4247 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4248 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D1_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4249 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4250 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D1_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4251 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D1_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4252 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4253 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4254 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D1_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4255 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4256 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4257 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D0_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4258 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4259 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D0_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4260 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D0_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4261 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4262 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4263 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4264 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4265 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D0_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4266 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4267 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4268 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D0_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4269 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D0_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4270 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4271 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4272 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4273 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4274 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4275 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4276 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4277 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4278 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4279 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4280 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4281 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4282 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4283 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4284 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4285 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4286 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4287 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4288 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4289 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4290 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4291 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4292 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4293 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4294 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4295 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4296 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D2_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4297 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4298 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D2_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4299 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D2_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4300 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4301 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4302 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D2_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4303 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4304 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4305 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4306 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4307 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4308 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4309 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4310 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4311 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4312 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4313 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4314 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4315 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4316 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4317 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4318 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4319 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4320 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4321 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4322 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4323 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4324 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4325 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4326 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4327 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4328 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4329 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4330 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4331 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4332 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4333 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4334 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4335 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4336 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4337 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4338 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4339 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4340 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4341 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4342 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4343 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4344 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4345 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4346 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4347 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4348 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4349 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4350 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4351 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4352 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4353 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4354 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4355 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4356 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4357 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4358 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4359 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4360 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D3_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4361 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4362 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D3_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4363 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D3_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4364 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4365 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4366 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D3_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4367 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4368 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4369 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4370 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4371 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4372 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4373 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4374 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4375 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4376 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4377 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4378 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4379 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4380 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4381 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4382 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4383 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4384 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4385 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4386 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4387 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4388 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4389 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4390 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4391 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4392 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4393 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4394 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4395 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4396 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4397 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4398 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4399 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4400 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4401 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4402 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4403 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4404 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4405 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4406 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4407 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4408 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4409 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4410 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4411 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4412 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4413 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4414 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4415 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4416 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4417 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4418 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4419 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4420 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4421 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4422 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4423 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4424 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4425 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4426 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4427 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4428 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4429 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4430 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4431 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4432 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4433 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4434 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4435 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4436 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4437 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4438 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4439 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4440 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4441 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4442 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4443 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4444 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4445 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4446 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4447 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4448 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4449 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4450 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4451 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4452 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4453 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4454 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4455 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4456 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4457 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4458 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4459 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4460 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4461 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4462 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4463 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4464 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4465 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4466 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4467 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4468 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4469 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4470 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4471 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4472 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4473 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4474 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4475 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4476 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4477 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4478 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4479 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4480 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4481 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4482 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4483 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4484 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4485 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4486 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4487 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4488 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D4_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4489 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4490 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D4_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4491 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D4_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4492 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4493 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4494 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D4_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4495 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4496 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4497 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4498 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4499 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4500 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4501 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4502 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4503 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4504 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4505 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4506 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4507 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4508 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4509 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4510 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4511 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4512 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4513 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4514 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4515 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4516 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4517 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4518 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4519 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4520 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4521 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4522 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4523 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4524 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4525 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4526 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4527 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4528 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4529 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4530 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4531 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4532 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4533 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4534 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4535 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4536 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4537 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4538 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4539 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4540 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4541 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4542 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4543 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4544 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4545 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4546 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4547 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4548 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4549 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4550 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4551 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4552 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4553 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4554 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4555 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4556 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4557 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4558 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4559 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4560 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4561 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4562 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4563 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4564 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4565 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4566 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4567 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4568 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4569 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4570 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4571 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4572 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4573 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4574 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4575 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4576 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4577 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4578 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4579 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4580 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4581 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4582 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4583 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4584 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4585 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4586 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4587 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4588 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4589 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4590 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4591 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4592 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4593 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4594 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4595 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4596 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4597 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4598 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4599 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4600 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4601 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4602 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4603 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4604 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4605 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4606 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4607 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4608 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4609 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4610 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4611 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4612 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4613 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4614 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4615 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4616 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4617 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4618 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4619 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4620 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4621 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4622 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4623 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4624 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4625 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4626 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4627 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4628 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4629 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4630 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4631 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4632 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4633 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4634 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4635 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4636 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4637 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4638 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4639 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4640 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4641 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4642 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4643 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4644 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4645 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4646 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4647 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4648 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4649 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4650 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4651 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4652 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4653 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4654 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4655 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4656 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4657 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4658 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4659 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4660 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4661 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4662 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4663 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4664 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4665 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4666 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4667 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4668 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4669 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4670 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4671 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4672 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4673 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4674 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4675 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4676 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4677 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4678 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4679 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4680 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4681 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4682 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4683 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4684 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4685 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4686 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4687 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4688 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4689 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4690 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4691 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4692 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4693 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4694 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4695 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4696 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4697 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4698 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4699 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4700 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4701 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4702 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4703 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4704 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4705 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4706 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4707 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4708 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4709 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4710 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4711 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4712 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4713 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4714 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4715 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4716 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4717 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4718 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4719 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4720 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4721 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4722 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4723 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4724 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4725 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4726 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4727 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4728 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4729 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4730 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4731 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4732 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4733 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4734 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4735 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4736 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4737 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4738 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4739 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4740 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4741 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4742 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4743 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4744 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4745 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4746 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4747 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4748 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4749 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4750 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4751 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4752 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4753 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4754 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4755 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4756 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4757 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4758 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4759 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4760 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4761 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4762 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4763 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4764 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4765 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4766 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4767 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4768 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4769 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4770 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4771 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4772 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4773 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4774 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4775 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4776 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4777 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4778 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4779 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4780 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4781 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4782 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4783 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4784 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4785 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4786 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4787 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4788 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4789 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4790 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4791 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4792 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4793 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4794 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4795 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4796 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4797 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4798 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4799 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4800 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4801 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4802 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4803 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4804 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4805 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4806 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4807 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4808 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4809 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4810 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4811 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4812 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4813 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4814 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4815 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4816 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4817 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4818 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4819 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4820 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4821 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4822 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4823 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4824 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4825 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4826 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4827 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4828 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4829 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4830 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4831 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4832 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4833 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4834 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4835 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4836 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4837 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4838 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4839 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4840 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4841 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4842 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4843 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4844 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4845 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4846 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4847 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4848 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4849 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4850 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4851 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4852 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4853 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4854 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4855 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4856 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4857 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4858 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4859 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4860 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4861 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4862 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4863 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4864 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4865 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4866 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4867 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4868 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4869 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4870 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4871 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4872 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4873 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4874 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4875 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4876 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4877 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4878 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4879 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4880 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4881 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4882 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4883 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4884 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4885 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4886 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4887 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4888 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4889 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4890 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4891 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4892 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4893 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4894 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4895 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4896 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4897 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4898 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4899 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4900 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4901 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4902 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4903 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4904 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4905 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4906 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4907 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4908 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4909 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4910 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4911 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4912 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4913 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4914 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4915 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4916 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4917 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4918 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4919 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4920 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4921 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4922 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4923 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4924 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4925 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4926 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4927 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4928 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4929 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4930 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4931 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4932 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4933 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4934 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4935 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4936 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4937 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4938 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4939 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4940 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4941 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4942 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4943 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4944 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4945 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4946 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4947 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4948 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4949 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4950 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4951 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4952 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X4953 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4954 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4955 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X4956 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4957 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4958 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4959 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4960 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4961 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4962 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4963 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4964 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4965 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4966 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4967 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4968 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X4969 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4970 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4971 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X4972 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X4973 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4974 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4975 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X4976 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4977 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4978 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4979 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4980 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4981 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4982 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4983 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4984 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X4985 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4986 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4987 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X4988 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4989 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4990 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4991 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4992 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4993 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4994 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X4995 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X4996 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4997 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X4998 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X4999 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5000 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5001 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5002 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5003 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5004 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5005 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5006 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5007 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5008 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5009 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5010 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5011 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5012 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5013 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5014 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5015 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5016 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5017 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5018 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5019 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5020 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5021 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5022 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5023 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5024 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5025 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5026 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5027 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5028 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5029 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5030 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5031 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5032 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5033 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5034 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5035 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5036 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5037 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5038 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5039 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5040 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5041 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5042 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5043 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5044 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5045 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5046 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5047 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5048 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5049 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5050 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5051 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5052 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5053 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5054 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5055 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5056 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5057 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5058 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5059 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5060 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5061 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5062 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5063 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5064 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5065 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5066 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5067 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5068 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5069 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5070 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5071 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5072 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5073 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5074 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5075 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5076 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5077 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5078 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5079 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5080 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5081 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5082 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5083 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5084 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5085 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5086 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5087 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5088 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5089 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5090 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5091 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5092 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5093 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5094 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5095 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5096 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5097 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5098 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5099 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5100 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5101 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5102 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5103 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5104 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5105 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5106 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5107 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5108 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5109 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5110 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5111 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5112 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5113 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5114 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5115 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5116 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5117 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5118 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5119 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5120 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5121 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5122 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5123 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5124 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5125 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5126 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5127 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5128 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5129 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5130 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5131 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5132 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5133 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5134 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5135 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5136 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5137 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5138 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5139 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5140 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5141 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5142 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5143 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5144 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5145 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5146 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5147 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5148 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5149 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5150 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5151 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5152 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5153 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5154 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5155 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5156 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5157 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5158 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5159 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5160 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5161 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5162 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5163 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5164 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5165 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5166 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5167 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5168 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5169 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5170 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5171 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5172 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5173 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5174 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5175 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5176 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5177 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5178 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5179 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5180 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5181 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5182 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5183 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5184 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5185 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5186 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5187 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5188 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5189 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5190 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5191 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5192 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5193 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5194 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5195 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5196 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5197 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5198 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5199 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5200 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5201 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5202 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5203 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5204 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5205 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5206 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5207 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5208 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5209 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5210 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5211 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5212 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5213 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5214 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5215 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5216 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5217 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5218 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5219 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5220 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5221 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5222 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5223 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5224 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5225 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5226 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5227 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5228 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5229 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5230 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5231 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5232 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5233 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5234 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5235 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5236 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5237 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5238 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5239 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5240 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5241 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5242 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5243 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5244 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5245 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5246 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5247 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5248 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D6_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5249 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/D6 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5250 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D6_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5251 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D6_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5252 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/D6 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5253 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5254 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D6_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5255 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5256 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5257 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5258 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5259 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5260 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5261 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5262 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5263 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5264 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5265 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5266 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5267 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5268 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5269 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5270 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5271 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5272 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5273 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5274 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5275 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5276 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5277 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5278 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5279 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5280 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5281 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5282 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5283 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5284 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5285 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5286 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5287 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5288 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5289 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5290 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5291 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5292 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5293 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5294 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5295 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5296 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5297 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5298 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5299 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5300 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5301 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5302 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5303 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5304 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5305 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5306 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5307 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5308 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5309 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5310 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5311 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5312 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5313 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5314 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5315 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5316 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5317 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5318 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5319 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5320 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5321 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5322 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5323 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5324 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5325 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5326 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5327 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5328 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5329 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5330 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5331 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5332 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5333 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5334 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5335 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5336 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5337 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5338 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5339 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5340 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5341 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5342 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5343 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5344 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5345 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5346 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5347 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5348 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5349 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5350 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5351 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5352 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5353 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5354 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5355 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5356 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5357 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5358 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5359 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5360 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5361 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5362 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5363 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5364 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5365 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5366 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5367 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5368 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5369 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5370 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5371 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5372 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5373 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5374 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5375 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5376 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5377 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5378 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5379 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5380 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5381 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5382 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5383 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5384 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5385 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5386 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5387 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5388 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5389 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5390 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5391 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5392 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5393 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5394 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5395 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5396 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5397 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5398 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5399 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5400 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5401 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5402 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5403 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5404 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5405 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5406 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5407 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5408 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5409 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5410 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5411 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5412 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5413 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5414 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5415 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5416 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5417 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5418 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5419 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5420 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5421 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5422 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5423 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5424 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5425 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5426 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5427 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5428 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5429 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5430 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5431 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5432 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5433 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5434 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5435 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5436 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5437 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5438 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5439 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5440 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5441 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5442 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5443 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5444 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5445 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5446 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5447 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5448 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5449 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5450 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5451 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5452 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5453 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5454 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5455 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5456 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5457 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5458 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5459 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5460 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5461 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5462 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5463 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5464 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5465 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5466 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5467 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5468 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5469 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5470 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5471 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5472 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5473 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5474 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5475 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5476 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5477 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5478 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5479 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5480 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5481 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5482 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5483 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5484 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5485 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5486 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5487 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5488 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5489 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5490 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5491 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5492 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5493 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5494 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5495 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5496 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5497 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5498 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5499 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5500 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5501 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5502 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5503 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5504 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5505 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5506 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5507 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5508 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5509 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5510 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5511 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5512 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5513 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5514 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5515 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5516 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5517 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5518 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5519 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5520 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5521 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5522 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5523 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5524 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5525 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5526 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5527 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5528 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5529 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5530 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5531 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5532 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5533 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5534 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5535 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5536 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5537 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5538 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5539 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5540 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5541 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5542 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5543 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5544 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5545 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5546 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5547 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5548 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5549 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5550 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5551 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5552 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5553 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5554 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5555 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5556 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5557 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5558 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5559 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5560 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5561 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5562 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5563 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5564 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5565 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5566 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5567 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5568 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5569 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5570 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5571 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5572 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5573 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5574 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5575 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5576 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5577 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5578 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5579 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5580 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5581 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5582 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5583 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5584 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5585 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5586 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5587 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5588 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5589 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5590 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5591 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5592 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5593 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5594 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5595 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5596 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5597 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5598 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5599 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5600 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5601 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5602 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5603 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5604 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5605 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5606 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5607 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5608 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5609 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5610 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5611 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5612 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5613 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5614 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5615 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5616 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5617 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5618 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5619 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5620 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5621 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5622 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5623 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5624 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5625 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5626 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5627 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5628 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5629 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5630 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5631 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5632 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5633 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5634 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5635 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5636 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5637 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5638 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5639 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5640 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5641 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5642 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5643 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5644 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5645 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5646 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5647 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5648 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5649 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5650 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5651 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5652 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5653 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5654 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5655 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5656 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5657 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5658 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5659 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5660 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5661 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5662 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5663 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5664 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5665 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5666 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5667 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5668 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5669 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5670 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5671 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5672 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5673 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5674 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5675 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5676 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5677 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5678 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5679 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5680 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5681 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5682 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5683 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5684 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5685 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5686 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5687 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5688 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5689 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5690 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5691 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5692 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5693 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5694 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5695 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5696 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5697 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5698 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5699 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5700 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5701 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5702 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5703 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5704 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5705 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5706 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5707 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5708 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5709 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5710 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5711 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5712 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5713 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5714 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5715 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5716 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5717 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5718 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5719 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5720 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5721 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5722 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5723 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5724 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5725 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5726 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5727 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5728 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5729 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5730 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5731 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5732 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5733 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5734 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5735 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5736 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5737 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5738 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5739 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5740 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5741 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5742 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5743 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5744 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5745 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5746 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5747 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5748 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5749 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5750 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5751 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5752 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5753 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5754 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5755 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5756 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5757 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5758 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5759 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5760 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5761 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5762 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5763 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5764 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5765 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5766 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5767 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5768 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5769 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5770 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5771 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5772 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5773 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5774 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5775 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5776 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5777 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5778 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5779 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5780 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5781 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5782 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5783 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5784 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5785 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5786 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5787 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5788 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5789 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5790 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5791 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5792 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5793 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5794 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5795 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5796 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5797 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5798 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5799 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5800 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5801 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5802 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5803 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5804 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5805 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5806 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5807 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5808 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5809 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5810 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5811 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5812 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5813 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5814 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5815 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5816 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5817 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5818 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5819 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5820 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5821 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5822 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5823 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5824 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5825 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5826 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5827 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5828 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5829 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5830 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5831 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5832 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5833 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5834 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5835 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5836 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5837 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5838 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5839 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5840 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5841 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5842 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5843 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5844 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5845 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5846 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5847 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5848 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5849 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5850 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5851 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5852 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5853 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5854 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5855 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5856 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5857 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5858 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5859 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5860 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5861 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5862 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5863 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5864 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5865 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5866 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5867 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5868 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5869 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5870 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5871 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5872 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5873 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5874 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5875 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5876 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5877 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5878 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5879 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5880 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5881 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5882 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5883 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5884 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5885 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5886 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5887 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5888 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5889 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5890 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5891 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5892 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5893 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5894 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5895 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5896 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5897 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5898 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5899 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5900 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5901 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5902 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5903 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5904 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5905 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5906 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5907 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5908 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5909 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5910 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5911 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5912 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5913 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5914 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5915 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5916 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5917 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5918 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5919 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5920 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5921 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5922 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5923 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5924 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5925 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5926 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5927 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5928 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5929 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5930 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5931 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5932 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5933 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5934 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5935 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5936 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5937 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5938 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5939 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5940 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5941 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5942 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5943 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X5944 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5945 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5946 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5947 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5948 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5949 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5950 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5951 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5952 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5953 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5954 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5955 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5956 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5957 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5958 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5959 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5960 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5961 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5962 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5963 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5964 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5965 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5966 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5967 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5968 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X5969 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5970 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5971 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X5972 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5973 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5974 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5975 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5976 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5977 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5978 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5979 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5980 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5981 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5982 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5983 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5984 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X5985 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5986 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5987 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5988 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X5989 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5990 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5991 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5992 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X5993 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5994 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X5995 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X5996 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5997 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X5998 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X5999 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6000 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6001 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6002 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6003 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6004 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6005 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6006 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6007 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6008 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6009 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6010 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6011 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6012 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6013 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6014 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6015 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6016 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6017 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6018 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6019 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6020 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6021 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6022 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6023 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6024 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6025 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6026 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6027 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6028 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6029 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6030 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6031 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6032 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6033 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6034 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6035 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6036 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6037 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6038 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6039 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6040 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6041 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6042 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6043 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6044 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6045 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6046 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6047 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6048 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6049 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6050 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6051 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6052 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6053 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6054 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6055 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6056 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6057 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6058 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6059 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6060 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6061 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6062 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6063 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6064 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6065 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6066 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6067 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6068 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6069 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6070 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6071 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6072 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6073 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6074 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6075 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6076 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6077 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6078 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6079 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6080 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6081 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6082 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6083 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6084 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6085 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6086 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6087 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6088 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6089 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6090 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6091 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6092 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6093 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6094 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6095 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6096 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6097 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6098 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6099 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6100 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6101 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6102 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6103 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6104 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6105 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6106 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6107 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6108 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6109 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6110 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6111 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6112 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6113 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6114 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6115 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6116 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6117 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6118 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6119 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6120 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6121 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6122 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6123 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6124 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6125 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6126 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6127 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6128 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6129 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6130 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6131 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6132 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6133 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6134 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6135 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6136 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6137 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6138 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6139 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6140 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6141 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6142 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6143 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6144 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6145 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6146 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6147 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6148 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6149 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6150 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6151 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6152 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6153 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6154 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6155 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6156 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6157 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6158 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6159 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6160 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6161 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6162 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6163 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6164 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6165 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6166 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6167 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6168 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6169 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6170 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6171 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6172 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6173 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6174 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6175 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6176 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6177 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6178 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6179 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6180 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6181 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6182 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6183 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6184 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6185 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6186 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6187 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6188 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6189 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6190 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6191 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6192 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6193 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6194 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6195 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6196 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6197 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6198 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6199 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6200 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6201 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6202 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6203 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6204 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6205 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6206 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6207 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6208 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6209 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6210 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6211 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6212 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6213 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6214 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6215 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6216 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6217 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6218 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6219 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6220 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6221 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6222 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6223 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6224 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6225 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6226 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6227 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6228 VSSA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6229 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6230 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6231 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6232 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6233 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6234 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6235 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6236 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6237 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6238 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6239 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6240 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6241 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6242 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6243 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6244 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6245 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6246 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6247 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6248 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6249 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6250 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6251 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6252 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6253 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6254 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6255 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6256 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6257 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6258 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6259 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6260 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6261 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6262 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6263 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6264 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/D6 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6265 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D6 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6266 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/D6 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6267 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/D6 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6268 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D6 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6269 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6270 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/D6 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6271 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6272 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D7_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=3.16 as=0 ps=0 w=0.5 l=0.5
X6273 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D7 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6274 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D7_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6275 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D7_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.5
X6276 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D7 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6277 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6278 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D7_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6279 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/7_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6280 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1423_1248# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6281 VSSD Din2[0] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X6282 VSSD Din2[0] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6283 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6284 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1353_675# Din2[0] VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X6285 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6286 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1423_1248# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6287 VSSD Din2[1] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X6288 VSSD Din2[1] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6289 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6290 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1353_675# Din2[1] VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X6291 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6292 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1423_1248# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6293 VSSD Din2[2] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X6294 VSSD Din2[2] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6295 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6296 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1353_675# Din2[2] VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X6297 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6298 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1423_1248# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6299 VSSD Din2[3] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X6300 VSSD Din2[3] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6301 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6302 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1353_675# Din2[3] VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X6303 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6304 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1423_1248# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6305 VSSD Din2[4] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X6306 VSSD Din2[4] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6307 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6308 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1353_675# Din2[4] VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X6309 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6310 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1423_1248# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6311 VSSD Din2[5] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X6312 VSSD Din2[5] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6313 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6314 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1353_675# Din2[5] VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X6315 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6316 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1423_1248# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D6 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6317 VSSD Din2[6] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X6318 VSSD Din2[6] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6319 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D6 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6320 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1353_675# Din2[6] VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X6321 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D6 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6322 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1423_1248# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D7 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6323 VSSD Din2[7] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X6324 VSSD Din2[7] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6325 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D7 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6326 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1353_675# Din2[7] VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X6327 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/8_bit_dac_0/D7 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6328 VSSA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_3246_n774# VOUT2 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=2.32 ps=17.2 w=4 l=1
X6329 VOUT2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_3246_n774# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4 l=1
X6330 VDDA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_1618_n334# VOUT2 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=4.64 ps=33.2 w=8 l=1
X6331 VDDA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_394_n920# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_1704_376# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=1.74 ps=13.2 w=2 l=1
X6332 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_1704_376# VOUT2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_1446_376# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=1
X6333 VDDA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_1618_n334# VOUT2 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=8 l=1
X6334 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_408_552# VSSA VSSA sky130_fd_pr__res_generic_nd__hv w=0.48 l=4.46
X6335 VSSA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_1022_n914# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_2158_n774# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.74 ps=13.2 w=4 l=1
X6336 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_2158_n774# VOUT2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_1900_n774# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.58 ps=4.58 w=2 l=1
X6337 VSSA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_2894_292# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_2894_292# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.58 ps=4.58 w=2 l=0.5
X6338 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_1022_n914# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_394_n920# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.6 as=0 ps=0 w=8 l=1
X6339 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_1776_n834# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_408_552# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_1618_n334# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=9.16 as=0.58 ps=4.58 w=2 l=0.5
X6340 VSSA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_1022_n914# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_1446_376# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=9.16 w=2 l=0.5
X6341 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_2894_292# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_408_552# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_1900_n774# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=1.74 ps=13.2 w=2 l=0.5
X6342 VDDA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_408_552# VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=8.32
X6343 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_2416_n774# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_394_n920# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=13.2 as=0 ps=0 w=4 l=1
X6344 VDDA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_394_n920# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_394_n920# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=2.32 ps=16.6 w=8 l=1
X6345 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_1446_376# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_408_552# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_1300_n354# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.58 ps=4.58 w=2 l=0.5
X6346 VOUT2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_3246_n774# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4 l=1
X6347 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_2416_n774# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_2158_n774# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=1
X6348 VOUT2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_1618_n334# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=8 l=1
X6349 VOUT2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_1618_n334# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=8 l=1
X6350 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_1776_n834# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_1704_376# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=1
X6351 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_1618_n334# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_1300_n354# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.6 as=0 ps=0 w=8 l=1
X6352 VSSA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_3246_n774# VOUT2 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4 l=1
X6353 VSSA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_1022_n914# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_1022_n914# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X6354 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_1776_n834# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_1022_n914# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=2 l=0.5
X6355 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_3246_n774# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_2894_292# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X6356 VSSA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_394_n920# VSSA sky130_fd_pr__res_generic_nd__hv w=0.41 l=15.7
X6357 VDDA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_394_n920# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_1900_n774# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4 l=1
X6358 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_3246_n774# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_408_552# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_2416_n774# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X6359 VDDA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_1300_n354# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[2]/opamp_0/a_1300_n354# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=2.32 ps=16.6 w=8 l=1
X6360 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D5_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6361 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6362 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D5_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6363 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D5_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6364 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6365 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6366 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D5_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6367 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6368 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D1_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6369 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6370 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D1_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6371 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D1_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6372 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6373 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6374 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D1_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6375 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6376 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6377 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D0_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6378 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6379 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D0_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6380 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D0_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6381 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6382 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6383 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6384 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6385 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D0_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6386 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6387 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6388 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D0_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6389 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D0_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6390 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6391 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6392 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6393 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6394 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6395 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6396 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6397 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6398 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6399 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6400 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6401 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6402 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6403 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6404 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6405 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6406 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6407 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6408 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6409 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6410 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6411 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6412 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6413 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6414 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6415 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6416 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D2_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6417 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6418 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D2_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6419 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D2_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6420 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6421 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6422 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D2_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6423 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6424 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6425 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6426 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6427 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6428 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6429 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6430 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6431 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6432 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6433 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6434 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6435 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6436 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6437 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6438 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6439 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6440 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6441 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6442 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6443 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6444 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6445 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6446 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6447 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6448 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6449 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6450 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6451 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6452 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6453 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6454 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6455 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6456 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6457 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6458 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6459 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6460 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6461 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6462 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6463 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6464 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6465 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6466 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6467 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6468 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6469 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6470 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6471 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6472 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6473 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6474 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6475 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6476 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6477 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6478 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6479 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6480 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D3_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6481 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6482 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D3_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6483 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D3_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6484 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6485 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6486 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D3_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6487 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6488 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6489 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6490 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6491 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6492 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6493 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6494 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6495 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6496 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6497 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6498 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6499 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6500 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6501 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6502 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6503 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6504 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6505 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6506 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6507 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6508 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6509 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6510 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6511 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6512 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6513 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6514 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6515 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6516 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6517 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6518 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6519 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6520 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6521 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6522 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6523 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6524 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6525 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6526 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6527 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6528 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6529 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6530 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6531 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6532 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6533 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6534 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6535 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6536 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6537 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6538 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6539 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6540 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6541 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6542 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6543 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6544 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6545 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6546 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6547 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6548 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6549 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6550 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6551 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6552 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6553 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6554 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6555 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6556 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6557 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6558 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6559 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6560 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6561 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6562 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6563 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6564 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6565 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6566 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6567 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6568 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6569 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6570 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6571 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6572 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6573 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6574 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6575 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6576 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6577 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6578 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6579 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6580 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6581 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6582 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6583 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6584 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6585 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6586 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6587 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6588 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6589 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6590 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6591 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6592 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6593 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6594 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6595 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6596 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6597 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6598 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6599 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6600 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6601 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6602 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6603 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6604 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6605 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6606 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6607 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6608 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D4_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6609 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6610 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D4_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6611 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D4_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6612 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6613 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6614 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D4_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6615 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6616 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6617 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6618 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6619 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6620 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6621 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6622 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6623 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6624 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6625 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6626 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6627 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6628 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6629 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6630 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6631 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6632 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6633 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6634 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6635 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6636 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6637 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6638 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6639 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6640 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6641 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6642 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6643 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6644 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6645 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6646 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6647 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6648 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6649 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6650 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6651 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6652 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6653 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6654 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6655 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6656 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6657 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6658 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6659 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6660 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6661 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6662 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6663 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6664 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6665 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6666 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6667 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6668 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6669 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6670 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6671 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6672 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6673 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6674 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6675 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6676 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6677 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6678 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6679 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6680 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6681 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6682 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6683 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6684 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6685 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6686 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6687 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6688 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6689 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6690 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6691 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6692 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6693 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6694 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6695 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6696 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6697 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6698 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6699 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6700 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6701 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6702 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6703 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6704 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6705 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6706 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6707 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6708 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6709 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6710 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6711 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6712 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6713 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6714 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6715 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6716 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6717 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6718 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6719 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6720 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6721 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6722 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6723 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6724 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6725 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6726 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6727 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6728 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6729 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6730 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6731 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6732 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6733 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6734 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6735 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6736 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6737 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6738 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6739 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6740 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6741 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6742 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6743 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6744 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6745 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6746 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6747 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6748 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6749 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6750 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6751 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6752 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6753 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6754 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6755 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6756 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6757 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6758 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6759 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6760 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6761 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6762 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6763 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6764 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6765 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6766 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6767 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6768 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6769 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6770 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6771 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6772 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6773 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6774 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6775 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6776 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6777 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6778 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6779 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6780 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6781 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6782 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6783 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6784 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6785 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6786 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6787 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6788 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6789 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6790 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6791 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6792 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6793 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6794 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6795 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6796 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6797 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6798 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6799 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6800 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6801 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6802 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6803 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6804 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6805 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6806 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6807 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6808 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6809 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6810 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6811 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6812 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6813 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6814 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6815 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6816 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6817 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6818 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6819 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6820 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6821 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6822 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6823 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6824 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6825 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6826 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6827 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6828 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6829 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6830 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6831 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6832 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6833 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6834 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6835 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6836 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6837 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6838 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6839 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6840 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6841 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6842 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6843 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6844 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6845 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6846 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6847 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6848 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6849 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6850 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6851 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6852 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6853 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6854 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6855 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6856 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6857 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6858 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6859 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6860 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6861 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6862 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6863 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6864 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6865 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6866 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6867 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6868 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6869 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6870 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6871 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6872 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6873 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6874 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6875 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6876 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6877 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6878 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6879 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6880 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6881 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6882 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6883 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6884 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6885 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6886 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6887 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6888 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6889 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6890 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6891 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6892 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6893 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6894 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6895 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6896 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6897 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6898 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6899 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6900 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6901 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6902 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6903 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6904 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6905 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6906 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6907 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6908 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6909 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6910 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6911 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6912 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6913 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6914 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6915 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6916 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6917 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6918 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6919 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6920 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6921 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6922 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6923 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6924 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6925 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6926 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6927 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6928 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6929 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6930 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6931 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6932 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6933 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6934 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6935 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6936 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6937 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6938 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6939 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6940 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6941 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6942 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6943 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6944 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6945 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6946 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6947 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6948 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6949 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6950 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6951 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6952 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6953 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6954 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6955 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6956 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6957 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6958 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6959 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6960 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6961 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6962 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6963 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6964 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6965 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6966 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6967 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6968 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X6969 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6970 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6971 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6972 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X6973 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6974 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6975 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X6976 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6977 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6978 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6979 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6980 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6981 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6982 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6983 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6984 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6985 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6986 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6987 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X6988 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6989 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X6990 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6991 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6992 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X6993 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6994 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X6995 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X6996 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6997 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X6998 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X6999 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7000 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7001 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7002 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7003 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7004 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7005 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7006 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7007 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7008 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7009 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7010 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7011 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7012 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7013 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7014 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7015 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7016 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7017 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7018 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7019 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7020 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7021 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7022 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7023 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7024 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7025 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7026 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7027 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7028 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7029 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7030 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7031 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7032 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7033 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7034 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7035 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7036 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7037 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7038 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7039 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7040 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7041 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7042 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7043 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7044 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7045 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7046 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7047 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7048 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7049 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7050 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7051 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7052 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7053 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7054 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7055 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7056 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7057 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7058 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7059 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7060 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7061 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7062 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7063 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7064 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7065 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7066 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7067 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7068 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7069 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7070 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7071 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7072 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7073 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7074 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7075 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7076 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7077 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7078 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7079 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7080 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7081 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7082 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7083 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7084 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7085 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7086 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7087 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7088 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7089 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7090 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7091 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7092 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7093 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7094 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7095 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7096 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7097 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7098 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7099 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7100 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7101 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7102 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7103 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7104 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7105 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7106 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7107 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7108 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7109 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7110 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7111 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7112 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7113 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7114 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7115 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7116 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7117 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7118 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7119 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7120 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7121 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7122 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7123 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7124 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7125 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7126 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7127 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7128 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7129 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7130 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7131 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7132 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7133 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7134 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7135 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7136 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7137 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7138 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7139 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7140 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7141 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7142 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7143 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7144 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7145 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7146 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7147 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7148 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7149 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7150 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7151 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7152 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7153 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7154 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7155 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7156 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7157 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7158 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7159 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7160 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7161 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7162 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7163 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7164 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7165 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7166 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7167 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7168 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7169 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7170 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7171 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7172 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7173 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7174 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7175 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7176 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7177 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7178 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7179 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7180 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7181 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7182 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7183 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7184 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7185 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7186 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7187 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7188 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7189 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7190 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7191 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7192 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7193 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7194 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7195 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7196 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7197 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7198 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7199 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7200 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7201 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7202 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7203 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7204 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7205 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7206 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7207 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7208 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7209 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7210 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7211 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7212 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7213 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7214 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7215 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7216 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7217 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7218 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7219 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7220 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7221 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7222 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7223 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7224 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7225 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7226 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7227 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7228 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7229 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7230 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7231 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7232 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7233 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7234 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7235 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7236 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7237 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7238 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7239 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7240 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7241 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7242 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7243 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7244 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7245 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7246 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7247 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7248 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7249 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7250 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7251 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7252 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7253 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7254 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7255 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7256 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7257 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7258 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7259 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7260 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7261 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7262 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7263 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7264 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7265 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7266 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7267 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7268 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7269 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7270 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7271 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7272 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7273 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7274 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7275 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7276 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7277 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7278 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7279 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7280 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7281 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7282 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7283 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7284 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7285 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7286 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7287 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7288 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7289 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7290 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7291 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7292 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7293 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7294 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7295 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7296 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7297 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7298 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7299 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7300 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7301 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7302 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7303 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7304 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7305 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7306 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7307 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7308 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7309 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7310 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7311 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7312 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7313 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7314 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7315 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7316 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7317 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7318 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7319 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7320 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7321 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7322 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7323 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7324 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7325 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7326 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7327 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7328 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7329 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7330 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7331 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7332 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7333 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7334 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7335 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7336 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7337 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7338 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7339 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7340 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7341 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7342 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7343 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7344 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7345 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7346 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7347 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7348 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7349 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7350 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7351 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7352 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7353 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7354 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7355 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7356 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7357 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7358 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7359 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7360 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7361 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7362 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7363 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7364 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7365 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7366 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7367 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7368 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D6_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7369 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/D6 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7370 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D6_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7371 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D6_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7372 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/D6 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7373 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7374 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D6_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7375 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7376 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7377 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7378 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7379 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7380 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7381 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7382 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7383 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7384 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7385 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7386 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7387 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7388 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7389 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7390 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7391 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7392 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7393 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7394 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7395 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7396 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7397 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7398 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7399 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7400 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7401 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7402 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7403 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7404 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7405 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7406 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7407 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7408 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7409 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7410 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7411 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7412 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7413 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7414 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7415 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7416 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7417 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7418 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7419 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7420 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7421 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7422 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7423 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7424 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7425 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7426 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7427 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7428 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7429 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7430 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7431 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7432 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7433 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7434 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7435 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7436 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7437 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7438 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7439 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7440 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7441 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7442 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7443 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7444 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7445 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7446 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7447 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7448 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7449 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7450 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7451 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7452 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7453 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7454 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7455 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7456 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7457 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7458 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7459 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7460 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7461 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7462 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7463 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7464 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7465 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7466 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7467 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7468 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7469 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7470 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7471 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7472 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7473 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7474 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7475 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7476 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7477 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7478 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7479 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7480 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7481 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7482 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7483 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7484 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7485 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7486 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7487 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7488 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7489 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7490 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7491 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7492 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7493 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7494 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7495 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7496 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7497 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7498 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7499 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7500 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7501 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7502 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7503 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7504 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7505 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7506 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7507 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7508 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7509 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7510 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7511 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7512 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7513 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7514 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7515 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7516 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7517 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7518 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7519 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7520 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7521 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7522 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7523 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7524 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7525 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7526 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7527 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7528 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7529 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7530 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7531 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7532 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7533 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7534 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7535 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7536 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7537 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7538 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7539 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7540 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7541 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7542 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7543 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7544 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7545 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7546 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7547 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7548 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7549 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7550 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7551 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7552 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7553 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7554 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7555 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7556 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7557 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7558 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7559 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7560 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7561 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7562 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7563 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7564 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7565 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7566 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7567 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7568 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7569 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7570 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7571 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7572 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7573 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7574 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7575 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7576 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7577 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7578 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7579 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7580 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7581 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7582 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7583 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7584 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7585 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7586 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7587 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7588 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7589 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7590 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7591 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7592 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7593 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7594 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7595 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7596 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7597 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7598 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7599 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7600 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7601 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7602 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7603 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7604 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7605 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7606 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7607 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7608 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7609 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7610 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7611 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7612 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7613 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7614 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7615 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7616 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7617 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7618 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7619 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7620 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7621 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7622 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7623 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7624 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7625 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7626 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7627 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7628 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7629 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7630 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7631 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7632 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7633 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7634 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7635 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7636 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7637 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7638 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7639 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7640 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7641 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7642 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7643 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7644 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7645 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7646 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7647 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7648 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7649 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7650 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7651 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7652 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7653 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7654 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7655 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7656 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7657 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7658 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7659 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7660 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7661 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7662 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7663 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7664 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7665 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7666 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7667 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7668 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7669 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7670 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7671 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7672 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7673 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7674 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7675 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7676 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7677 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7678 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7679 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7680 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7681 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7682 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7683 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7684 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7685 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7686 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7687 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7688 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7689 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7690 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7691 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7692 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7693 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7694 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7695 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7696 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7697 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7698 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7699 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7700 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7701 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7702 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7703 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7704 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7705 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7706 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7707 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7708 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7709 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7710 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7711 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7712 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7713 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7714 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7715 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7716 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7717 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7718 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7719 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7720 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7721 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7722 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7723 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7724 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7725 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7726 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7727 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7728 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7729 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7730 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7731 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7732 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7733 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7734 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7735 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7736 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7737 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7738 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7739 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7740 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7741 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7742 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7743 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7744 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7745 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7746 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7747 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7748 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7749 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7750 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7751 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7752 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7753 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7754 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7755 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7756 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7757 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7758 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7759 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7760 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7761 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7762 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7763 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7764 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7765 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7766 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7767 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7768 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7769 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7770 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7771 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7772 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7773 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7774 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7775 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7776 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7777 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7778 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7779 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7780 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7781 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7782 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7783 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7784 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7785 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7786 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7787 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7788 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7789 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7790 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7791 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7792 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7793 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7794 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7795 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7796 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7797 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7798 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7799 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7800 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7801 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7802 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7803 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7804 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7805 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7806 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7807 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7808 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7809 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7810 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7811 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7812 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7813 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7814 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7815 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7816 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7817 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7818 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7819 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7820 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7821 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7822 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7823 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7824 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7825 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7826 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7827 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7828 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7829 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7830 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7831 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7832 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7833 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7834 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7835 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7836 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7837 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7838 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7839 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7840 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7841 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7842 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7843 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7844 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7845 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7846 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7847 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7848 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7849 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7850 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7851 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7852 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7853 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7854 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7855 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7856 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7857 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7858 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7859 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7860 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7861 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7862 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7863 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7864 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7865 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7866 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7867 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7868 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7869 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7870 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7871 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7872 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7873 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7874 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7875 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7876 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7877 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7878 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7879 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7880 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7881 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7882 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7883 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7884 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7885 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7886 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7887 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7888 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7889 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7890 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7891 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7892 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7893 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7894 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7895 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7896 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7897 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7898 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7899 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7900 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7901 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7902 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7903 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7904 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7905 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7906 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7907 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7908 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7909 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7910 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7911 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7912 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7913 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7914 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7915 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7916 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7917 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7918 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7919 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7920 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7921 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7922 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7923 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7924 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7925 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7926 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7927 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7928 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7929 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7930 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7931 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7932 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7933 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7934 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7935 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7936 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7937 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7938 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7939 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7940 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7941 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7942 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7943 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X7944 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7945 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7946 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7947 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7948 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7949 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7950 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7951 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7952 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7953 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7954 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7955 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7956 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7957 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7958 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7959 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7960 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7961 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7962 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7963 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7964 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7965 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7966 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7967 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7968 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X7969 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7970 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7971 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X7972 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7973 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7974 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7975 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7976 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7977 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7978 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7979 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7980 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7981 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7982 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7983 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7984 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X7985 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7986 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7987 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X7988 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X7989 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7990 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7991 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7992 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X7993 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7994 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X7995 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X7996 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7997 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X7998 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X7999 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8000 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8001 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8002 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8003 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8004 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8005 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X8006 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8007 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8008 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X8009 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8010 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8011 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X8012 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8013 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8014 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8015 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8016 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8017 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8018 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8019 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8020 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8021 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8022 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8023 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8024 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8025 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8026 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8027 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8028 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8029 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8030 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8031 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8032 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X8033 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8034 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8035 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X8036 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8037 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8038 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8039 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8040 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8041 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8042 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8043 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8044 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8045 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8046 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8047 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8048 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8049 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8050 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8051 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8052 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8053 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8054 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8055 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8056 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8057 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8058 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8059 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8060 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8061 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X8062 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8063 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8064 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X8065 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8066 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8067 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X8068 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8069 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8070 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8071 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8072 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8073 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8074 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8075 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8076 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8077 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8078 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8079 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8080 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8081 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8082 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8083 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8084 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8085 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8086 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8087 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8088 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X8089 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8090 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8091 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X8092 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8093 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8094 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8095 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8096 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8097 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8098 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8099 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8100 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8101 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8102 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8103 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8104 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8105 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8106 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8107 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8108 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8109 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8110 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8111 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8112 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8113 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8114 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8115 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8116 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8117 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X8118 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8119 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8120 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8121 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8122 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8123 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8124 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8125 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X8126 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8127 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8128 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X8129 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8130 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8131 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8132 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8133 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X8134 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8135 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8136 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X8137 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8138 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8139 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X8140 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8141 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8142 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8143 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8144 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8145 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8146 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8147 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8148 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8149 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8150 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8151 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8152 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8153 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8154 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8155 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8156 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8157 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8158 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8159 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8160 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X8161 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8162 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8163 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X8164 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8165 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8166 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8167 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8168 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8169 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8170 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8171 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8172 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8173 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8174 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8175 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8176 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8177 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8178 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8179 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8180 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8181 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8182 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8183 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8184 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8185 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8186 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8187 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8188 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8189 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X8190 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8191 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8192 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X8193 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8194 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8195 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X8196 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8197 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8198 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8199 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8200 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8201 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8202 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8203 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8204 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8205 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8206 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8207 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8208 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8209 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8210 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8211 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8212 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8213 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8214 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8215 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8216 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X8217 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8218 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8219 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X8220 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8221 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8222 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8223 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8224 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8225 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8226 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8227 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8228 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8229 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8230 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8231 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8232 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8233 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8234 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8235 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8236 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8237 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8238 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8239 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8240 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8241 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8242 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8243 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8244 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8245 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X8246 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8247 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8248 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8249 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8250 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8251 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8252 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8253 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X8254 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8255 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8256 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X8257 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8258 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8259 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X8260 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8261 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8262 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8263 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8264 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8265 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8266 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8267 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8268 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8269 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8270 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8271 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8272 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8273 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8274 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8275 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8276 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8277 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8278 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8279 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8280 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X8281 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8282 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8283 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X8284 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8285 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8286 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8287 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8288 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8289 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8290 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8291 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8292 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8293 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8294 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8295 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8296 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8297 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8298 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8299 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8300 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8301 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8302 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8303 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8304 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8305 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8306 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8307 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8308 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8309 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X8310 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8311 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8312 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X8313 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8314 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8315 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X8316 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8317 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8318 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8319 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8320 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8321 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8322 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8323 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8324 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8325 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8326 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8327 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8328 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8329 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8330 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8331 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8332 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8333 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8334 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8335 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8336 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X8337 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8338 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8339 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X8340 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8341 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8342 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8343 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8344 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8345 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8346 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8347 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8348 VSSA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8349 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8350 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8351 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X8352 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X8353 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8354 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8355 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X8356 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X8357 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8358 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8359 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8360 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8361 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8362 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8363 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8364 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8365 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X8366 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8367 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8368 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8369 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8370 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8371 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8372 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8373 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X8374 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8375 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8376 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X8377 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8378 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8379 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8380 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8381 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X8382 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8383 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8384 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/D6 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X8385 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D6 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8386 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/D6 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8387 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/D6 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X8388 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D6 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8389 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X8390 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/D6 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8391 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8392 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D7_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=3.16 as=0 ps=0 w=0.5 l=0.5
X8393 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D7 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8394 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D7_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8395 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D7_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.5
X8396 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D7 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8397 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[1]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X8398 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D7_BUF 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8399 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/7_bit_dac_0[0]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/switch_n_3v3_1/DX_ 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X8400 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1423_1248# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8401 VSSD Din3[0] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X8402 VSSD Din3[0] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8403 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8404 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1353_675# Din3[0] VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X8405 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D0 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[0]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8406 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1423_1248# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8407 VSSD Din3[1] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X8408 VSSD Din3[1] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8409 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8410 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1353_675# Din3[1] VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X8411 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D1 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[1]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8412 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1423_1248# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8413 VSSD Din3[2] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X8414 VSSD Din3[2] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8415 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8416 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1353_675# Din3[2] VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X8417 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D2 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[2]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8418 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1423_1248# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8419 VSSD Din3[3] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X8420 VSSD Din3[3] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8421 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8422 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1353_675# Din3[3] VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X8423 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[3]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8424 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1423_1248# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8425 VSSD Din3[4] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X8426 VSSD Din3[4] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8427 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8428 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1353_675# Din3[4] VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X8429 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D4 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[4]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8430 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1423_1248# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8431 VSSD Din3[5] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X8432 VSSD Din3[5] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8433 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8434 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1353_675# Din3[5] VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X8435 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D5 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[5]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8436 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1423_1248# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D6 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8437 VSSD Din3[6] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X8438 VSSD Din3[6] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8439 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D6 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8440 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1353_675# Din3[6] VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X8441 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D6 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[6]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8442 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1423_1248# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D7 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8443 VSSD Din3[7] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X8444 VSSD Din3[7] 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X8445 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D7 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X8446 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1353_675# Din3[7] VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X8447 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/8_bit_dac_0/D7 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/level_tx_8bit_0/level_tx_1bit_0[7]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X8448 VSSA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_3246_n774# VOUT3 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=2.32 ps=17.2 w=4 l=1
X8449 VOUT3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_3246_n774# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4 l=1
X8450 VDDA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_1618_n334# VOUT3 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=4.64 ps=33.2 w=8 l=1
X8451 VDDA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_394_n920# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_1704_376# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=1.74 ps=13.2 w=2 l=1
X8452 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_1704_376# VOUT3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_1446_376# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=1
X8453 VDDA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_1618_n334# VOUT3 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=8 l=1
X8454 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_408_552# VSSA VSSA sky130_fd_pr__res_generic_nd__hv w=0.48 l=4.46
X8455 VSSA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_1022_n914# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_2158_n774# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.74 ps=13.2 w=4 l=1
X8456 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_2158_n774# VOUT3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_1900_n774# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.58 ps=4.58 w=2 l=1
X8457 VSSA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_2894_292# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_2894_292# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.58 ps=4.58 w=2 l=0.5
X8458 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_1022_n914# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_394_n920# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.6 as=0 ps=0 w=8 l=1
X8459 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_1776_n834# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_408_552# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_1618_n334# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=9.16 as=0.58 ps=4.58 w=2 l=0.5
X8460 VSSA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_1022_n914# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_1446_376# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=9.16 w=2 l=0.5
X8461 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_2894_292# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_408_552# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_1900_n774# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=1.74 ps=13.2 w=2 l=0.5
X8462 VDDA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_408_552# VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=8.32
X8463 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_2416_n774# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_394_n920# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=13.2 as=0 ps=0 w=4 l=1
X8464 VDDA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_394_n920# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_394_n920# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=2.32 ps=16.6 w=8 l=1
X8465 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_1446_376# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_408_552# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_1300_n354# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.58 ps=4.58 w=2 l=0.5
X8466 VOUT3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_3246_n774# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4 l=1
X8467 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_2416_n774# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_2158_n774# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=1
X8468 VOUT3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_1618_n334# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=8 l=1
X8469 VOUT3 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_1618_n334# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=8 l=1
X8470 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_1776_n834# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/VOUT 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_1704_376# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0 ps=0 w=4 l=1
X8471 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_1618_n334# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_1300_n354# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.6 as=0 ps=0 w=8 l=1
X8472 VSSA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_3246_n774# VOUT3 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4 l=1
X8473 VSSA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_1022_n914# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_1022_n914# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=1.16 ps=8.58 w=4 l=0.5
X8474 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_1776_n834# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_1022_n914# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=2 l=0.5
X8475 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_3246_n774# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_2894_292# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X8476 VSSA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_394_n920# VSSA sky130_fd_pr__res_generic_nd__hv w=0.41 l=15.7
X8477 VDDA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_394_n920# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_1900_n774# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=4 l=1
X8478 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_3246_n774# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_408_552# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_2416_n774# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X8479 VDDA 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_1300_n354# 4x8_bit_dac_0/8_bit_dac_tx_buffer_0[3]/opamp_0/a_1300_n354# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=2.32 ps=16.6 w=8 l=1
.ends

**********************************************************************************
X1 VDDA VSSA VCCD VSSD VREFH Din0[0] Din0[1] Din0[2] Din0[3] Din0[4]
+ Din0[5] Din0[6] Din0[7] VOUT0 Din1[0] Din1[1] Din1[2] Din1[3] Din1[4] Din1[5] Din1[6]
+ Din1[7] VOUT1 Din2[0] Din2[1] Din2[2] Din2[3] Din2[4] Din2[5] Din2[6] Din2[7] VOUT2
+ Din3[0] Din3[1] Din3[2] Din3[3] Din3[4] Din3[5] Din3[6] Din3[7] VOUT3
+ dac_top
**********************************************************************************

.param mc_mm_switch=0
.param mc_pr_switch=0
.lib "/foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice.tt.red" tt


V1 VDDA 0 dc 3.3
V2 VSSA 0 dc 0
V3 VCCD 0 dc 1.8
V4 VSSD 0 dc 0
V6 VREFH 0 dc 3

V7  Din0[0] 0 pulse(0 1.8 0ns 0.1ns 0.1ns 1us 2us)
V8  Din0[1] 0 pulse(0 1.8 0ns 0.1ns 0.1ns 2us 4us)
V9  Din0[2] 0 pulse(0 1.8 0ns 0.1ns 0.1ns 4us 8us)
V10 Din0[3] 0 pulse(0 1.8 0ns 0.1ns 0.1ns 8us 16us)
V11 Din0[4] 0 pulse(0 1.8 0ns 0.1ns 0.1ns 16us 32us)
V12 Din0[5] 0 pulse(0 1.8 0ns 0.1ns 0.1ns 32us 64us)
V13 Din0[6] 0 pulse(0 1.8 0ns 0.1ns 0.1ns 64us 128us)
V14 Din0[7] 0 pulse(0 1.8 0ns 0.1ns 0.1ns 128us 256us)

V15 Din1[0] 0 pulse(0 1.8 1us 0.1ns 0.1ns 1us 2us)
V16 Din1[1] 0 pulse(0 1.8 2us 0.1ns 0.1ns 2us 4us)
V17 Din1[2] 0 pulse(0 1.8 4us 0.1ns 0.1ns 4us 8us)
V18 Din1[3] 0 pulse(0 1.8 8us 0.1ns 0.1ns 8us 16us)
V19 Din1[4] 0 pulse(0 1.8 16us 0.1ns 0.1ns 16us 32us)
V20 Din1[5] 0 pulse(0 1.8 32us 0.1ns 0.1ns 32us 64us)
V21 Din1[6] 0 pulse(0 1.8 64us 0.1ns 0.1ns 64us 128us)
V22 Din1[7] 0 pulse(0 1.8 128us 0.1ns 0.1ns 128us 256us)

V23 Din2[0] 0 pulse(0 1.8 0ns 0.1ns 0.1ns 1us 2us)
V24 Din2[1] 0 pulse(0 1.8 0ns 0.1ns 0.1ns 2us 4us)
V25 Din2[2] 0 pulse(0 1.8 0ns 0.1ns 0.1ns 4us 8us)
V26 Din2[3] 0 pulse(0 1.8 0ns 0.1ns 0.1ns 8us 16us)
V27 Din2[4] 0 pulse(0 1.8 0ns 0.1ns 0.1ns 16us 32us)
V28 Din2[5] 0 pulse(0 1.8 0ns 0.1ns 0.1ns 32us 64us)
V29 Din2[6] 0 pulse(0 1.8 0ns 0.1ns 0.1ns 64us 128us)
V30 Din2[7] 0 pulse(0 1.8 0ns 0.1ns 0.1ns 128us 256us)

V31 Din3[0] 0 pulse(0 1.8 1us 0.1ns 0.1ns 1us 2us)
V32 Din3[1] 0 pulse(0 1.8 2us 0.1ns 0.1ns 2us 4us)
V33 Din3[2] 0 pulse(0 1.8 4us 0.1ns 0.1ns 4us 8us)
V34 Din3[3] 0 pulse(0 1.8 8us 0.1ns 0.1ns 8us 16us)
V35 Din3[4] 0 pulse(0 1.8 16us 0.1ns 0.1ns 16us 32us)
V36 Din3[5] 0 pulse(0 1.8 32us 0.1ns 0.1ns 32us 64us)
V37 Din3[6] 0 pulse(0 1.8 64us 0.1ns 0.1ns 64us 128us)
V38 Din3[7] 0 pulse(0 1.8 128us 0.1ns 0.1ns 128us 256us)

.tran 5u 10u
.control
run
set xbrushwidth=2
set hcopydevtype = svg
plot VOUT0 VOUT1 VOUT2 VOUT3
hardcopy dac_top.svg VOUT0 VOUT1 VOUT2 VOUT3
.endc
.end
