VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO dac_top
  CLASS BLOCK ;
  FOREIGN dac_top ;
  ORIGIN 2.500 2.500 ;
  SIZE 217.500 BY 434.450 ;
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.450 212.020 6.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 11.590 212.020 12.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 17.730 212.020 18.430 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 23.870 212.020 24.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 30.010 212.020 30.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 36.150 212.020 36.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 42.290 212.020 42.990 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 48.430 212.020 49.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 54.570 212.020 55.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 60.710 212.020 61.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 66.850 212.020 67.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 72.990 212.020 73.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 79.130 212.020 79.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 85.270 212.020 85.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 91.410 212.020 92.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 97.550 212.020 98.250 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 103.690 212.020 104.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 109.830 212.020 110.530 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 115.970 212.020 116.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 122.110 212.020 122.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 128.250 212.020 128.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 134.390 212.020 135.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 140.530 212.020 141.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 146.670 212.020 147.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 152.810 212.020 153.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 158.950 212.020 159.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 165.090 212.020 165.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 171.230 212.020 171.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 177.370 212.020 178.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 183.510 212.020 184.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 189.650 212.020 190.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 195.790 212.020 196.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 201.930 212.020 202.630 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 208.070 212.020 208.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 214.210 212.020 214.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 220.350 212.020 221.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 226.490 212.020 227.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 232.630 212.020 233.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 238.770 212.020 239.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 244.910 212.020 245.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 251.050 212.020 251.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 257.190 212.020 257.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 263.330 212.020 264.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 269.470 212.020 270.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 275.610 212.020 276.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 281.750 212.020 282.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 287.890 212.020 288.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 294.030 212.020 294.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 300.170 212.020 300.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 306.310 212.020 307.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 312.450 212.020 313.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 318.590 212.020 319.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 324.730 212.020 325.430 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 330.870 212.020 331.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 337.010 212.020 337.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 343.150 212.020 343.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 349.290 212.020 349.990 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 355.430 212.020 356.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 361.570 212.020 362.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 367.710 212.020 368.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 373.850 212.020 374.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 379.990 212.020 380.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 386.130 212.020 386.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 392.270 212.020 392.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 404.470 212.020 404.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 426.945 212.020 427.445 ;
    END
  END VDDA
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.000 212.020 2.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 8.140 212.020 8.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 14.280 212.020 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 20.420 212.020 21.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 26.560 212.020 27.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 32.700 212.020 33.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 38.840 212.020 39.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 44.980 212.020 45.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 51.120 212.020 51.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 57.260 212.020 57.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 63.400 212.020 64.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 69.540 212.020 70.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 75.680 212.020 76.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 81.820 212.020 82.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 87.960 212.020 88.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 94.100 212.020 94.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 100.240 212.020 100.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 106.380 212.020 107.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 112.520 212.020 113.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 118.660 212.020 119.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 124.800 212.020 125.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 130.940 212.020 131.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 137.080 212.020 137.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 143.220 212.020 143.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 149.360 212.020 150.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 155.500 212.020 156.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 161.640 212.020 162.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 167.780 212.020 168.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 173.920 212.020 174.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 180.060 212.020 180.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 186.200 212.020 186.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 192.340 212.020 193.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 198.480 212.020 199.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 204.620 212.020 205.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 210.760 212.020 211.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 216.900 212.020 217.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 223.040 212.020 223.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 229.180 212.020 229.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 212.020 236.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 241.460 212.020 242.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 247.600 212.020 248.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 253.740 212.020 254.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 259.880 212.020 260.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 266.020 212.020 266.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 272.160 212.020 272.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 278.300 212.020 279.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 284.440 212.020 285.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 290.580 212.020 291.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 296.720 212.020 297.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 302.860 212.020 303.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 309.000 212.020 309.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 315.140 212.020 315.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 321.280 212.020 321.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 327.420 212.020 328.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 333.560 212.020 334.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 339.700 212.020 340.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 345.840 212.020 346.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 351.980 212.020 352.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 358.120 212.020 358.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 364.260 212.020 364.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 370.400 212.020 371.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 376.540 212.020 377.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 382.680 212.020 383.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 388.820 212.020 389.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 408.190 212.020 408.690 ;
    END
  END VSSA
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.000 400.635 212.020 401.135 ;
    END
  END VCCD
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.000 396.975 212.020 397.475 ;
    END
  END VSSD
  PIN VREFH
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -4.000 0.000 -0.030 0.700 ;
    END
  END VREFH
  PIN Din0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.725 405.755 3.895 434.000 ;
    END
  END Din0[0]
  PIN Din0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.240 405.395 4.410 434.000 ;
    END
  END Din0[1]
  PIN Din0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.730 405.715 4.900 434.000 ;
    END
  END Din0[2]
  PIN Din0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.250 406.035 5.420 434.000 ;
    END
  END Din0[3]
  PIN Din0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.790 406.355 5.960 434.000 ;
    END
  END Din0[4]
  PIN Din0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.290 406.675 6.460 434.000 ;
    END
  END Din0[5]
  PIN Din0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.830 406.995 7.000 434.000 ;
    END
  END Din0[6]
  PIN Din0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.390 407.315 7.560 434.000 ;
    END
  END Din0[7]
  PIN Din1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.730 405.755 56.900 434.000 ;
    END
  END Din1[0]
  PIN Din1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.245 405.395 57.415 434.000 ;
    END
  END Din1[1]
  PIN Din1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.735 405.715 57.905 434.000 ;
    END
  END Din1[2]
  PIN Din1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.255 406.035 58.425 434.000 ;
    END
  END Din1[3]
  PIN Din1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.795 406.355 58.965 434.000 ;
    END
  END Din1[4]
  PIN Din1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.295 406.675 59.465 434.000 ;
    END
  END Din1[5]
  PIN Din1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.835 406.995 60.005 434.000 ;
    END
  END Din1[6]
  PIN Din1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.395 407.315 60.565 434.000 ;
    END
  END Din1[7]
  PIN Din2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.735 405.755 109.905 434.000 ;
    END
  END Din2[0]
  PIN Din2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.250 405.395 110.420 434.000 ;
    END
  END Din2[1]
  PIN Din2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.740 405.715 110.910 434.000 ;
    END
  END Din2[2]
  PIN Din2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.260 406.035 111.430 434.000 ;
    END
  END Din2[3]
  PIN Din2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.800 406.355 111.970 434.000 ;
    END
  END Din2[4]
  PIN Din2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.300 406.675 112.470 434.000 ;
    END
  END Din2[5]
  PIN Din2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.840 406.995 113.010 434.000 ;
    END
  END Din2[6]
  PIN Din2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.400 407.315 113.570 434.000 ;
    END
  END Din2[7]
  PIN Din3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.740 405.755 162.910 434.000 ;
    END
  END Din3[0]
  PIN Din3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.255 405.395 163.425 434.000 ;
    END
  END Din3[1]
  PIN Din3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.745 405.715 163.915 434.000 ;
    END
  END Din3[2]
  PIN Din3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.265 406.035 164.435 434.000 ;
    END
  END Din3[3]
  PIN Din3[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.805 406.355 164.975 434.000 ;
    END
  END Din3[4]
  PIN Din3[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.305 406.675 165.475 434.000 ;
    END
  END Din3[5]
  PIN Din3[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.845 406.995 166.015 434.000 ;
    END
  END Din3[6]
  PIN Din3[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.405 407.315 166.575 434.000 ;
    END
  END Din3[7]
  PIN VOUT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.325 423.830 46.865 434.000 ;
    END
  END VOUT0
  PIN VOUT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.330 423.830 99.870 434.000 ;
    END
  END VOUT1
  PIN VOUT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.335 423.830 152.875 434.000 ;
    END
  END VOUT2
  PIN VOUT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.340 423.830 205.880 434.000 ;
    END
  END VOUT3
  OBS
      LAYER li1 ;
        RECT 0.000 0.000 212.020 427.735 ;
      LAYER met1 ;
        RECT -0.060 -0.060 207.290 427.745 ;
      LAYER met2 ;
        RECT -0.030 405.475 3.445 427.720 ;
        RECT 7.840 423.550 46.045 427.720 ;
        RECT 47.145 423.550 56.450 427.720 ;
        RECT 7.840 407.035 56.450 423.550 ;
        RECT 60.845 423.550 99.050 427.720 ;
        RECT 100.150 423.550 109.455 427.720 ;
        RECT 60.845 407.035 109.455 423.550 ;
        RECT 113.850 423.550 152.055 427.720 ;
        RECT 153.155 423.550 162.460 427.720 ;
        RECT 113.850 407.035 162.460 423.550 ;
        RECT 166.855 423.550 205.060 427.720 ;
        RECT 206.160 423.550 211.310 427.720 ;
        RECT 166.855 407.035 211.310 423.550 ;
        RECT 7.280 406.715 56.450 407.035 ;
        RECT 60.285 406.715 109.455 407.035 ;
        RECT 113.290 406.715 162.460 407.035 ;
        RECT 166.295 406.715 211.310 407.035 ;
        RECT 6.740 406.395 56.450 406.715 ;
        RECT 59.745 406.395 109.455 406.715 ;
        RECT 112.750 406.395 162.460 406.715 ;
        RECT 165.755 406.395 211.310 406.715 ;
        RECT 6.240 406.075 56.450 406.395 ;
        RECT 59.245 406.075 109.455 406.395 ;
        RECT 112.250 406.075 162.460 406.395 ;
        RECT 165.255 406.075 211.310 406.395 ;
        RECT 5.700 405.755 56.450 406.075 ;
        RECT 58.705 405.755 109.455 406.075 ;
        RECT 111.710 405.755 162.460 406.075 ;
        RECT 164.715 405.755 211.310 406.075 ;
        RECT 5.180 405.475 56.450 405.755 ;
        RECT 58.185 405.475 109.455 405.755 ;
        RECT 111.190 405.475 162.460 405.755 ;
        RECT -0.030 405.115 3.960 405.475 ;
        RECT 5.180 405.435 56.965 405.475 ;
        RECT 58.185 405.435 109.970 405.475 ;
        RECT 111.190 405.435 162.975 405.475 ;
        RECT 164.195 405.435 211.310 405.755 ;
        RECT 4.690 405.115 56.965 405.435 ;
        RECT 57.695 405.115 109.970 405.435 ;
        RECT 110.700 405.115 162.975 405.435 ;
        RECT 163.705 405.115 211.310 405.435 ;
        RECT -0.030 0.980 211.310 405.115 ;
        RECT 0.250 -0.060 211.310 0.980 ;
      LAYER met3 ;
        RECT 21.670 409.090 206.470 426.545 ;
        RECT 21.670 405.370 206.470 407.790 ;
        RECT 21.670 401.535 206.470 404.070 ;
        RECT 21.670 397.875 206.470 400.235 ;
        RECT 21.670 393.370 206.470 396.575 ;
        RECT 21.670 389.920 206.470 391.870 ;
        RECT 21.670 387.230 206.470 388.420 ;
        RECT 21.670 383.780 206.470 385.730 ;
        RECT 21.670 381.090 206.470 382.280 ;
        RECT 21.670 377.640 206.470 379.590 ;
        RECT 21.670 374.950 206.470 376.140 ;
        RECT 21.670 371.500 206.470 373.450 ;
        RECT 21.670 368.810 206.470 370.000 ;
        RECT 21.670 365.360 206.470 367.310 ;
        RECT 21.670 362.670 206.470 363.860 ;
        RECT 21.670 359.220 206.470 361.170 ;
        RECT 21.670 356.530 206.470 357.720 ;
        RECT 21.670 353.080 206.470 355.030 ;
        RECT 21.670 350.390 206.470 351.580 ;
        RECT 21.670 346.940 206.470 348.890 ;
        RECT 21.670 344.250 206.470 345.440 ;
        RECT 21.670 340.800 206.470 342.750 ;
        RECT 21.670 338.110 206.470 339.300 ;
        RECT 21.670 334.660 206.470 336.610 ;
        RECT 21.670 331.970 206.470 333.160 ;
        RECT 21.670 328.520 206.470 330.470 ;
        RECT 21.670 325.830 206.470 327.020 ;
        RECT 21.670 322.380 206.470 324.330 ;
        RECT 21.670 319.690 206.470 320.880 ;
        RECT 21.670 316.240 206.470 318.190 ;
        RECT 21.670 313.550 206.470 314.740 ;
        RECT 21.670 310.100 206.470 312.050 ;
        RECT 21.670 307.410 206.470 308.600 ;
        RECT 21.670 303.960 206.470 305.910 ;
        RECT 21.670 301.270 206.470 302.460 ;
        RECT 21.670 297.820 206.470 299.770 ;
        RECT 21.670 295.130 206.470 296.320 ;
        RECT 21.670 291.680 206.470 293.630 ;
        RECT 21.670 288.990 206.470 290.180 ;
        RECT 21.670 285.540 206.470 287.490 ;
        RECT 21.670 282.850 206.470 284.040 ;
        RECT 21.670 279.400 206.470 281.350 ;
        RECT 21.670 276.710 206.470 277.900 ;
        RECT 21.670 273.260 206.470 275.210 ;
        RECT 21.670 270.570 206.470 271.760 ;
        RECT 21.670 267.120 206.470 269.070 ;
        RECT 21.670 264.430 206.470 265.620 ;
        RECT 21.670 260.980 206.470 262.930 ;
        RECT 21.670 258.290 206.470 259.480 ;
        RECT 21.670 254.840 206.470 256.790 ;
        RECT 21.670 252.150 206.470 253.340 ;
        RECT 21.670 248.700 206.470 250.650 ;
        RECT 21.670 246.010 206.470 247.200 ;
        RECT 21.670 242.560 206.470 244.510 ;
        RECT 21.670 239.870 206.470 241.060 ;
        RECT 21.670 236.420 206.470 238.370 ;
        RECT 21.670 233.730 206.470 234.920 ;
        RECT 21.670 230.280 206.470 232.230 ;
        RECT 21.670 227.590 206.470 228.780 ;
        RECT 21.670 224.140 206.470 226.090 ;
        RECT 21.670 221.450 206.470 222.640 ;
        RECT 21.670 218.000 206.470 219.950 ;
        RECT 21.670 215.310 206.470 216.500 ;
        RECT 21.670 211.860 206.470 213.810 ;
        RECT 21.670 209.170 206.470 210.360 ;
        RECT 21.670 205.720 206.470 207.670 ;
        RECT 21.670 203.030 206.470 204.220 ;
        RECT 21.670 199.580 206.470 201.530 ;
        RECT 21.670 196.890 206.470 198.080 ;
        RECT 21.670 193.440 206.470 195.390 ;
        RECT 21.670 190.750 206.470 191.940 ;
        RECT 21.670 187.300 206.470 189.250 ;
        RECT 21.670 184.610 206.470 185.800 ;
        RECT 21.670 181.160 206.470 183.110 ;
        RECT 21.670 178.470 206.470 179.660 ;
        RECT 21.670 175.020 206.470 176.970 ;
        RECT 21.670 172.330 206.470 173.520 ;
        RECT 21.670 168.880 206.470 170.830 ;
        RECT 21.670 166.190 206.470 167.380 ;
        RECT 21.670 162.740 206.470 164.690 ;
        RECT 21.670 160.050 206.470 161.240 ;
        RECT 21.670 156.600 206.470 158.550 ;
        RECT 21.670 153.910 206.470 155.100 ;
        RECT 21.670 150.460 206.470 152.410 ;
        RECT 21.670 147.770 206.470 148.960 ;
        RECT 21.670 144.320 206.470 146.270 ;
        RECT 21.670 141.630 206.470 142.820 ;
        RECT 21.670 138.180 206.470 140.130 ;
        RECT 21.670 135.490 206.470 136.680 ;
        RECT 21.670 132.040 206.470 133.990 ;
        RECT 21.670 129.350 206.470 130.540 ;
        RECT 21.670 125.900 206.470 127.850 ;
        RECT 21.670 123.210 206.470 124.400 ;
        RECT 21.670 119.760 206.470 121.710 ;
        RECT 21.670 117.070 206.470 118.260 ;
        RECT 21.670 113.620 206.470 115.570 ;
        RECT 21.670 110.930 206.470 112.120 ;
        RECT 21.670 107.480 206.470 109.430 ;
        RECT 21.670 104.790 206.470 105.980 ;
        RECT 21.670 101.340 206.470 103.290 ;
        RECT 21.670 98.650 206.470 99.840 ;
        RECT 21.670 95.200 206.470 97.150 ;
        RECT 21.670 92.510 206.470 93.700 ;
        RECT 21.670 89.060 206.470 91.010 ;
        RECT 21.670 86.370 206.470 87.560 ;
        RECT 21.670 82.920 206.470 84.870 ;
        RECT 21.670 80.230 206.470 81.420 ;
        RECT 21.670 76.780 206.470 78.730 ;
        RECT 21.670 74.090 206.470 75.280 ;
        RECT 21.670 70.640 206.470 72.590 ;
        RECT 21.670 67.950 206.470 69.140 ;
        RECT 21.670 64.500 206.470 66.450 ;
        RECT 21.670 61.810 206.470 63.000 ;
        RECT 21.670 58.360 206.470 60.310 ;
        RECT 21.670 55.670 206.470 56.860 ;
        RECT 21.670 52.220 206.470 54.170 ;
        RECT 21.670 49.530 206.470 50.720 ;
        RECT 21.670 46.080 206.470 48.030 ;
        RECT 21.670 43.390 206.470 44.580 ;
        RECT 21.670 39.940 206.470 41.890 ;
        RECT 21.670 37.250 206.470 38.440 ;
        RECT 21.670 33.800 206.470 35.750 ;
        RECT 21.670 31.110 206.470 32.300 ;
        RECT 21.670 27.660 206.470 29.610 ;
        RECT 21.670 24.970 206.470 26.160 ;
        RECT 21.670 21.520 206.470 23.470 ;
        RECT 21.670 18.830 206.470 20.020 ;
        RECT 21.670 15.380 206.470 17.330 ;
        RECT 21.670 12.690 206.470 13.880 ;
        RECT 21.670 9.240 206.470 11.190 ;
        RECT 21.670 6.550 206.470 7.740 ;
        RECT 21.670 3.100 206.470 5.050 ;
  END
END dac_top
END LIBRARY

