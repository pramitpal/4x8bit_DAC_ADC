** sch_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/z_stuff/All_schematic/dac_top.sch
.subckt dac_top Din0[0] Din0[1] Din0[2] Din0[3] Din0[4] Din0[5] Din0[6] Din0[7] Din1[0] Din1[1]
+ Din1[2] Din1[3] Din1[4] Din1[5] Din1[6] Din1[7] Din2[0] Din2[1] Din2[2] Din2[3] Din2[4] Din2[5] Din2[6]
+ Din2[7] Din3[0] Din3[1] Din3[2] Din3[3] Din3[4] Din3[5] Din3[6] Din3[7] VREFH VDDA VSSA VCCD VSSD VOUT0
+ VOUT1 VOUT2 VOUT3
*.PININFO Din0[0]:I Din0[1]:I Din0[2]:I Din0[3]:I Din0[4]:I Din0[5]:I Din0[6]:I Din0[7]:I Din1[0]:I
*+ Din1[1]:I Din1[2]:I Din1[3]:I Din1[4]:I Din1[5]:I Din1[6]:I Din1[7]:I Din2[0]:I Din2[1]:I Din2[2]:I Din2[3]:I
*+ Din2[4]:I Din2[5]:I Din2[6]:I Din2[7]:I Din3[0]:I Din3[1]:I Din3[2]:I Din3[3]:I Din3[4]:I Din3[5]:I Din3[6]:I
*+ Din3[7]:I VREFH:I VDDA:B VSSA:B VCCD:B VSSD:B VOUT0:O VOUT1:O VOUT2:O VOUT3:O
x1 VREFH VDDA Din0[0] VSSA Din0[1] VCCD Din0[2] VSSD Din0[3] VOUT0 Din0[4] Din0[5] Din0[6] Din0[7]
+ Din1[0] Din1[1] Din1[2] Din1[3] VOUT1 Din1[4] Din1[5] Din1[6] Din1[7] Din2[0] Din2[1] Din2[2] Din2[3]
+ Din2[4] VOUT2 Din2[5] Din2[6] Din2[7] Din3[0] Din3[1] Din3[2] Din3[3] VOUT3 Din3[4] Din3[5] Din3[6] Din3[7]
+ 4x8_bit_dac
.ends

* expanding   symbol:
*+  /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/z_stuff/All_schematic/4x8_bit_dac.sym # of pins=41
** sym_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/z_stuff/All_schematic/4x8_bit_dac.sym
** sch_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/z_stuff/All_schematic/4x8_bit_dac.sch
.subckt 4x8_bit_dac VREFH VDDA Din0[0] VSSA Din0[1] VCCD Din0[2] VSSD Din0[3] VOUT0 Din0[4] Din0[5]
+ Din0[6] Din0[7] Din1[0] Din1[1] Din1[2] Din1[3] VOUT1 Din1[4] Din1[5] Din1[6] Din1[7] Din2[0] Din2[1]
+ Din2[2] Din2[3] Din2[4] VOUT2 Din2[5] Din2[6] Din2[7] Din3[0] Din3[1] Din3[2] Din3[3] VOUT3 Din3[4] Din3[5]
+ Din3[6] Din3[7]
*.PININFO VREFH:I VOUT0:O VDDA:B Din0[0]:I Din0[1]:I Din0[2]:I Din0[3]:I Din0[4]:I Din0[5]:I
*+ Din0[6]:I Din0[7]:I Din1[0]:I Din1[1]:I Din1[2]:I Din1[3]:I Din1[4]:I Din1[5]:I Din1[6]:I Din1[7]:I Din2[0]:I
*+ Din2[1]:I Din2[2]:I Din2[3]:I Din2[4]:I Din2[5]:I Din2[6]:I Din2[7]:I Din3[0]:I Din3[1]:I Din3[2]:I Din3[3]:I
*+ Din3[4]:I Din3[5]:I Din3[6]:I Din3[7]:I VOUT1:O VOUT2:O VOUT3:O VSSA:B VCCD:B VSSD:B
x1 Din0[0] VREFH VCCD Din0[1] VSSD Din0[2] Din0[3] Din0[4] VDDA Din0[5] VSSA Din0[6] Din0[7] net1
+ VOUT0 8_bit_dac_tx_buffer
x2 Din1[0] VREFH VCCD Din1[1] VSSD Din1[2] Din1[3] Din1[4] VDDA Din1[5] VSSA Din1[6] Din1[7] net2
+ VOUT1 8_bit_dac_tx_buffer
x3 Din2[0] VREFH VCCD Din2[1] VSSD Din2[2] Din2[3] Din2[4] VDDA Din2[5] VSSA Din2[6] Din2[7] net3
+ VOUT2 8_bit_dac_tx_buffer
x4 Din3[0] VREFH VCCD Din3[1] VSSD Din3[2] Din3[3] Din3[4] VDDA Din3[5] VSSA Din3[6] Din3[7] net4
+ VOUT3 8_bit_dac_tx_buffer
.ends


* expanding   symbol:
*+  /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/z_stuff/All_schematic/8_bit_dac_tx_buffer.sym # of pins=15
** sym_path:
*+ /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/z_stuff/All_schematic/8_bit_dac_tx_buffer.sym
** sch_path:
*+ /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/z_stuff/All_schematic/8_bit_dac_tx_buffer.sch
.subckt 8_bit_dac_tx_buffer D0 VREFH VCCD D1 VSSD D2 D3 D4 VDDA D5 VSSA D6 D7 VOUT VOUT_BUF
*.PININFO VSSD:B VCCD:B VDDA:B VSSA:B VOUT_BUF:O D0:I D1:I D2:I D3:I D4:I D5:I D6:I D7:I VREFH:I
*+ VOUT:O
x1 VDDA VREFH VSSA net9 net10 net11 net12 net13 net14 net15 net8 net16 VOUT net1 net2 net3 net4 net5
+ net6 net7 VSSA 8_bit_dac
x2 VDDA VSSA VOUT VOUT_BUF opamp
x3 VSSD VCCD VDDA D0 D4 net5 net1 D1 D5 net6 net2 D2 D6 net3 net7 D7 D3 net8 net4 level_tx_8bit
.ends


* expanding   symbol:  8_bit_dac.sym # of pins=21
** sym_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/z_stuff/All_schematic/8_bit_dac.sym
** sch_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/z_stuff/All_schematic/8_bit_dac.sch
.subckt 8_bit_dac VCC VREFH VSS D0_BUF D1_BUF D2_BUF D3_BUF D4_BUF D5_BUF D6_BUF D7 D7_BUF VOUT D0
+ D1 D2 D3 D4 D5 D6 VREFL
*.PININFO D0:I D1:I D2:I D7:I VREFH:I VREFL:I D0_BUF:O D1_BUF:O D2_BUF:O D7_BUF:O VOUT:O VCC:B VSS:B
*+ D3:I D3_BUF:O D4:I D4_BUF:O D5:I D5_BUF:O D6_BUF:O D6:I
x1 VCC VREFH VSS D0_BUF D1_BUF D2_BUF D3_BUF D4_BUF D5_BUF BUF6 D6_BUF VINH BUF0 BUF1 BUF2 BUF3 BUF4
+ BUF5 VINT 7_bit_dac
x2 VCC VINT VSS BUF0 BUF1 BUF2 BUF3 BUF4 BUF5 D6 BUF6 VINL D0 D1 D2 D3 D4 D5 VREFL 7_bit_dac
x3 VCC D7 D7_BUF VSS VINH VOUT VINL switch_n_3v3
.ends


* expanding   symbol:  opamp.sym # of pins=4
** sym_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/z_stuff/All_schematic/opamp.sym
** sch_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/z_stuff/All_schematic/opamp.sch
.subckt opamp VDDA VSSA VIN VOUT
*.PININFO VOUT:O VIN:I VSSA:B VDDA:B
XM1 net1 net1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=8 nf=1 m=1
XM2 net2 net1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=8 nf=1 m=1
XM3 net2 net2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM4 net3 net1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=1
XM5 net6 VOUT net3 VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=1
XM6 net5 VIN net3 VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=1
XM7 out net4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=8 nf=1 m=1
XM8 net4 net4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=8 nf=1 m=1
XM9 net4 Vb1 net6 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM10 out Vb1 net5 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM11 net6 net2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM12 net5 net2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM13 net7 net1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=1
XM14 net8 net1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=1
XM17 net9 net9 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM18 out2 net9 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM15 out2 Vb1 net7 VDDA sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM16 net9 Vb1 net8 VDDA sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM19 net10 net2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=1 W=4 nf=1 m=1
XM20 net8 VOUT net10 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=1
XM21 net7 VIN net10 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=1
XM22 VOUT out VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=50 nf=1 m=1
XM23 VOUT out2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 nf=1 m=1
XR3 VSSA net1 VSSA sky130_fd_pr__res_generic_nd__hv W=1 L=1 mult=1 m=1
XR1 Vb1 VDDA VSSA sky130_fd_pr__res_generic_nd__hv W=1 L=1 mult=1 m=1
XR2 VSSA Vb1 VSSA sky130_fd_pr__res_generic_nd__hv W=1 L=1 mult=1 m=1
XM24 VOUT out VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=50 nf=1 m=1
XM25 VOUT out2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 nf=1 m=1
XM26 VOUT out VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=50 nf=1 m=1
XM27 VOUT out2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 nf=1 m=1
XM28 VOUT out VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=50 nf=1 m=1
XM29 VOUT out2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 nf=1 m=1
.ends


* expanding   symbol:  level_tx_8bit.sym # of pins=19
** sym_path:
*+ /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/z_stuff/All_schematic/level_tx_8bit.sym
** sch_path:
*+ /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/z_stuff/All_schematic/level_tx_8bit.sch
.subckt level_tx_8bit VSSD VCCD VDDA VIN0 VIN4 VOUT4 VOUT0 VIN1 VIN5 VOUT5 VOUT1 VIN2 VIN6 VOUT2
+ VOUT6 VIN7 VIN3 VOUT7 VOUT3
*.PININFO VDDA:B VCCD:B VSSD:B VIN0:I VOUT0:O VIN1:I VOUT1:O VIN2:I VOUT2:O VIN3:I VOUT3:O VIN4:I
*+ VOUT4:O VIN5:I VOUT5:O VIN6:I VOUT6:O VIN7:I VOUT7:O
x1 VDDA VOUT0 VCCD VIN0 VSSD level_tx_1bit
x2 VDDA VOUT1 VCCD VIN1 VSSD level_tx_1bit
x3 VDDA VOUT2 VCCD VIN2 VSSD level_tx_1bit
x4 VDDA VOUT3 VCCD VIN3 VSSD level_tx_1bit
x5 VDDA VOUT4 VCCD VIN4 VSSD level_tx_1bit
x6 VDDA VOUT5 VCCD VIN5 VSSD level_tx_1bit
x7 VDDA VOUT6 VCCD VIN6 VSSD level_tx_1bit
x8 VDDA VOUT7 VCCD VIN7 VSSD level_tx_1bit
.ends


* expanding   symbol:  7_bit_dac.sym # of pins=19
** sym_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/z_stuff/All_schematic/7_bit_dac.sym
** sch_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/z_stuff/All_schematic/7_bit_dac.sch
.subckt 7_bit_dac VCC VREFH VSS D0_BUF D1_BUF D2_BUF D3_BUF D4_BUF D5_BUF D6 D6_BUF VOUT D0 D1 D2 D3
+ D4 D5 VREFL
*.PININFO D0:I D1:I D2:I D6:I VREFH:I VREFL:I D0_BUF:O D1_BUF:O D2_BUF:O D6_BUF:O VOUT:O VCC:B VSS:B
*+ D3:I D3_BUF:O D4:I D4_BUF:O D5:I D5_BUF:O
x1 VCC VREFH VSS D0_BUF D1_BUF D2_BUF D3_BUF D4_BUF BUF5 D5_BUF VINH BUF0 BUF1 BUF2 BUF3 BUF4 VINT
+ 6_bit_dac
x2 VCC VINT VSS BUF0 BUF1 BUF2 BUF3 BUF4 D5 BUF5 VINL D0 D1 D2 D3 D4 VREFL 6_bit_dac
x3 VCC D6 D6_BUF VSS VINH VOUT VINL switch_n_3v3
.ends


* expanding   symbol:  switch_n_3v3.sym # of pins=7
** sym_path:
*+ /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/z_stuff/All_schematic/switch_n_3v3.sym
** sch_path:
*+ /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/z_stuff/All_schematic/switch_n_3v3.sch
.subckt switch_n_3v3 VCC DX DX_BUF VSS VREFH VOUT VREFL
*.PININFO VCC:B VSS:B DX_BUF:O VOUT:O DX:I VREFH:I VREFL:I
XM1 net1 DX VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM2 net1 DX VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM3 DX_BUF net1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM4 DX_BUF net1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM5 VOUT net1 VREFL VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM6 VOUT net1 VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM7 VREFL DX_BUF VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM8 VREFH DX_BUF VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
.ends


* expanding   symbol:  level_tx_1bit.sym # of pins=5
** sym_path:
*+ /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/z_stuff/All_schematic/level_tx_1bit.sym
** sch_path:
*+ /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/z_stuff/All_schematic/level_tx_1bit.sch
.subckt level_tx_1bit VDDA VOUT VCCD VIN VSSD
*.PININFO VDDA:B VIN:I VOUT:O VCCD:B VSSD:B
XM4 net2 VOUT VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM5 net1 VIN VCCD VCCD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM6 net1 VIN VSSD VSSD sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM7 net2 VIN VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM8 VOUT net1 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM9 VOUT net2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
.ends


* expanding   symbol:  6_bit_dac.sym # of pins=17
** sym_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/z_stuff/All_schematic/6_bit_dac.sym
** sch_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/z_stuff/All_schematic/6_bit_dac.sch
.subckt 6_bit_dac VCC VREFH VSS D0_BUF D1_BUF D2_BUF D3_BUF D4_BUF D5 D5_BUF VOUT D0 D1 D2 D3 D4
+ VREFL
*.PININFO D0:I D1:I D2:I D5:I VREFH:I VREFL:I D0_BUF:O D1_BUF:O D2_BUF:O D5_BUF:O VOUT:O VCC:B VSS:B
*+ D3:I D3_BUF:O D4:I D4_BUF:O
X1 VCC VREFH VSS D0_BUF D1_BUF D2_BUF D3_BUF BUF4 D4_BUF VINH BUF0 BUF1 BUF2 BUF3 VINT 5_bit_dac
X2 VCC VINT VSS BUF0 BUF1 BUF2 BUF3 D4 BUF4 VINL D0 D1 D2 D3 VREFL 5_bit_dac
x3 VCC D5 D5_BUF VSS VINH VOUT VINL switch_n_3v3
.ends


* expanding   symbol:  5_bit_dac.sym # of pins=15
** sym_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/z_stuff/All_schematic/5_bit_dac.sym
** sch_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/z_stuff/All_schematic/5_bit_dac.sch
.subckt 5_bit_dac VCC VREFH VSS D0_BUF D1_BUF D2_BUF D3_BUF D4 D4_BUF VOUT D0 D1 D2 D3 VREFL
*.PININFO D0:I D1:I D2:I D4:I VREFH:I VREFL:I D0_BUF:O D1_BUF:O D2_BUF:O D4_BUF:O VOUT:O VCC:B VSS:B
*+ D3:I D3_BUF:O
X1 VCC VREFH VSS D0_BUF D1_BUF D2_BUF BUF3 D3_BUF VINH BUF0 BUF1 BUF2 VINT 4_bit_dac
X2 VCC VINT VSS BUF0 BUF1 BUF2 D3 BUF3 VINL D0 D1 D2 VREFL 4_bit_dac
x3 VCC D4 D4_BUF VSS VINH VOUT VINL switch_n_3v3
.ends


* expanding   symbol:  4_bit_dac.sym # of pins=13
** sym_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/z_stuff/All_schematic/4_bit_dac.sym
** sch_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/z_stuff/All_schematic/4_bit_dac.sch
.subckt 4_bit_dac VCC VREFH VSS D0_BUF D1_BUF D2_BUF D3 D3_BUF VOUT D0 D1 D2 VREFL
*.PININFO D0:I D1:I D2:I D3:I VREFH:I VREFL:I D0_BUF:O D1_BUF:O D2_BUF:O D3_BUF:O VOUT:O VCC:B VSS:B
X1 VCC VSS VREFH D0_BUF D1_BUF BUF2 D2_BUF VINH BUF0 BUF1 VINT 3_bit_dac
X2 VCC VSS VINT BUF0 BUF1 D2 BUF2 VINL D0 D1 VREFL 3_bit_dac
x3 VCC D3 D3_BUF VSS VINH VOUT VINL switch_n_3v3
.ends


* expanding   symbol:  3_bit_dac.sym # of pins=11
** sym_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/z_stuff/All_schematic/3_bit_dac.sym
** sch_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/z_stuff/All_schematic/3_bit_dac.sch
.subckt 3_bit_dac VCC VSS VREFH D0_BUF D1_BUF D2 D2_BUF VOUT D0 D1 VREFL
*.PININFO D2:I D0_BUF:O D2_BUF:O VOUT:O VREFH:I VCC:B VSS:B D1_BUF:O D1:I VREFL:I D0:I
x2 VCC D2 D2_BUF VSS VINH VOUT VINL switch_n_3v3
X1 VCC VSS BUF0 BUF1 VREFH D0_BUF D1_BUF VINT VINH 2_bit_dac
X3 VCC VSS D0 D1 VINT BUF0 BUF1 VREFL VINL 2_bit_dac
.ends


* expanding   symbol:  2_bit_dac.sym # of pins=9
** sym_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/z_stuff/All_schematic/2_bit_dac.sym
** sch_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/z_stuff/All_schematic/2_bit_dac.sch
.subckt 2_bit_dac VCC VSS D0 D1 VREFH D0_BUF D1_BUF VREFL VOUT
*.PININFO D1:I D0:I D0_BUF:O D1_BUF:O VOUT:O VREFL:I VREFH:I VCC:B VSS:B
x1 VCC D0_BUF D0 VREFH VSS VINL VINH VREFL switch2n_3v3
x2 VCC D1 D1_BUF VSS VINH VOUT VINL switch_n_3v3
.ends


* expanding   symbol:  switch2n_3v3.sym # of pins=8
** sym_path:
*+ /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/z_stuff/All_schematic/switch2n_3v3.sym
** sch_path:
*+ /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/z_stuff/All_schematic/switch2n_3v3.sch
.subckt switch2n_3v3 VCC DX_BUF DX VREFH VSS VOUTL VOUTH VREFL
*.PININFO VCC:B VSS:B VOUTL:O DX:I VOUTH:O DX_BUF:O VREFH:I VREFL:I
XM1 net1 DX VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM2 net1 DX VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM3 DX_BUF net1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM4 DX_BUF net1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM5 VOUTL net1 VREFL VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM6 VOUTL net1 net2 VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM7 VREFL DX_BUF VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM8 net2 DX_BUF VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM9 VOUTH net1 net3 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM10 VOUTH net1 net4 VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM11 net3 DX_BUF VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM12 net4 DX_BUF VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XR1 net3 net4 VSS sky130_fd_pr__res_generic_nd__hv W=1 L=1 mult=1 m=1
XR2 net2 net3 VSS sky130_fd_pr__res_generic_nd__hv W=1 L=1 mult=1 m=1
XR3 VREFL net2 VSS sky130_fd_pr__res_generic_nd__hv W=1 L=1 mult=1 m=1
XR4 net4 VREFH VSS sky130_fd_pr__res_generic_nd__hv W=1 L=1 mult=1 m=1
.ends

.end
