** sch_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/opamp/opamp.sch
.subckt opamp VOUT VIN VSSA VDDA
*.PININFO VOUT:O VIN:I VSSA:B VDDA:B
XM1 net1 net1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=8 nf=1 m=1
XM2 net2 net1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=8 nf=1 m=1
XM3 net2 net2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=1 m=1
XM4 net3 net1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 m=1
XM5 net6 VOUT net3 VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=1
XM6 net5 VIN net3 VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=1
XM7 out net4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=8 nf=1 m=1
XM8 net4 net4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=8 nf=1 m=1
XM9 net4 Vb1 net6 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM10 out Vb1 net5 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM11 net6 net2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM12 net5 net2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM13 net7 net1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=1
XM14 net8 net1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=1 W=4 nf=1 m=1
XM17 net9 net9 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM18 out2 net9 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM15 out2 Vb1 net7 VDDA sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM16 net9 Vb1 net8 VDDA sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM19 net10 net2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=1 W=4 nf=1 m=1
XM20 net8 VOUT net10 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=1
XM21 net7 VIN net10 VSSA sky130_fd_pr__nfet_g5v0d10v5 L=1 W=2 nf=1 m=1
XM22 VOUT out VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=50 nf=1 m=1
XM23 VOUT out2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 nf=1 m=1
XR3 VSSA net1 VSSA sky130_fd_pr__res_generic_nd__hv W=1 L=1 mult=1 m=1
XR1 Vb1 VDDA VSSA sky130_fd_pr__res_generic_nd__hv W=1 L=1 mult=1 m=1
XR2 VSSA Vb1 VSSA sky130_fd_pr__res_generic_nd__hv W=1 L=1 mult=1 m=1
XM24 VOUT out VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=50 nf=1 m=1
XM25 VOUT out2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 nf=1 m=1
XM26 VOUT out VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=50 nf=1 m=1
XM27 VOUT out2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 nf=1 m=1
XM28 VOUT out VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=50 nf=1 m=1
XM29 VOUT out2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 nf=1 m=1
.ends
.end
