magic
tech sky130A
magscale 1 2
timestamp 1686405580
<< locali >>
rect 5769 85181 5842 85343
rect -2409 78873 8192 78908
rect -2409 78768 460 78873
rect 600 78768 8192 78873
rect -2409 -65 8192 -40
rect -2409 -113 336 -65
rect 476 -113 8192 -65
rect -2409 -180 8192 -113
<< viali >>
rect 460 78768 600 78873
rect 336 -113 476 -65
<< metal1 >>
rect 5716 85415 7851 85508
rect 5716 85343 5809 85415
rect 5540 85181 5546 85343
rect 5708 85181 5842 85343
rect 6856 84586 6964 84592
rect 6856 83138 6964 84478
rect 6720 83030 6964 83138
rect 3143 82158 3222 82447
rect 3143 82073 3222 82079
rect 2145 81430 2151 81592
rect 2313 81430 2443 81592
rect 4086 81227 4179 81559
rect 4086 81134 7618 81227
rect 448 78873 612 78879
rect 448 78867 460 78873
rect 600 78867 612 78873
rect 448 78762 454 78867
rect 606 78762 612 78867
rect 454 78756 606 78762
rect 7525 77711 7618 81134
rect 7758 78385 7851 85415
rect 7752 78292 7758 78385
rect 7851 78292 7857 78385
rect 7519 77618 7525 77711
rect 7618 77618 7624 77711
rect 330 -59 482 -53
rect 324 -111 330 -59
rect 482 -111 488 -59
rect 324 -113 336 -111
rect 476 -113 488 -111
rect 324 -119 488 -113
<< via1 >>
rect 5546 85181 5708 85343
rect 6856 84478 6964 84586
rect 3143 82079 3222 82158
rect 2151 81430 2313 81592
rect 454 78768 460 78867
rect 460 78768 600 78867
rect 600 78768 606 78867
rect 454 78762 606 78768
rect 7758 78292 7851 78385
rect 7525 77618 7618 77711
rect 330 -65 482 -59
rect 330 -111 336 -65
rect 336 -111 476 -65
rect 476 -111 482 -65
<< metal2 >>
rect -1664 81005 -1630 85648
rect -2118 80971 -1630 81005
rect -2118 80869 -2084 80971
rect -1561 80933 -1527 85648
rect -1463 80997 -1429 85648
rect -1359 81061 -1325 85648
rect -1251 81125 -1217 85648
rect -1151 81189 -1117 85648
rect -1043 81253 -1009 85648
rect -931 81317 -897 85648
rect 5546 85343 5708 85349
rect 5537 85181 5546 85343
rect 5708 85181 5717 85343
rect 5546 85175 5708 85181
rect 6856 84586 6964 85648
rect 6850 84478 6856 84586
rect 6964 84478 6970 84586
rect 3137 82079 3143 82158
rect 3222 82079 3228 82158
rect 3143 82000 3222 82079
rect 6847 82000 8050 82001
rect 3143 81922 8050 82000
rect 3143 81921 6847 81922
rect 2151 81592 2313 81598
rect 2142 81430 2151 81592
rect 2313 81430 2322 81592
rect 2151 81424 2313 81430
rect -931 81283 6029 81317
rect -1043 81219 4870 81253
rect -1151 81155 3711 81189
rect -1251 81091 2552 81125
rect -1359 81027 1393 81061
rect -1463 80963 234 80997
rect -1561 80899 -925 80933
rect -959 80869 -925 80899
rect 200 80869 234 80963
rect 1359 80869 1393 81027
rect 2518 80869 2552 81091
rect 3677 80869 3711 81155
rect 4836 80867 4870 81219
rect 5995 80869 6029 81283
rect -2251 80725 -2242 80793
rect -2174 80725 -2165 80793
rect -2242 78676 -2174 80725
rect -2038 79224 -1920 79310
rect -1107 78807 -1052 79427
rect 52 78960 93 79154
rect 52 78919 821 78960
rect -1107 78752 329 78807
rect 448 78762 454 78867
rect 606 78762 612 78867
rect -2242 78608 109 78676
rect 41 78260 109 78608
rect 274 78533 329 78752
rect 478 78599 583 78762
rect 780 78660 821 78919
rect 1212 78780 1253 79166
rect 2374 78880 2415 79176
rect 3533 78960 3574 79154
rect 4691 79040 4732 79152
rect 4691 78999 5403 79040
rect 3533 78919 5323 78960
rect 2374 78839 5243 78880
rect 1212 78739 5163 78780
rect 780 78619 3605 78660
rect 378 78537 583 78599
rect 3564 78551 3605 78619
rect 5122 78551 5163 78739
rect 5202 78551 5243 78839
rect 5282 78551 5323 78919
rect 5362 78551 5403 78999
rect 5849 78680 5890 79160
rect 5442 78639 5890 78680
rect 5442 78539 5483 78639
rect 7009 78592 7050 79160
rect 5522 78551 7050 78592
rect 7758 78385 7851 78391
rect 7749 78292 7758 78385
rect 7851 78292 7860 78385
rect 7758 78286 7851 78292
rect 7525 77711 7618 77717
rect 7516 77618 7525 77711
rect 7618 77618 7627 77711
rect 7525 77612 7618 77618
rect 144 77306 212 77500
rect 7971 40257 8050 81922
rect 7200 40213 8050 40257
rect 7193 40178 8050 40213
rect 378 -59 433 86
rect 324 -111 330 -59
rect 482 -111 488 -59
<< via2 >>
rect 5546 85181 5708 85343
rect 2151 81430 2313 81592
rect -2242 80725 -2174 80793
rect 7758 78292 7851 78385
rect 7525 77618 7618 77711
<< metal3 >>
rect 5541 85343 5713 85348
rect 5541 85309 5546 85343
rect -2409 85209 5546 85309
rect 5541 85181 5546 85209
rect 5708 85309 5713 85343
rect 5708 85209 8192 85309
rect 5708 85181 5713 85209
rect 5541 85176 5713 85181
rect 2146 81592 2318 81597
rect 2146 81558 2151 81592
rect -2409 81458 2151 81558
rect 2146 81430 2151 81458
rect 2313 81558 2318 81592
rect 2313 81458 8192 81558
rect 2313 81430 2318 81458
rect 2146 81425 2318 81430
rect -2409 80793 -2056 80814
rect -2409 80725 -2242 80793
rect -2174 80725 -2056 80793
rect -2409 80714 -2056 80725
rect 7019 80714 8192 80811
rect -2409 79947 -2056 80047
rect 7016 79947 8192 80047
rect -2409 79215 -2056 79315
rect 7016 79215 8192 79315
rect -2409 78274 187 78414
rect 6966 78385 8192 78414
rect 6966 78292 7758 78385
rect 7851 78292 8192 78385
rect 6966 78274 8192 78292
rect -2409 77584 0 77724
rect 6986 77711 8192 77724
rect 6986 77618 7525 77711
rect 7618 77618 8192 77711
rect 6986 77584 8192 77618
rect -2409 77046 0 77186
rect 7082 77046 8192 77186
rect -2409 76356 0 76496
rect 7082 76356 8192 76496
rect -2409 75818 0 75958
rect 7082 75818 8192 75958
rect -2409 75128 0 75268
rect 7082 75128 8192 75268
rect -2409 74590 0 74730
rect 7082 74590 8192 74730
rect -2409 73900 0 74040
rect 7082 73900 8192 74040
rect -2409 73362 0 73502
rect 7082 73362 8192 73502
rect -2409 72672 0 72812
rect 7082 72672 8192 72812
rect -2409 72134 0 72274
rect 7082 72134 8192 72274
rect -2409 71444 0 71584
rect 7082 71444 8192 71584
rect -2409 70906 0 71046
rect 7082 70906 8192 71046
rect -2409 70216 0 70356
rect 7082 70216 8192 70356
rect -2409 69678 0 69818
rect 7082 69678 8192 69818
rect -2409 68988 0 69128
rect 7082 68988 8192 69128
rect -2409 68450 0 68590
rect 7082 68450 8192 68590
rect -2409 67760 0 67900
rect 7082 67760 8192 67900
rect -2409 67222 0 67362
rect 7082 67222 8192 67362
rect -2409 66532 0 66672
rect 7082 66532 8192 66672
rect -2409 65994 0 66134
rect 7082 65994 8192 66134
rect -2409 65304 0 65444
rect 7082 65304 8192 65444
rect -2409 64766 0 64906
rect 7082 64766 8192 64906
rect -2409 64076 0 64216
rect 7082 64076 8192 64216
rect -2409 63538 0 63678
rect 7082 63538 8192 63678
rect -2409 62848 0 62988
rect 7082 62848 8192 62988
rect -2409 62310 0 62450
rect 7082 62310 8192 62450
rect -2409 61620 0 61760
rect 7082 61620 8192 61760
rect -2409 61082 0 61222
rect 7082 61082 8192 61222
rect -2409 60392 0 60532
rect 7082 60392 8192 60532
rect -2409 59854 0 59994
rect 7082 59854 8192 59994
rect -2409 59164 0 59304
rect 7082 59164 8192 59304
rect -2409 58626 0 58766
rect 7082 58626 8192 58766
rect -2409 57936 0 58076
rect 7082 57936 8192 58076
rect -2409 57398 0 57538
rect 7082 57398 8192 57538
rect -2409 56708 0 56848
rect 7082 56708 8192 56848
rect -2409 56170 0 56310
rect 7082 56170 8192 56310
rect -2409 55480 0 55620
rect 7082 55480 8192 55620
rect -2409 54942 0 55082
rect 7082 54942 8192 55082
rect -2409 54252 0 54392
rect 7082 54252 8192 54392
rect -2409 53714 0 53854
rect 7082 53714 8192 53854
rect -2409 53024 0 53164
rect 7082 53024 8192 53164
rect -2409 52486 0 52626
rect 7082 52486 8192 52626
rect -2409 51796 0 51936
rect 7082 51796 8192 51936
rect -2409 51258 0 51398
rect 7082 51258 8192 51398
rect -2409 50568 0 50708
rect 7082 50568 8192 50708
rect -2409 50030 0 50170
rect 7082 50030 8192 50170
rect -2409 49340 0 49480
rect 7082 49340 8192 49480
rect -2409 48802 0 48942
rect 7082 48802 8192 48942
rect -2409 48112 0 48252
rect 7082 48112 8192 48252
rect -2409 47574 0 47714
rect 7082 47574 8192 47714
rect -2409 46884 0 47024
rect 7082 46884 8192 47024
rect -2409 46346 0 46486
rect 7082 46346 8192 46486
rect -2409 45656 0 45796
rect 7082 45656 8192 45796
rect -2409 45118 0 45258
rect 7082 45118 8192 45258
rect -2409 44428 0 44568
rect 7082 44428 8192 44568
rect -2409 43890 0 44030
rect 7082 43890 8192 44030
rect -2409 43200 0 43340
rect 7082 43200 8192 43340
rect -2409 42662 0 42802
rect 7082 42662 8192 42802
rect -2409 41972 0 42112
rect 7082 41972 8192 42112
rect -2409 41434 0 41574
rect 7082 41434 8192 41574
rect -2409 40744 0 40884
rect 7082 40744 8192 40884
rect -2409 40206 0 40346
rect 7082 40206 8192 40346
rect -2409 39516 0 39656
rect 7082 39516 8192 39656
rect -2409 38978 0 39118
rect 7082 38978 8192 39118
rect -2409 38288 0 38428
rect 7082 38288 8192 38428
rect -2409 37750 0 37890
rect 7082 37750 8192 37890
rect -2409 37060 0 37200
rect 7082 37060 8192 37200
rect -2409 36522 0 36662
rect 7082 36522 8192 36662
rect -2409 35832 0 35972
rect 7082 35832 8192 35972
rect -2409 35294 0 35434
rect 7082 35294 8192 35434
rect -2409 34604 0 34744
rect 7082 34604 8192 34744
rect -2409 34066 0 34206
rect 7082 34066 8192 34206
rect -2409 33376 0 33516
rect 7082 33376 8192 33516
rect -2409 32838 0 32978
rect 7082 32838 8192 32978
rect -2409 32148 0 32288
rect 7082 32148 8192 32288
rect -2409 31610 0 31750
rect 7082 31610 8192 31750
rect -2409 30920 0 31060
rect 7082 30920 8192 31060
rect -2409 30382 0 30522
rect 7082 30382 8192 30522
rect -2409 29692 0 29832
rect 7082 29692 8192 29832
rect -2409 29154 0 29294
rect 7082 29154 8192 29294
rect -2409 28464 0 28604
rect 7082 28464 8192 28604
rect -2409 27926 0 28066
rect 7082 27926 8192 28066
rect -2409 27236 0 27376
rect 7082 27236 8192 27376
rect -2409 26698 0 26838
rect 7082 26698 8192 26838
rect -2409 26008 0 26148
rect 7082 26008 8192 26148
rect -2409 25470 0 25610
rect 7082 25470 8192 25610
rect -2409 24780 0 24920
rect 7082 24780 8192 24920
rect -2409 24242 0 24382
rect 7082 24242 8192 24382
rect -2409 23552 0 23692
rect 7082 23552 8192 23692
rect -2409 23014 0 23154
rect 7082 23014 8192 23154
rect -2409 22324 0 22464
rect 7082 22324 8192 22464
rect -2409 21786 0 21926
rect 7082 21786 8192 21926
rect -2409 21096 0 21236
rect 7082 21096 8192 21236
rect -2409 20558 0 20698
rect 7082 20558 8192 20698
rect -2409 19868 0 20008
rect 7082 19868 8192 20008
rect -2409 19330 0 19470
rect 7082 19330 8192 19470
rect -2409 18640 0 18780
rect 7082 18640 8192 18780
rect -2409 18102 0 18242
rect 7082 18102 8192 18242
rect -2409 17412 0 17552
rect 7082 17412 8192 17552
rect -2409 16874 0 17014
rect 7082 16874 8192 17014
rect -2409 16184 0 16324
rect 7082 16184 8192 16324
rect -2409 15646 0 15786
rect 7082 15646 8192 15786
rect -2409 14956 0 15096
rect 7082 14956 8192 15096
rect -2409 14418 0 14558
rect 7082 14418 8192 14558
rect -2409 13728 0 13868
rect 7082 13728 8192 13868
rect -2409 13190 0 13330
rect 7082 13190 8192 13330
rect -2409 12500 0 12640
rect 7082 12500 8192 12640
rect -2409 11962 0 12102
rect 7082 11962 8192 12102
rect -2409 11272 0 11412
rect 7082 11272 8192 11412
rect -2409 10734 0 10874
rect 7082 10734 8192 10874
rect -2409 10044 0 10184
rect 7082 10044 8192 10184
rect -2409 9506 0 9646
rect 7082 9506 8192 9646
rect -2409 8816 0 8956
rect 7082 8816 8192 8956
rect -2409 8278 0 8418
rect 7082 8278 8192 8418
rect -2409 7588 0 7728
rect 7082 7588 8192 7728
rect -2409 7050 0 7190
rect 7082 7050 8192 7190
rect -2409 6360 0 6500
rect 7082 6360 8192 6500
rect -2409 5822 0 5962
rect 7082 5822 8192 5962
rect -2409 5132 0 5272
rect 7082 5132 8192 5272
rect -2409 4594 0 4734
rect 7082 4594 8192 4734
rect -2409 3904 0 4044
rect 7082 3904 8192 4044
rect -2409 3366 0 3506
rect 7082 3366 8192 3506
rect -2409 2676 0 2816
rect 7082 2676 8192 2816
rect -2409 2138 0 2278
rect 7082 2138 8192 2278
rect -2409 1448 0 1588
rect 7082 1448 8192 1588
rect -2409 910 0 1050
rect 5037 910 8192 1050
rect -2409 220 0 360
rect 5076 220 8192 360
use 8_bit_dac  8_bit_dac_0
timestamp 1686024185
transform 1 0 0 0 1 0
box 0 0 8026 78592
use level_tx_8bit  level_tx_8bit_0
timestamp 1686240839
transform 1 0 -2156 0 1 79110
box 0 0 9272 1793
use opamp  opamp_0
timestamp 1686247030
transform 1 0 3066 0 1 81434
box -812 -4 3699 3985
<< labels >>
rlabel metal2 6008 80936 6008 80936 3 D7
rlabel metal2 4852 80953 4852 80953 3 D6
rlabel metal2 3691 80954 3691 80954 3 D5
rlabel metal2 2533 80939 2533 80939 3 D4
rlabel metal2 1379 80939 1379 80939 3 D3
rlabel metal2 222 80939 222 80939 3 D2
rlabel metal2 -2103 80938 -2103 80938 3 D0
rlabel metal2 -946 80916 -946 80916 3 D1
rlabel metal3 -2347 85262 -2347 85262 3 VDDA
rlabel metal3 -2374 79987 -2374 79987 3 VCCD
rlabel metal2 -1548 85638 -1548 85638 3 D1
rlabel metal2 -1446 85638 -1446 85638 3 D2
rlabel metal2 -1340 85633 -1340 85633 3 D3
rlabel metal2 -1235 85634 -1235 85634 3 D4
rlabel metal2 -1134 85633 -1134 85633 3 D5
rlabel metal2 -1022 85631 -1022 85631 3 D6
rlabel metal2 -912 85638 -912 85638 3 D7
rlabel metal2 6911 85596 6911 85596 3 VOUT
rlabel locali -2342 -117 -2342 -117 3 VREFH
rlabel locali -2339 78836 -2339 78836 3 VREFL
rlabel metal2 178 77378 178 77378 3 VSSA
flabel metal3 s -2360 79260 -2360 79260 7 FreeSans 800 0 0 0 VSSD
flabel metal2 s -1646 85632 -1646 85632 1 FreeSans 1600 0 0 0 D0
port 1 n signal input
<< end >>
