magic
tech sky130A
timestamp 1692509756
<< properties >>
string FIXED_BBOX -520 -520 520 520
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 10.00 l 10.00 val 207.6 carea 2.00 cperi 0.19 nx {} ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
