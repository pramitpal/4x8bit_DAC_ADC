.subckt dac_top DIN0 DIN1
.ends
