* NGSPICE file created from level_tx_1bit.ext - technology: sky130A

.subckt level_tx_1bit VIN VOUT VCCD VSSD VDDA
X0 a_n1423_1248# VOUT VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1 VSSD VIN a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.2
X2 VSSD VIN a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X3 VOUT a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4 a_n1353_675# VIN VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.2
X5 VOUT a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
.ends

