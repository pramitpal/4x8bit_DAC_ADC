magic
tech sky130A
magscale 1 2
timestamp 1688648239
<< metal1 >>
rect 0 -121 236 -21
<< metal2 >>
rect 642 84958 682 85090
rect 780 84928 820 85090
rect 916 84948 956 85090
rect 1050 84968 1090 85090
rect 1182 84952 1222 85090
rect 1314 84950 1354 85090
rect 1446 84954 1486 85090
rect 1580 84954 1620 85090
rect 6408 84928 6456 85090
rect 8368 84974 8408 85090
rect 8506 84974 8546 85090
rect 8642 84964 8682 85090
rect 8776 84986 8816 85090
rect 8908 84992 8948 85090
rect 9040 84988 9080 85090
rect 9172 84978 9212 85090
rect 9306 84980 9346 85090
rect 14134 84926 14182 85090
rect 16094 84998 16134 85090
rect 16232 84994 16272 85090
rect 16368 84974 16408 85090
rect 16502 84986 16542 85090
rect 16634 84990 16674 85090
rect 16766 84984 16806 85090
rect 16898 84992 16938 85090
rect 17032 84978 17072 85090
rect 21860 84952 21908 85090
rect 23820 85020 23860 85090
rect 23958 85014 23998 85090
rect 24094 85008 24134 85090
rect 24228 85014 24268 85090
rect 24360 85012 24400 85090
rect 24492 84994 24532 85090
rect 24624 85014 24664 85090
rect 24758 84996 24798 85090
rect 29586 84954 29634 85090
<< metal3 >>
rect 244 84602 792 84902
rect 56 81392 654 81692
rect 16 80262 254 80362
rect 0 79392 264 79492
rect 0 78932 228 79032
use 8_bit_dac_tx_buffer  8_bit_dac_tx_buffer_0
array 0 3 7726 0 0 85090
timestamp 1688642502
transform 1 0 0 0 1 0
box 0 -121 7726 85090
<< labels >>
flabel metal2 s 658 85056 658 85056 0 FreeSans 320 0 0 0 Din0[0]
flabel metal2 s 798 85058 798 85058 0 FreeSans 320 0 0 0 Din0[1]
flabel metal2 s 932 85058 932 85058 0 FreeSans 320 0 0 0 Din0[2]
flabel metal2 s 1070 85076 1070 85076 0 FreeSans 320 0 0 0 Din0[3]
flabel metal2 s 1198 85068 1198 85068 0 FreeSans 320 0 0 0 Din0[4]
flabel metal2 s 1342 85056 1342 85056 0 FreeSans 320 0 0 0 Din0[5]
flabel metal2 s 1472 85056 1472 85056 0 FreeSans 320 0 0 0 Din0[6]
flabel metal2 s 1598 85058 1598 85058 0 FreeSans 320 0 0 0 Din0[7]
flabel metal2 s 6430 85058 6430 85058 0 FreeSans 320 0 0 0 VOUT0
flabel metal2 s 8390 85064 8390 85064 0 FreeSans 320 0 0 0 Din1[0]
flabel metal2 s 8524 85064 8524 85064 0 FreeSans 320 0 0 0 Din1[1]
flabel metal2 s 8660 85070 8660 85070 0 FreeSans 320 0 0 0 Din1[2]
flabel metal2 s 8796 85076 8796 85076 0 FreeSans 320 0 0 0 Din1[3]
flabel metal2 s 8924 85062 8924 85062 0 FreeSans 320 0 0 0 Din1[4]
flabel metal2 s 9062 85068 9062 85068 0 FreeSans 320 0 0 0 Din1[5]
flabel metal2 s 9190 85064 9190 85064 0 FreeSans 320 0 0 0 Din1[6]
flabel metal2 s 9326 85076 9326 85076 0 FreeSans 320 0 0 0 Din1[7]
flabel metal2 s 14158 85064 14158 85064 0 FreeSans 320 0 0 0 VOUT1
flabel metal2 s 16116 85068 16116 85068 0 FreeSans 320 0 0 0 Din2[0]
flabel metal2 s 16250 85064 16250 85064 0 FreeSans 320 0 0 0 Din2[1]
flabel metal2 s 16388 85062 16388 85062 0 FreeSans 320 0 0 0 Din2[2]
flabel metal2 s 16524 85066 16524 85066 0 FreeSans 320 0 0 0 Din2[3]
flabel metal2 s 16654 85070 16654 85070 0 FreeSans 320 0 0 0 Din2[4]
flabel metal2 s 16784 85070 16784 85070 0 FreeSans 320 0 0 0 Din2[5]
flabel metal2 s 16924 85068 16924 85068 0 FreeSans 320 0 0 0 Din2[6]
flabel metal2 s 17056 85070 17056 85070 0 FreeSans 320 0 0 0 Din2[7]
flabel metal2 s 21888 85060 21888 85060 0 FreeSans 320 0 0 0 VOUT2
flabel metal2 s 23842 85074 23842 85074 0 FreeSans 320 0 0 0 Din3[0]
flabel metal2 s 23972 85074 23972 85074 0 FreeSans 320 0 0 0 Din3[1]
flabel metal2 s 24116 85066 24116 85066 0 FreeSans 320 0 0 0 Din3[2]
flabel metal2 s 24246 85064 24246 85064 0 FreeSans 320 0 0 0 Din3[3]
flabel metal2 s 24380 85068 24380 85068 0 FreeSans 320 0 0 0 Din3[4]
flabel metal2 s 24518 85074 24518 85074 0 FreeSans 320 0 0 0 Din3[5]
flabel metal2 s 24648 85066 24648 85066 0 FreeSans 320 0 0 0 Din3[6]
flabel metal2 s 24776 85070 24776 85070 0 FreeSans 320 0 0 0 Din3[7]
flabel metal2 s 29612 85062 29612 85062 0 FreeSans 320 0 0 0 VOUT3
flabel metal3 s 350 84762 350 84762 0 FreeSans 320 0 0 0 VDDA
flabel metal3 s 226 81540 226 81540 0 FreeSans 320 0 0 0 VSSA
flabel metal3 s 170 80316 170 80316 0 FreeSans 320 0 0 0 VDDA
flabel metal3 s 50 79440 50 79440 0 FreeSans 320 0 0 0 VSSD
flabel metal3 s 106 78986 106 78986 0 FreeSans 320 0 0 0 VCCD
flabel metal1 s 88 -66 88 -66 0 FreeSans 320 0 0 0 VREFH
<< end >>
