magic
tech sky130A
magscale 1 2
timestamp 1687539450
<< metal1 >>
rect 1138 77675 1182 77791
rect 1138 77631 1379 77675
rect 6968 40453 6974 40505
rect 7026 40453 7032 40505
rect 6808 40395 6814 40402
rect 6516 40356 6814 40395
rect 6808 40350 6814 40356
rect 6866 40350 6872 40402
rect 6985 40361 7015 40453
rect 5511 39865 5517 39917
rect 5569 39910 5575 39917
rect 5569 39903 5601 39910
rect 5569 39871 5628 39903
rect 5569 39865 5575 39871
rect 5510 39411 5516 39463
rect 5568 39456 5574 39463
rect 5568 39417 5594 39456
rect 5568 39411 5574 39417
rect 6908 39394 6936 39470
rect 6890 39342 6896 39394
rect 6948 39342 6954 39394
<< via1 >>
rect 6974 40453 7026 40505
rect 6814 40350 6866 40402
rect 5517 39865 5569 39917
rect 5516 39411 5568 39463
rect 6896 39342 6948 39394
<< metal2 >>
rect 274 78445 329 78592
rect 378 78447 433 78592
rect 3564 78478 3605 78592
rect 5122 78460 5163 78592
rect 5202 78460 5243 78592
rect 5282 78460 5323 78592
rect 5362 78460 5403 78592
rect 5442 78440 5483 78592
rect 5522 78460 5563 78592
rect 7421 60006 7521 60045
rect 6974 40505 7026 40511
rect 42 38810 110 40465
rect 5122 40407 5164 40480
rect 5202 40399 5244 40481
rect 5282 40401 5324 40483
rect 5362 40405 5404 40483
rect 5442 40411 5484 40483
rect 5522 40401 5564 40480
rect 7482 40494 7521 60006
rect 7026 40464 7521 40494
rect 6974 40447 7026 40453
rect 6814 40406 6866 40408
rect 6814 40402 7245 40406
rect 6866 40354 7245 40402
rect 6814 40344 6866 40350
rect 7193 40246 7245 40354
rect 7604 40246 7656 78470
rect 7193 40194 7656 40246
rect 5517 39917 5569 39923
rect 144 38148 212 39752
rect 5122 39707 5163 39861
rect 5202 39712 5243 39861
rect 5282 39703 5323 39861
rect 5362 39715 5403 39861
rect 5442 39715 5483 39861
rect 5517 39859 5569 39865
rect 5516 39463 5568 39469
rect 5516 39405 5568 39411
rect 6896 39394 6948 39400
rect 6948 39354 7523 39382
rect 6896 39336 6948 39342
rect 5122 39163 5164 39301
rect 5202 39165 5244 39285
rect 5282 39163 5324 39289
rect 5362 39141 5404 39287
rect 5442 39167 5484 39281
rect 5522 39171 5564 39295
rect 7484 20749 7523 39354
rect 7431 20710 7523 20749
rect 5122 1143 5163 1354
rect 5202 1141 5243 1363
rect 5282 1141 5323 1356
rect 5362 1141 5403 1356
rect 5442 1141 5483 1363
rect 5522 1141 5563 1364
rect 277 0 332 212
rect 378 0 433 224
rect 3564 0 3605 111
use 7_bit_dac  7_bit_dac_0
array 0 0 7470 0 1 39296
timestamp 1687539450
transform 1 0 0 0 1 0
box -2 0 7724 39296
use switch_n_3v3  switch_n_3v3_1
timestamp 1687539450
transform 1 0 12004 0 1 40200
box -6932 -990 -4922 236
<< labels >>
rlabel metal2 5138 78553 5138 78553 3 D2
rlabel metal2 5216 78558 5216 78558 3 D3
rlabel metal2 5305 78568 5305 78568 3 D4
rlabel metal2 5376 78572 5376 78572 3 D5
rlabel metal2 5468 78571 5468 78571 3 D6
rlabel metal2 5538 78578 5538 78578 3 D7
rlabel metal2 3591 78565 3591 78565 3 D1
rlabel metal2 290 78583 290 78583 3 D0
rlabel metal2 399 78576 399 78576 3 VREFL
rlabel metal2 297 52 297 52 3 D0_BUF
rlabel metal2 409 46 409 46 3 VREFH
rlabel metal2 3589 32 3589 32 3 D1_BUF
rlabel metal2 5137 1174 5137 1174 3 D2_BUF
rlabel metal2 5217 1169 5217 1169 3 D3_BUF
rlabel metal2 5295 1165 5295 1165 3 D4_BUF
rlabel metal2 5374 1161 5374 1161 3 D5_BUF
rlabel metal2 5449 1164 5449 1164 3 D6_BUF
rlabel metal2 5535 1161 5535 1161 3 D7_BUF
rlabel metal2 70 39257 70 39257 3 VCC
rlabel metal2 176 39252 176 39252 3 VSS
rlabel metal2 7578 40220 7578 40220 3 VOUT
flabel metal2 s 7626 78438 7626 78438 0 FreeSans 480 0 0 0 VOUT
<< end >>
