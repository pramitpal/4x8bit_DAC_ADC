magic
tech sky130A
magscale 1 2
timestamp 1692270715
<< metal3 >>
rect -3492 3172 -120 3200
rect -3492 148 -204 3172
rect -140 148 -120 3172
rect -3492 120 -120 148
rect 120 3172 3492 3200
rect 120 148 3408 3172
rect 3472 148 3492 3172
rect 120 120 3492 148
rect -3492 -148 -120 -120
rect -3492 -3172 -204 -148
rect -140 -3172 -120 -148
rect -3492 -3200 -120 -3172
rect 120 -148 3492 -120
rect 120 -3172 3408 -148
rect 3472 -3172 3492 -148
rect 120 -3200 3492 -3172
<< via3 >>
rect -204 148 -140 3172
rect 3408 148 3472 3172
rect -204 -3172 -140 -148
rect 3408 -3172 3472 -148
<< mimcap >>
rect -3452 3120 -452 3160
rect -3452 200 -3412 3120
rect -492 200 -452 3120
rect -3452 160 -452 200
rect 160 3120 3160 3160
rect 160 200 200 3120
rect 3120 200 3160 3120
rect 160 160 3160 200
rect -3452 -200 -452 -160
rect -3452 -3120 -3412 -200
rect -492 -3120 -452 -200
rect -3452 -3160 -452 -3120
rect 160 -200 3160 -160
rect 160 -3120 200 -200
rect 3120 -3120 3160 -200
rect 160 -3160 3160 -3120
<< mimcapcontact >>
rect -3412 200 -492 3120
rect 200 200 3120 3120
rect -3412 -3120 -492 -200
rect 200 -3120 3120 -200
<< metal4 >>
rect -2004 3121 -1900 3320
rect -224 3172 -120 3320
rect -3413 3120 -491 3121
rect -3413 200 -3412 3120
rect -492 200 -491 3120
rect -3413 199 -491 200
rect -2004 -199 -1900 199
rect -224 148 -204 3172
rect -140 148 -120 3172
rect 1608 3121 1712 3320
rect 3388 3172 3492 3320
rect 199 3120 3121 3121
rect 199 200 200 3120
rect 3120 200 3121 3120
rect 199 199 3121 200
rect -224 -148 -120 148
rect -3413 -200 -491 -199
rect -3413 -3120 -3412 -200
rect -492 -3120 -491 -200
rect -3413 -3121 -491 -3120
rect -2004 -3320 -1900 -3121
rect -224 -3172 -204 -148
rect -140 -3172 -120 -148
rect 1608 -199 1712 199
rect 3388 148 3408 3172
rect 3472 148 3492 3172
rect 3388 -148 3492 148
rect 199 -200 3121 -199
rect 199 -3120 200 -200
rect 3120 -3120 3121 -200
rect 199 -3121 3121 -3120
rect -224 -3320 -120 -3172
rect 1608 -3320 1712 -3121
rect 3388 -3172 3408 -148
rect 3472 -3172 3492 -148
rect 3388 -3320 3492 -3172
<< properties >>
string FIXED_BBOX 120 120 3200 3200
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 15.00 l 15.00 val 461.4 carea 2.00 cperi 0.19 nx 2 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
