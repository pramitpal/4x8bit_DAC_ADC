* NGSPICE file created from 5_bit_dac.ext - technology: sky130A

.subckt switch_n_3v3_v2 VREFH DX_BUF DX VCC VSS VOUT VREFL
X0 VOUT DX_BUF VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1 DX_ DX VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2 DX_BUF DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X3 VOUT DX_BUF VREFL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X4 DX_ DX VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5 VREFL DX_ VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6 DX_BUF DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7 VREFH DX_ VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt switch2n_3v3 VOUTH VOUTL DX_BUF DX VREFL VREFH VCC VSS
X0 VOUTH a_n6524_n498# a_n7536_n67# VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1 a_n7536_n67# DX_BUF VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2 a_n7536_n67# a_n7390_n590# VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3 DX_BUF a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4 VREFL DX_BUF VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X5 a_n7536_n67# VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6 a_n6524_n498# DX VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7 VOUTL a_n6524_n498# VREFL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8 VOUTH a_n6524_n498# a_n7390_n590# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9 a_n7390_n590# DX_BUF VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X10 a_n7390_n590# a_n7246_n584# VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X11 a_n7246_n584# VREFL VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X12 a_n7246_n584# DX_BUF VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X13 DX_BUF a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X14 a_n6524_n498# DX VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X15 VOUTL a_n6524_n498# a_n7246_n584# VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt x2_bit_dac VREFH D1_BUF D1 D0 VCC D0_BUF VOUT VREFL VSS
Xswitch_n_3v3_v2_0 switch2n_3v3_0/VOUTH D1_BUF D1 VCC VSS VOUT switch2n_3v3_0/VOUTL
+ switch_n_3v3_v2
Xswitch2n_3v3_0 switch2n_3v3_0/VOUTH switch2n_3v3_0/VOUTL D0_BUF D0 VREFL VREFH VCC
+ VSS switch2n_3v3
.ends

.subckt switch_n_3v3 VREFH DX_BUF m2_n6802_n990# m2_n6562_n990# D7 D6 D5 D4 DX m2_n6722_n990#
+ D3 D2 m2_n6482_n990# m2_n6882_n990# VCC VSS VOUT m2_n6642_n990# VREFL
X0 VOUT DX_BUF VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1 DX_ DX VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2 DX_BUF DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X3 VOUT DX_BUF VREFL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X4 DX_ DX VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5 VREFL DX_ VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6 DX_BUF DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7 VREFH DX_ VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt x3_bit_dac VREFH D1_BUF switch_n_3v3_1/D6 switch_n_3v3_1/D7 switch_n_3v3_1/D3
+ D2_BUF switch_n_3v3_1/D4 D2 D1 D0 D0_BUF VCC VOUT VREFL switch_n_3v3_1/D5 VSS
X2_bit_dac_0[0] VREFH D1_BUF 2_bit_dac_0[0]/D1 2_bit_dac_0[0]/D0 VCC D0_BUF 2_bit_dac_0[0]/VOUT
+ 2_bit_dac_0[1]/VREFH VSS x2_bit_dac
X2_bit_dac_0[1] 2_bit_dac_0[1]/VREFH 2_bit_dac_0[0]/D1 D1 D0 VCC 2_bit_dac_0[0]/D0
+ 2_bit_dac_0[1]/VOUT VREFL VSS x2_bit_dac
Xswitch_n_3v3_1 2_bit_dac_0[0]/VOUT D2_BUF switch_n_3v3_1/D3 switch_n_3v3_1/D6 switch_n_3v3_1/D7
+ switch_n_3v3_1/D6 switch_n_3v3_1/D5 switch_n_3v3_1/D4 D2 switch_n_3v3_1/D4 switch_n_3v3_1/D3
+ D2 switch_n_3v3_1/D7 D2_BUF VCC VSS VOUT switch_n_3v3_1/D5 2_bit_dac_0[1]/VOUT switch_n_3v3
.ends

.subckt x4_bit_dac VREFH D1_BUF D2_BUF D3 D2 switch_n_3v3_0/D7 D1 switch_n_3v3_0/D6
+ D0 switch_n_3v3_0/D5 switch_n_3v3_0/D4 D3_BUF D0_BUF VCC VOUT VREFL VSS
X3_bit_dac_0[0] VREFH D1_BUF switch_n_3v3_0/D6 switch_n_3v3_0/D7 D3_BUF D2_BUF switch_n_3v3_0/D4
+ switch_n_3v3_0/D2 3_bit_dac_0[0]/D1 3_bit_dac_0[0]/D0 D0_BUF VCC 3_bit_dac_0[0]/VOUT
+ 3_bit_dac_0[1]/VREFH switch_n_3v3_0/D5 VSS x3_bit_dac
X3_bit_dac_0[1] 3_bit_dac_0[1]/VREFH 3_bit_dac_0[0]/D1 switch_n_3v3_0/D6 switch_n_3v3_0/D7
+ D3 switch_n_3v3_0/D2 switch_n_3v3_0/D4 D2 D1 D0 3_bit_dac_0[0]/D0 VCC 3_bit_dac_0[1]/VOUT
+ VREFL switch_n_3v3_0/D5 VSS x3_bit_dac
Xswitch_n_3v3_0 3_bit_dac_0[0]/VOUT D3_BUF D3_BUF switch_n_3v3_0/D6 switch_n_3v3_0/D7
+ switch_n_3v3_0/D6 switch_n_3v3_0/D5 switch_n_3v3_0/D4 D3 switch_n_3v3_0/D4 D3 switch_n_3v3_0/D2
+ switch_n_3v3_0/D7 switch_n_3v3_0/D2 VCC VSS VOUT switch_n_3v3_0/D5 3_bit_dac_0[1]/VOUT
+ switch_n_3v3
.ends

.subckt x5_bit_dac VCC VSS D0 VREFL D0_BUF VREFH D1_BUF D1 D2 D3 D4 D2_BUF D3_BUF
+ D4_BUF VOUT
X4_bit_dac_0[0] VREFH D1_BUF D2_BUF switch_n_3v3_0/D3 switch_n_3v3_0/D2 switch_n_3v3_0/D7
+ 4_bit_dac_0[0]/D1 switch_n_3v3_0/D6 4_bit_dac_0[0]/D0 switch_n_3v3_0/D5 D4_BUF D3_BUF
+ D0_BUF VCC 4_bit_dac_0[0]/VOUT 4_bit_dac_0[1]/VREFH VSS x4_bit_dac
X4_bit_dac_0[1] 4_bit_dac_0[1]/VREFH 4_bit_dac_0[0]/D1 switch_n_3v3_0/D2 D3 D2 switch_n_3v3_0/D7
+ D1 switch_n_3v3_0/D6 D0 switch_n_3v3_0/D5 D4 switch_n_3v3_0/D3 4_bit_dac_0[0]/D0
+ VCC 4_bit_dac_0[1]/VOUT VREFL VSS x4_bit_dac
Xswitch_n_3v3_0 4_bit_dac_0[0]/VOUT D4_BUF switch_n_3v3_0/D3 switch_n_3v3_0/D6 switch_n_3v3_0/D7
+ switch_n_3v3_0/D6 switch_n_3v3_0/D5 D4 D4 D4_BUF switch_n_3v3_0/D3 switch_n_3v3_0/D2
+ switch_n_3v3_0/D7 switch_n_3v3_0/D2 VCC VSS VOUT switch_n_3v3_0/D5 4_bit_dac_0[1]/VOUT
+ switch_n_3v3
.ends

