* SPICE3 file created from 8_bit_dac_tx_buffer.ext - technology: sky130A

.subckt x8_bit_dac_tx_buffer VDDA VSSD VCCD VSSA D0 D1 D2 D3 D4 D5 D6 D7 VOUT VREFH
+ VOUT_BUF
X0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT 8_bit_dac_0/D5_BUF 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2 8_bit_dac_0/D5_BUF 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X3 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT 8_bit_dac_0/D5_BUF 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X4 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6 8_bit_dac_0/D5_BUF 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X8 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/D1_BUF 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X10 8_bit_dac_0/D1_BUF 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X11 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/D1_BUF 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X12 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X13 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X14 8_bit_dac_0/D1_BUF 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X15 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X16 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X17 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/D0_BUF 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X18 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X19 8_bit_dac_0/D0_BUF 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X20 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 8_bit_dac_0/D0_BUF 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X21 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X22 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X23 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X24 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X25 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/D0_BUF 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X26 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X27 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X28 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/D0_BUF 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X29 8_bit_dac_0/D0_BUF 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X30 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X31 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X32 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X33 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=126 ps=1.11k w=1 l=0.5
X34 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X35 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X36 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=63.2 ps=663 w=0.5 l=0.5
X37 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X38 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X39 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X40 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X41 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X42 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X43 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X44 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X45 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X46 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X47 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X48 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X49 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X50 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X51 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X52 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X53 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X54 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X55 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X56 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/D2_BUF 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X57 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X58 8_bit_dac_0/D2_BUF 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X59 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/D2_BUF 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X60 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X61 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X62 8_bit_dac_0/D2_BUF 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X63 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X64 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X65 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X66 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X67 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X68 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X69 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X70 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X71 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X72 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X73 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X74 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X75 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X76 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X77 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X78 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X79 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X80 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X81 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X82 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X83 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X84 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X85 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X86 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X87 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X88 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X89 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X90 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X91 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X92 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X93 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X94 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X95 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X96 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X97 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X98 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X99 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X100 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X101 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X102 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X103 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X104 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X105 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X106 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X107 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X108 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X109 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X110 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X111 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X112 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X113 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X114 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X115 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X116 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X117 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X118 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X119 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X120 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 8_bit_dac_0/D3_BUF 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X121 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X122 8_bit_dac_0/D3_BUF 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X123 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 8_bit_dac_0/D3_BUF 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X124 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X125 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X126 8_bit_dac_0/D3_BUF 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X127 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X128 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X129 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X130 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X131 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X132 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X133 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X134 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X135 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X136 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X137 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X138 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X139 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X140 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X141 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X142 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X143 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X144 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X145 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X146 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X147 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X148 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X149 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X150 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X151 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X152 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X153 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X154 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X155 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X156 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X157 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X158 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X159 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X160 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X161 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X162 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X163 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X164 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X165 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X166 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X167 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X168 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X169 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X170 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X171 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X172 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X173 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X174 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X175 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X176 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X177 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X178 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X179 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X180 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X181 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X182 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X183 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X184 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X185 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X186 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X187 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X188 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X189 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X190 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X191 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X192 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X193 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X194 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X195 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X196 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X197 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X198 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X199 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X200 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X201 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X202 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X203 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X204 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X205 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X206 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X207 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X208 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X209 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X210 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X211 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X212 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X213 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X214 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X215 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X216 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X217 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X218 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X219 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X220 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X221 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X222 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X223 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X224 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X225 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X226 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X227 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X228 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X229 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X230 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X231 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X232 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X233 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X234 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X235 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X236 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X237 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X238 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X239 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X240 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X241 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X242 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X243 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X244 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X245 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X246 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X247 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X248 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 8_bit_dac_0/D4_BUF 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X249 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X250 8_bit_dac_0/D4_BUF 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X251 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 8_bit_dac_0/D4_BUF 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X252 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X253 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X254 8_bit_dac_0/D4_BUF 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X255 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X256 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X257 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X258 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X259 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X260 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X261 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X262 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X263 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X264 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X265 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X266 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X267 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X268 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X269 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X270 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X271 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X272 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X273 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X274 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X275 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X276 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X277 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X278 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X279 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X280 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X281 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X282 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X283 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X284 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X285 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X286 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X287 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X288 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X289 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X290 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X291 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X292 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X293 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X294 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X295 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X296 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X297 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X298 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X299 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X300 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X301 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X302 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X303 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X304 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X305 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X306 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X307 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X308 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X309 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X310 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X311 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X312 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X313 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X314 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X315 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X316 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X317 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X318 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X319 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X320 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X321 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X322 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X323 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X324 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X325 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X326 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X327 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X328 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X329 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X330 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X331 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X332 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X333 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X334 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X335 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X336 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X337 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X338 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X339 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X340 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X341 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X342 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X343 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X344 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X345 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X346 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X347 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X348 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X349 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X350 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X351 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X352 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X353 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X354 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X355 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X356 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X357 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X358 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X359 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X360 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X361 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X362 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X363 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X364 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X365 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X366 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X367 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X368 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X369 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X370 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X371 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X372 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X373 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X374 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X375 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X376 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X377 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X378 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X379 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X380 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X381 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X382 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X383 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X384 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X385 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X386 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X387 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X388 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X389 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X390 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X391 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X392 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X393 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X394 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X395 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X396 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X397 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X398 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X399 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X400 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X401 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X402 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X403 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X404 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X405 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X406 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X407 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X408 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X409 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X410 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X411 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X412 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X413 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X414 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X415 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X416 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X417 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X418 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X419 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X420 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X421 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X422 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X423 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X424 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X425 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X426 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X427 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X428 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X429 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X430 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X431 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X432 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X433 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X434 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X435 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X436 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X437 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X438 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X439 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X440 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X441 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X442 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X443 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X444 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X445 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X446 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X447 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X448 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X449 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X450 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X451 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X452 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X453 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X454 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X455 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X456 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X457 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X458 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X459 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X460 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X461 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X462 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X463 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X464 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X465 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X466 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X467 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X468 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X469 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X470 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X471 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X472 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X473 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X474 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X475 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X476 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X477 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X478 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X479 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X480 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X481 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X482 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X483 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X484 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X485 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X486 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X487 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X488 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X489 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X490 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X491 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X492 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X493 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X494 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X495 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X496 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X497 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X498 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X499 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X500 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X501 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X502 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/switch_n_3v3_0/D4 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X503 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X504 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X505 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/switch_n_3v3_1/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X506 8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X507 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X508 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/switch_n_3v3_1/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X509 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X510 8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D5 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X511 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X512 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X513 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X514 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X515 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X516 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X517 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X518 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X519 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X520 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X521 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X522 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X523 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X524 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X525 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X526 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X527 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X528 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X529 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X530 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X531 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X532 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X533 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X534 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X535 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X536 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X537 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X538 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X539 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X540 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X541 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X542 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X543 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X544 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X545 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X546 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X547 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X548 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X549 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X550 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X551 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X552 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X553 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X554 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X555 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X556 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X557 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X558 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X559 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X560 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X561 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X562 8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X563 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X564 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X565 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X566 8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X567 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X568 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X569 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X570 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X571 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X572 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X573 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X574 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X575 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X576 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X577 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X578 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X579 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X580 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X581 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X582 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X583 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X584 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X585 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X586 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X587 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X588 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X589 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X590 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X591 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X592 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X593 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X594 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X595 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X596 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X597 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X598 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X599 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X600 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X601 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X602 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X603 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X604 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X605 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X606 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X607 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X608 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X609 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X610 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X611 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X612 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X613 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X614 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X615 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X616 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X617 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X618 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X619 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X620 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X621 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X622 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X623 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X624 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X625 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X626 8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X627 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X628 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X629 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X630 8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D3 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X631 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X632 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X633 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X634 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X635 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X636 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X637 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X638 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X639 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X640 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X641 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X642 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X643 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X644 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X645 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X646 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X647 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X648 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X649 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X650 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X651 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X652 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X653 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X654 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X655 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X656 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X657 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X658 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X659 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X660 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X661 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X662 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X663 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X664 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X665 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X666 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X667 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X668 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X669 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X670 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X671 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X672 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X673 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X674 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X675 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X676 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X677 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X678 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X679 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X680 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X681 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X682 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X683 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X684 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X685 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X686 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X687 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X688 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X689 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X690 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X691 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X692 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X693 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X694 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X695 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X696 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X697 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X698 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X699 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X700 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X701 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X702 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X703 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X704 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X705 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X706 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X707 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X708 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X709 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X710 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X711 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X712 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X713 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X714 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X715 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X716 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X717 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X718 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X719 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X720 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X721 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X722 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X723 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X724 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X725 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X726 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X727 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X728 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X729 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X730 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X731 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X732 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X733 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X734 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X735 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X736 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X737 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X738 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X739 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X740 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X741 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X742 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X743 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X744 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X745 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X746 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X747 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X748 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X749 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X750 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X751 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X752 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X753 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X754 8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X755 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X756 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X757 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X758 8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/D4 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X759 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X760 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X761 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X762 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X763 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X764 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X765 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X766 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X767 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X768 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X769 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X770 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X771 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X772 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X773 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X774 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X775 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X776 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X777 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X778 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X779 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X780 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X781 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X782 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X783 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X784 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X785 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X786 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X787 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X788 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X789 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X790 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X791 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X792 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X793 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X794 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X795 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X796 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X797 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X798 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X799 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X800 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X801 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X802 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X803 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X804 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X805 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X806 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X807 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X808 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X809 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X810 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X811 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X812 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X813 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X814 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X815 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X816 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X817 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X818 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X819 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X820 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X821 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X822 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X823 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X824 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X825 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X826 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X827 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X828 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X829 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X830 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X831 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X832 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X833 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X834 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X835 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X836 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X837 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X838 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X839 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X840 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X841 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X842 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X843 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X844 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X845 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X846 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X847 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X848 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X849 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X850 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X851 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X852 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X853 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X854 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X855 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X856 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X857 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X858 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X859 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X860 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X861 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X862 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X863 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X864 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X865 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X866 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X867 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X868 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X869 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X870 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X871 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X872 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X873 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X874 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X875 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X876 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X877 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X878 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X879 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X880 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X881 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X882 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X883 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X884 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X885 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X886 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X887 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X888 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X889 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X890 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X891 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X892 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X893 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X894 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X895 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X896 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X897 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X898 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X899 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X900 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X901 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X902 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X903 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X904 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X905 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X906 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X907 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X908 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X909 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X910 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X911 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X912 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X913 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X914 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X915 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X916 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X917 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X918 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X919 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X920 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X921 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X922 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X923 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X924 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X925 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X926 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X927 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X928 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X929 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X930 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X931 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X932 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X933 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X934 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X935 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X936 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X937 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X938 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X939 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X940 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X941 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X942 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X943 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X944 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X945 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X946 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X947 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X948 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X949 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X950 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X951 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X952 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X953 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X954 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X955 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X956 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X957 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X958 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X959 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X960 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X961 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X962 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X963 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X964 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X965 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X966 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X967 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X968 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X969 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X970 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X971 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X972 8_bit_dac_0/7_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X973 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X974 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X975 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X976 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X977 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X978 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X979 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X980 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X981 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X982 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X983 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X984 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X985 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/switch_n_3v3_1/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X986 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X987 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X988 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/switch_n_3v3_1/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X989 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X990 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X991 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X992 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X993 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/switch_n_3v3_1/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X994 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X995 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X996 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/switch_n_3v3_1/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X997 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X998 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X999 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1000 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1001 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/switch_n_3v3_1/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1002 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1003 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1004 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/switch_n_3v3_1/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1005 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1006 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/switch_n_3v3_0/D4 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1007 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1008 8_bit_dac_0/7_bit_dac_0[0]/VOUT 8_bit_dac_0/D6_BUF 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1009 8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/switch_n_3v3_1/D6 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1010 8_bit_dac_0/D6_BUF 8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1011 8_bit_dac_0/7_bit_dac_0[0]/VOUT 8_bit_dac_0/D6_BUF 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1012 8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/switch_n_3v3_1/D6 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1013 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1014 8_bit_dac_0/D6_BUF 8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1015 8_bit_dac_0/7_bit_dac_0[0]/6_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1016 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT 8_bit_dac_0/switch_n_3v3_1/D5 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1017 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1018 8_bit_dac_0/switch_n_3v3_1/D5 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1019 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT 8_bit_dac_0/switch_n_3v3_1/D5 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1020 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1021 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1022 8_bit_dac_0/switch_n_3v3_1/D5 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1023 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1024 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1025 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1026 8_bit_dac_0/7_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1027 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1028 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1029 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1030 8_bit_dac_0/7_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1031 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1032 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1033 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1034 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1035 8_bit_dac_0/7_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1036 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1037 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1038 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1039 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1040 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1041 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1042 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1043 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1044 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1045 8_bit_dac_0/7_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1046 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1047 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1048 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1049 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1050 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1051 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1052 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1053 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1054 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1055 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1056 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1057 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1058 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1059 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1060 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1061 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1062 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1063 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1064 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1065 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1066 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1067 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1068 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1069 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1070 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1071 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1072 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/switch_n_3v3_1/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1073 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1074 8_bit_dac_0/switch_n_3v3_1/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1075 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/switch_n_3v3_1/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1076 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1077 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1078 8_bit_dac_0/switch_n_3v3_1/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1079 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1080 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1081 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1082 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1083 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1084 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1085 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1086 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1087 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1088 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1089 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1090 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1091 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1092 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1093 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1094 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1095 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1096 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1097 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1098 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1099 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1100 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1101 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1102 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1103 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1104 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1105 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1106 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1107 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1108 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1109 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1110 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1111 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1112 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1113 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1114 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1115 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1116 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1117 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1118 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1119 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1120 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1121 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1122 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1123 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1124 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1125 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1126 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1127 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1128 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1129 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1130 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1131 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1132 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1133 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1134 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1135 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1136 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 8_bit_dac_0/switch_n_3v3_1/D3 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1137 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1138 8_bit_dac_0/switch_n_3v3_1/D3 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1139 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 8_bit_dac_0/switch_n_3v3_1/D3 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1140 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1141 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1142 8_bit_dac_0/switch_n_3v3_1/D3 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1143 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1144 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1145 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1146 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1147 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1148 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1149 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1150 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1151 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1152 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1153 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1154 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1155 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1156 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1157 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1158 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1159 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1160 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1161 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1162 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1163 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1164 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1165 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1166 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1167 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1168 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1169 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1170 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1171 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1172 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1173 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1174 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1175 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1176 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1177 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1178 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1179 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1180 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1181 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1182 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1183 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1184 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1185 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1186 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1187 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1188 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1189 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1190 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1191 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1192 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1193 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1194 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1195 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1196 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1197 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1198 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1199 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1200 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1201 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1202 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1203 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1204 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1205 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1206 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1207 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1208 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1209 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1210 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1211 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1212 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1213 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1214 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1215 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1216 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1217 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1218 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1219 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1220 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1221 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1222 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1223 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1224 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1225 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1226 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1227 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1228 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1229 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1230 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1231 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1232 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1233 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1234 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1235 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1236 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1237 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1238 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1239 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1240 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1241 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1242 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1243 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1244 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1245 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1246 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1247 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1248 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1249 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1250 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1251 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1252 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1253 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1254 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1255 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1256 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1257 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1258 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1259 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1260 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1261 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1262 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1263 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1264 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 8_bit_dac_0/switch_n_3v3_1/D4 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1265 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1266 8_bit_dac_0/switch_n_3v3_1/D4 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1267 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 8_bit_dac_0/switch_n_3v3_1/D4 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1268 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1269 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1270 8_bit_dac_0/switch_n_3v3_1/D4 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1271 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1272 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1273 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1274 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1275 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1276 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1277 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1278 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1279 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1280 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1281 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1282 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1283 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1284 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1285 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1286 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1287 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1288 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1289 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1290 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1291 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1292 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1293 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1294 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1295 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1296 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1297 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1298 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1299 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1300 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1301 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1302 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1303 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1304 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1305 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1306 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1307 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1308 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1309 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1310 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1311 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1312 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1313 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1314 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1315 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1316 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1317 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1318 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1319 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1320 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1321 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1322 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1323 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1324 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1325 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1326 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1327 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1328 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1329 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1330 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1331 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1332 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1333 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1334 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1335 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1336 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1337 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1338 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1339 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1340 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1341 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1342 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1343 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1344 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1345 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1346 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1347 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1348 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1349 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1350 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1351 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1352 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1353 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1354 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1355 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1356 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1357 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1358 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1359 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1360 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1361 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1362 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1363 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1364 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1365 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1366 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1367 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1368 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1369 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1370 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1371 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1372 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1373 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1374 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1375 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1376 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1377 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1378 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1379 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1380 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1381 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1382 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1383 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1384 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1385 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1386 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1387 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1388 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1389 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1390 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1391 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1392 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1393 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1394 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1395 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1396 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1397 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1398 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1399 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1400 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1401 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1402 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1403 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1404 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1405 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1406 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1407 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1408 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1409 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1410 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1411 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1412 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1413 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1414 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1415 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1416 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1417 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1418 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1419 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1420 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1421 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1422 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1423 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1424 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1425 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1426 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1427 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1428 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1429 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1430 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1431 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1432 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1433 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1434 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1435 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1436 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1437 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1438 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1439 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1440 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1441 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1442 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1443 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1444 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1445 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1446 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1447 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1448 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1449 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1450 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1451 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1452 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1453 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1454 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1455 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1456 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1457 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1458 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1459 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1460 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1461 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1462 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1463 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1464 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1465 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1466 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1467 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1468 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1469 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1470 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1471 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1472 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1473 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1474 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1475 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1476 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1477 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1478 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1479 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1480 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1481 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1482 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1483 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1484 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1485 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1486 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1487 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1488 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1489 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1490 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1491 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1492 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1493 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1494 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1495 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1496 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1497 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1498 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1499 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1500 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1501 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1502 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1503 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1504 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1505 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1506 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1507 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1508 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1509 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1510 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1511 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1512 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1513 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1514 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1515 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1516 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1517 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1518 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/switch_n_3v3_0/D4 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1519 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1520 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1521 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1522 8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1523 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1524 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/D5 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1525 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1526 8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D5 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1527 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1528 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1529 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1530 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1531 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1532 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1533 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1534 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1535 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1536 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1537 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1538 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1539 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1540 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1541 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1542 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1543 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1544 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1545 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1546 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1547 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1548 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1549 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1550 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1551 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1552 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1553 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1554 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1555 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1556 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1557 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1558 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1559 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1560 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1561 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1562 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1563 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1564 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1565 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1566 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1567 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1568 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1569 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1570 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1571 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1572 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1573 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1574 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1575 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1576 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1577 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1578 8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1579 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1580 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1581 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1582 8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1583 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1584 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1585 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1586 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1587 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1588 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1589 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1590 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1591 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1592 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1593 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1594 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1595 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1596 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1597 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1598 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1599 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1600 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1601 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1602 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1603 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1604 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1605 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1606 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1607 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1608 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1609 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1610 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1611 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1612 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1613 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1614 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1615 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1616 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1617 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1618 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1619 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1620 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1621 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1622 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1623 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1624 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1625 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1626 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1627 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1628 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1629 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1630 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1631 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1632 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1633 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1634 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1635 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1636 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1637 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1638 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1639 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1640 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1641 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1642 8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1643 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1644 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1645 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1646 8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D3 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1647 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1648 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1649 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1650 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1651 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1652 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1653 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1654 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1655 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1656 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1657 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1658 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1659 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1660 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1661 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1662 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1663 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1664 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1665 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1666 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1667 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1668 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1669 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1670 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1671 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1672 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1673 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1674 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1675 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1676 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1677 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1678 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1679 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1680 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1681 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1682 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1683 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1684 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1685 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1686 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1687 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1688 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1689 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1690 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1691 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1692 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1693 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1694 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1695 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1696 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1697 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1698 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1699 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1700 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1701 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1702 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1703 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1704 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1705 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1706 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1707 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1708 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1709 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1710 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1711 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1712 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1713 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1714 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1715 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1716 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1717 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1718 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1719 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1720 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1721 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1722 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1723 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1724 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1725 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1726 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1727 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1728 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1729 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1730 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1731 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1732 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1733 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1734 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1735 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1736 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1737 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1738 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1739 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1740 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1741 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1742 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1743 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1744 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1745 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1746 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1747 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1748 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1749 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1750 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1751 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1752 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1753 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1754 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1755 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1756 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1757 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1758 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1759 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1760 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1761 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1762 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1763 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1764 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1765 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1766 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1767 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1768 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1769 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1770 8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1771 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1772 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1773 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1774 8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/D4 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1775 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1776 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1777 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1778 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1779 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1780 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1781 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1782 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1783 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1784 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1785 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1786 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1787 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1788 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1789 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1790 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1791 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1792 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1793 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1794 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1795 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1796 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1797 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1798 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1799 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1800 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1801 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1802 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1803 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1804 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1805 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1806 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1807 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1808 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1809 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1810 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1811 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1812 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1813 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1814 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1815 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1816 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1817 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1818 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1819 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1820 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1821 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1822 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1823 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1824 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1825 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1826 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1827 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1828 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1829 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1830 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1831 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1832 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1833 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1834 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1835 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1836 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1837 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1838 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1839 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1840 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1841 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1842 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1843 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1844 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1845 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1846 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1847 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1848 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1849 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1850 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1851 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1852 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1853 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1854 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1855 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1856 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1857 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1858 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1859 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1860 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1861 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1862 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1863 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1864 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1865 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1866 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1867 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1868 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1869 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1870 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1871 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1872 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1873 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1874 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1875 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1876 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1877 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1878 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1879 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1880 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1881 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1882 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1883 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1884 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1885 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1886 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1887 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1888 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1889 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1890 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1891 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1892 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1893 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1894 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1895 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1896 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1897 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1898 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1899 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1900 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1901 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1902 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1903 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1904 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1905 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1906 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1907 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1908 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1909 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1910 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1911 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1912 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1913 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1914 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1915 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1916 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1917 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1918 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1919 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1920 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1921 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1922 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1923 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1924 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1925 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1926 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1927 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1928 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1929 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1930 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1931 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1932 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1933 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1934 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1935 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1936 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1937 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1938 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1939 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1940 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1941 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1942 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1943 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1944 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1945 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1946 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1947 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1948 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1949 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1950 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1951 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1952 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1953 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1954 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1955 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1956 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1957 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1958 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1959 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1960 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1961 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1962 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1963 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1964 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1965 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1966 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1967 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1968 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1969 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1970 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1971 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1972 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1973 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1974 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1975 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1976 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X1977 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1978 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1979 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X1980 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/D1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1981 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X1982 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1983 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X1984 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X1985 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1986 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1987 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1988 VSSA 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=23.8 pd=36.9 as=0 ps=0 w=1 l=0.5
X1989 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1990 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/D0 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1991 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1992 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X1993 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1994 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1995 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSSA VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1996 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X1997 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1998 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1999 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2000 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2001 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2002 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2003 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2004 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/D2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2005 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2006 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2007 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2008 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2009 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2010 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2011 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2012 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/D3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2013 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2014 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2015 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2016 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2017 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2018 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2019 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2020 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/D4 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2021 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2022 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/switch_n_3v3_0/D4 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2023 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2024 8_bit_dac_0/7_bit_dac_0[1]/VOUT 8_bit_dac_0/switch_n_3v3_1/D6 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X2025 8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/D6 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2026 8_bit_dac_0/switch_n_3v3_1/D6 8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2027 8_bit_dac_0/7_bit_dac_0[1]/VOUT 8_bit_dac_0/switch_n_3v3_1/D6 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X2028 8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/D6 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2029 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[1]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2030 8_bit_dac_0/switch_n_3v3_1/D6 8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2031 8_bit_dac_0/7_bit_dac_0[1]/6_bit_dac_0[0]/VOUT 8_bit_dac_0/7_bit_dac_0[1]/switch_n_3v3_1/DX_ 8_bit_dac_0/7_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2032 VOUT 8_bit_dac_0/D7_BUF 8_bit_dac_0/7_bit_dac_0[0]/VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=3.16 as=0 ps=0 w=0.5 l=0.5
X2033 8_bit_dac_0/switch_n_3v3_1/DX_ 8_bit_dac_0/D7 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2034 8_bit_dac_0/D7_BUF 8_bit_dac_0/switch_n_3v3_1/DX_ VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2035 VOUT 8_bit_dac_0/D7_BUF 8_bit_dac_0/7_bit_dac_0[1]/VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.5
X2036 8_bit_dac_0/switch_n_3v3_1/DX_ 8_bit_dac_0/D7 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2037 8_bit_dac_0/7_bit_dac_0[1]/VOUT 8_bit_dac_0/switch_n_3v3_1/DX_ VOUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X2038 8_bit_dac_0/D7_BUF 8_bit_dac_0/switch_n_3v3_1/DX_ VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2039 8_bit_dac_0/7_bit_dac_0[0]/VOUT 8_bit_dac_0/switch_n_3v3_1/DX_ VOUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X2040 level_tx_8bit_0/level_tx_1bit_0[0]/a_n1423_1248# 8_bit_dac_0/D0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2041 VSSD D0 level_tx_8bit_0/level_tx_1bit_0[0]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.2
X2042 VSSD D0 level_tx_8bit_0/level_tx_1bit_0[0]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X2043 8_bit_dac_0/D0 level_tx_8bit_0/level_tx_1bit_0[0]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2044 level_tx_8bit_0/level_tx_1bit_0[0]/a_n1353_675# D0 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.2
X2045 8_bit_dac_0/D0 level_tx_8bit_0/level_tx_1bit_0[0]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X2046 level_tx_8bit_0/level_tx_1bit_0[1]/a_n1423_1248# 8_bit_dac_0/D1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2047 VSSD D1 level_tx_8bit_0/level_tx_1bit_0[1]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0.974 pd=11.4 as=0.122 ps=1.42 w=0.42 l=0.2
X2048 VSSD D1 level_tx_8bit_0/level_tx_1bit_0[1]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=2.32 pd=20.6 as=0.29 ps=2.58 w=1 l=0.5
X2049 8_bit_dac_0/D1 level_tx_8bit_0/level_tx_1bit_0[1]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2050 level_tx_8bit_0/level_tx_1bit_0[1]/a_n1353_675# D1 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=1.16 ps=12.6 w=0.5 l=0.2
X2051 8_bit_dac_0/D1 level_tx_8bit_0/level_tx_1bit_0[1]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2052 level_tx_8bit_0/level_tx_1bit_0[2]/a_n1423_1248# 8_bit_dac_0/D2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2053 VSSD D2 level_tx_8bit_0/level_tx_1bit_0[2]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X2054 VSSD D2 level_tx_8bit_0/level_tx_1bit_0[2]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2055 8_bit_dac_0/D2 level_tx_8bit_0/level_tx_1bit_0[2]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2056 level_tx_8bit_0/level_tx_1bit_0[2]/a_n1353_675# D2 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X2057 8_bit_dac_0/D2 level_tx_8bit_0/level_tx_1bit_0[2]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2058 level_tx_8bit_0/level_tx_1bit_0[3]/a_n1423_1248# 8_bit_dac_0/D3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2059 VSSD D3 level_tx_8bit_0/level_tx_1bit_0[3]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X2060 VSSD D3 level_tx_8bit_0/level_tx_1bit_0[3]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2061 8_bit_dac_0/D3 level_tx_8bit_0/level_tx_1bit_0[3]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2062 level_tx_8bit_0/level_tx_1bit_0[3]/a_n1353_675# D3 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X2063 8_bit_dac_0/D3 level_tx_8bit_0/level_tx_1bit_0[3]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2064 level_tx_8bit_0/level_tx_1bit_0[4]/a_n1423_1248# 8_bit_dac_0/D4 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2065 VSSD D4 level_tx_8bit_0/level_tx_1bit_0[4]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X2066 VSSD D4 level_tx_8bit_0/level_tx_1bit_0[4]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2067 8_bit_dac_0/D4 level_tx_8bit_0/level_tx_1bit_0[4]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2068 level_tx_8bit_0/level_tx_1bit_0[4]/a_n1353_675# D4 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X2069 8_bit_dac_0/D4 level_tx_8bit_0/level_tx_1bit_0[4]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2070 level_tx_8bit_0/level_tx_1bit_0[5]/a_n1423_1248# 8_bit_dac_0/D5 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2071 VSSD D5 level_tx_8bit_0/level_tx_1bit_0[5]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X2072 VSSD D5 level_tx_8bit_0/level_tx_1bit_0[5]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2073 8_bit_dac_0/D5 level_tx_8bit_0/level_tx_1bit_0[5]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2074 level_tx_8bit_0/level_tx_1bit_0[5]/a_n1353_675# D5 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X2075 8_bit_dac_0/D5 level_tx_8bit_0/level_tx_1bit_0[5]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2076 level_tx_8bit_0/level_tx_1bit_0[6]/a_n1423_1248# 8_bit_dac_0/D6 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2077 VSSD D6 level_tx_8bit_0/level_tx_1bit_0[6]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X2078 VSSD D6 level_tx_8bit_0/level_tx_1bit_0[6]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2079 8_bit_dac_0/D6 level_tx_8bit_0/level_tx_1bit_0[6]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2080 level_tx_8bit_0/level_tx_1bit_0[6]/a_n1353_675# D6 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X2081 8_bit_dac_0/D6 level_tx_8bit_0/level_tx_1bit_0[6]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2082 level_tx_8bit_0/level_tx_1bit_0[7]/a_n1423_1248# 8_bit_dac_0/D7 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2083 VSSD D7 level_tx_8bit_0/level_tx_1bit_0[7]/a_n1353_675# VSSD sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.122 ps=1.42 w=0.42 l=0.2
X2084 VSSD D7 level_tx_8bit_0/level_tx_1bit_0[7]/a_n1423_1248# VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X2085 8_bit_dac_0/D7 level_tx_8bit_0/level_tx_1bit_0[7]/a_n1423_1248# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X2086 level_tx_8bit_0/level_tx_1bit_0[7]/a_n1353_675# D7 VCCD VCCD sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.2
X2087 8_bit_dac_0/D7 level_tx_8bit_0/level_tx_1bit_0[7]/a_n1353_675# VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X2088 VSSA opamp_0/a_3246_n774# VOUT_BUF VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=1
X2089 VOUT_BUF opamp_0/a_3246_n774# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X2090 VDDA opamp_0/a_1618_n334# VOUT_BUF VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X2091 VDDA opamp_0/a_394_n920# opamp_0/a_1704_376# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=1
X2092 opamp_0/a_1704_376# VOUT_BUF opamp_0/a_1446_376# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=1
X2093 VDDA opamp_0/a_1618_n334# VOUT_BUF VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.6 as=1.16 ps=8.29 w=8 l=1
X2094 opamp_0/a_408_552# VSSA VSSA sky130_fd_pr__res_generic_nd__hv w=0.48 l=4.46
X2095 VSSA opamp_0/a_1022_n914# opamp_0/a_2158_n774# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
X2096 opamp_0/a_2158_n774# VOUT_BUF opamp_0/a_1900_n774# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=1
X2097 VSSA opamp_0/a_2894_292# opamp_0/a_2894_292# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X2098 opamp_0/a_1022_n914# opamp_0/a_394_n920# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.6 as=1.16 ps=8.29 w=8 l=1
X2099 opamp_0/a_1776_n834# opamp_0/a_408_552# opamp_0/a_1618_n334# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X2100 VSSA opamp_0/a_1022_n914# opamp_0/a_1446_376# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X2101 opamp_0/a_2894_292# opamp_0/a_408_552# opamp_0/a_1900_n774# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X2102 VDDA opamp_0/a_408_552# VSSA sky130_fd_pr__res_generic_nd__hv w=0.42 l=8.32
X2103 opamp_0/a_2416_n774# opamp_0/a_394_n920# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=1
X2104 VDDA opamp_0/a_394_n920# opamp_0/a_394_n920# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.29 as=2.32 ps=16.6 w=8 l=1
X2105 opamp_0/a_1446_376# opamp_0/a_408_552# opamp_0/a_1300_n354# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X2106 VOUT_BUF opamp_0/a_3246_n774# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=1
X2107 opamp_0/a_2416_n774# VOUT opamp_0/a_2158_n774# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=1
X2108 VOUT_BUF opamp_0/a_1618_n334# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.29 as=2.32 ps=16.6 w=8 l=1
X2109 VOUT_BUF opamp_0/a_1618_n334# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.29 as=1.16 ps=8.29 w=8 l=1
X2110 opamp_0/a_1776_n834# VOUT opamp_0/a_1704_376# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=1
X2111 opamp_0/a_1618_n334# opamp_0/a_1300_n354# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.6 as=1.16 ps=8.29 w=8 l=1
X2112 VSSA opamp_0/a_3246_n774# VOUT_BUF VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=0.58 ps=4.29 w=4 l=1
X2113 VSSA opamp_0/a_1022_n914# opamp_0/a_1022_n914# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
X2114 opamp_0/a_1776_n834# opamp_0/a_1022_n914# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X2115 opamp_0/a_3246_n774# opamp_0/a_2894_292# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X2116 VSSA opamp_0/a_394_n920# VSSA sky130_fd_pr__res_generic_nd__hv w=0.41 l=15.7
X2117 VDDA opamp_0/a_394_n920# opamp_0/a_1900_n774# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=1
X2118 opamp_0/a_3246_n774# opamp_0/a_408_552# opamp_0/a_2416_n774# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X2119 VDDA opamp_0/a_1300_n354# opamp_0/a_1300_n354# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.29 as=2.32 ps=16.6 w=8 l=1
.ends

X1 VDDA VSSD VCCD VSSA D0 D1 D2 D3 D4 D5 D6 D7 VOUT VREFH VOUT_BUF x8_bit_dac_tx_buffer
   
.param mc_mm_switch=0
.param mc_pr_switch=0
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

V1 VSSA 0 dc 0
V2 VDDA 0 dc 3.3

V3 VSSD 0 dc 0
V4 VCCD 0 dc 1.8

V5 VREFH 0 dc 3.3

V6  D0 0 PULSE(0 1.8 0 1n 1n 1u 2u)
V7  D1 0 PULSE(0 1.8 0 1n 1n 2u 4u)
V8  D2 0 PULSE(0 1.8 0 1n 1n 4u 8u)
V9  D3 0 PULSE(0 1.8 0 1n 1n 8u 16u)
V10 D4 0 PULSE(0 1.8 0 1n 1n 16u 32u)
V11 D5 0 PULSE(0 1.8 0 1n 1n 32u 64u)
V12 D6 0 PULSE(0 1.8 0 1n 1n 64u 128u)
V13 D7 0 PULSE(0 1.8 0 1n 1n 128u 256u)

.tran 5u 60u
.control
run
plot VOUT VOUT_BUF
.endc
.end
