** sch_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/2_bit_dac/2_bit_dac.sch
.subckt 2_bit_dac D1 D0 D0_BUF D1_BUF VOUT VREFL VREFH VCC VSS
*.PININFO D1:I D0:I D0_BUF:O D1_BUF:O VOUT:O VREFL:I VREFH:I VCC:B VSS:B
R2 VREFH net1 sky130_fd_pr__res_generic_po W=1 L=1 m=1
x1 VCC D0_BUF D0 net1 VSS VINL VINH VREFL switch_2n
x2 VCC D1 D1_BUF VSS VINH VOUT VINL switch_n
.ends

* expanding   symbol:  /foss/designs/8_bit_dac/Switch_2n/switch_2n.sym # of pins=8
** sym_path: /foss/designs/8_bit_dac/Switch_2n/switch_2n.sym
** sch_path: /foss/designs/8_bit_dac/Switch_2n/switch_2n.sch
.subckt switch_2n VCC DX_BUF DX VREFH VSS VOUTL VOUTH VREFL
*.PININFO VCC:B VSS:B VOUTL:O DX:I VOUTH:O DX_BUF:O VREFH:I VREFL:I
XM1 net1 DX VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM2 net1 DX VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM3 DX_BUF net1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM4 DX_BUF net1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM5 VOUTL net1 VREFL VREFL sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM6 VOUTL net1 net2 net2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM7 VREFL DX_BUF VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM8 net2 DX_BUF VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM9 VOUTH net1 net3 net3 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM10 VOUTH net1 VREFH VREFH sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM11 net3 DX_BUF VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM12 VREFH DX_BUF VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
R1 net3 VREFH sky130_fd_pr__res_generic_po W=1 L=1 m=1
R2 net2 net3 sky130_fd_pr__res_generic_po W=1 L=1 m=1
R3 VREFL net2 sky130_fd_pr__res_generic_po W=1 L=1 m=1
.ends


* expanding   symbol:  /foss/designs/8_bit_dac/Switch_n/switch_n.sym # of pins=7
** sym_path: /foss/designs/8_bit_dac/Switch_n/switch_n.sym
** sch_path: /foss/designs/8_bit_dac/Switch_n/switch_n.sch
.subckt switch_n VCC DX DX_BUF VSS VREFH VOUT VREFL
*.PININFO VCC:B VSS:B DX_BUF:O VOUT:O DX:I VREFH:I VREFL:I
XM1 net1 DX VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM2 net1 DX VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM3 DX_BUF net1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM4 DX_BUF net1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM5 VOUT net1 VREFL VREFL sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM6 VOUT net1 VREFH VREFH sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM7 VREFL DX_BUF VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM8 VREFH DX_BUF VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
.ends

.end
