magic
tech sky130A
magscale 1 2
timestamp 1690460648
<< nwell >>
rect 7755 5346 8777 5703
rect 7755 5340 8243 5346
rect 7755 5300 8224 5340
rect 7755 5296 8243 5300
rect 8311 5296 8777 5346
rect 7755 5165 8777 5296
<< psubdiff >>
rect 7859 4910 8294 4943
rect 7859 4828 7892 4910
rect 8264 4828 8294 4910
rect 7859 4803 8294 4828
<< mvnsubdiff >>
rect 7824 5602 8710 5633
rect 7824 5516 7850 5602
rect 8686 5516 8710 5602
rect 7824 5493 8710 5516
<< psubdiffcont >>
rect 7892 4828 8264 4910
<< mvnsubdiffcont >>
rect 7850 5516 8686 5602
<< poly >>
rect 7933 5190 8033 5229
rect 7933 5156 7968 5190
rect 8002 5156 8033 5190
rect 7933 5082 8033 5156
rect 8221 5195 8321 5229
rect 8221 5161 8250 5195
rect 8284 5161 8321 5195
rect 8221 5082 8321 5161
rect 8509 5193 8609 5229
rect 8509 5159 8547 5193
rect 8581 5159 8609 5193
rect 8509 5092 8609 5159
<< polycont >>
rect 7968 5156 8002 5190
rect 8250 5161 8284 5195
rect 8547 5159 8581 5193
<< locali >>
rect 7824 5602 8710 5633
rect 7824 5516 7850 5602
rect 8686 5516 8710 5602
rect 7824 5493 8710 5516
rect 7968 5190 8002 5206
rect 8234 5161 8250 5195
rect 8284 5161 8300 5195
rect 8531 5159 8547 5193
rect 8581 5159 8597 5193
rect 7968 5140 8002 5156
rect 7859 4910 8294 4943
rect 7859 4828 7892 4910
rect 8264 4828 8294 4910
rect 7859 4803 8294 4828
<< viali >>
rect 7850 5516 8686 5602
rect 7968 5156 8002 5190
rect 8250 5161 8284 5195
rect 8547 5159 8581 5193
rect 7892 4828 8264 4910
<< metal1 >>
rect 7824 5602 8710 5633
rect 7824 5516 7850 5602
rect 8686 5516 8710 5602
rect 7824 5493 8710 5516
rect 7881 5409 7927 5493
rect 8463 5351 8497 5364
rect 8166 5345 8218 5351
rect 8166 5287 8218 5293
rect 8454 5345 8506 5351
rect 8454 5287 8506 5293
rect 7962 5199 8008 5202
rect 7953 5147 7959 5199
rect 8011 5147 8017 5199
rect 8045 5195 8079 5284
rect 8175 5274 8209 5287
rect 8606 5284 8612 5336
rect 8664 5284 8670 5336
rect 8234 5195 8298 5204
rect 8045 5161 8250 5195
rect 8284 5161 8298 5195
rect 7962 5144 8008 5147
rect 8045 5049 8079 5161
rect 8234 5152 8298 5161
rect 8166 5070 8218 5076
rect 7881 4943 7927 5029
rect 8166 5012 8218 5018
rect 8175 5011 8209 5012
rect 8333 4968 8367 5284
rect 8401 5150 8407 5202
rect 8459 5193 8465 5202
rect 8531 5193 8595 5202
rect 8459 5159 8547 5193
rect 8581 5159 8599 5193
rect 8459 5150 8465 5159
rect 8531 5150 8595 5159
rect 8463 5086 8497 5094
rect 8621 5086 8655 5115
rect 8454 5080 8506 5086
rect 8621 5084 8656 5086
rect 8454 5022 8506 5028
rect 8612 5078 8664 5084
rect 8612 5020 8664 5026
rect 8621 4968 8655 5020
rect 7859 4910 8294 4943
rect 8333 4934 8655 4968
rect 7859 4828 7892 4910
rect 8264 4828 8294 4910
rect 7859 4803 8294 4828
<< via1 >>
rect 7850 5516 8686 5602
rect 8166 5293 8218 5345
rect 8454 5293 8506 5345
rect 7959 5190 8011 5199
rect 7959 5156 7968 5190
rect 7968 5156 8002 5190
rect 8002 5156 8011 5190
rect 7959 5147 8011 5156
rect 8612 5284 8664 5336
rect 8166 5018 8218 5070
rect 8407 5150 8459 5202
rect 8454 5028 8506 5080
rect 8612 5026 8664 5078
rect 7892 4828 8264 4910
<< metal2 >>
rect 7824 5602 8710 5633
rect 7824 5516 7850 5602
rect 8686 5516 8710 5602
rect 7824 5493 8710 5516
rect 8176 5420 8576 5454
rect 8176 5345 8210 5420
rect 8160 5336 8166 5345
rect 7764 5302 8166 5336
rect 8160 5293 8166 5302
rect 8218 5293 8224 5345
rect 8448 5336 8454 5345
rect 8253 5302 8454 5336
rect 7959 5203 8011 5205
rect 7946 5190 7955 5203
rect 7870 5156 7955 5190
rect 7946 5143 7955 5156
rect 8015 5143 8024 5203
rect 7959 5141 8011 5143
rect 8253 5134 8287 5302
rect 8448 5293 8454 5302
rect 8506 5293 8512 5345
rect 8407 5206 8459 5208
rect 8394 5146 8403 5206
rect 8463 5146 8472 5206
rect 8407 5144 8459 5146
rect 8175 5100 8287 5134
rect 8175 5070 8209 5100
rect 8160 5061 8166 5070
rect 7753 5027 8166 5061
rect 8160 5018 8166 5027
rect 8218 5018 8224 5070
rect 8448 5028 8454 5080
rect 8506 5071 8512 5080
rect 8542 5071 8576 5420
rect 8612 5336 8664 5342
rect 8664 5294 8777 5328
rect 8612 5278 8664 5284
rect 8621 5078 8655 5278
rect 8506 5037 8576 5071
rect 8506 5028 8512 5037
rect 8606 5026 8612 5078
rect 8664 5026 8670 5078
rect 7859 4910 8294 4943
rect 7859 4828 7892 4910
rect 8264 4828 8294 4910
rect 7859 4803 8294 4828
<< via2 >>
rect 7850 5516 8686 5602
rect 7955 5199 8015 5203
rect 7955 5147 7959 5199
rect 7959 5147 8011 5199
rect 8011 5147 8015 5199
rect 7955 5143 8015 5147
rect 8403 5202 8463 5206
rect 8403 5150 8407 5202
rect 8407 5150 8459 5202
rect 8459 5150 8463 5202
rect 8403 5146 8463 5150
rect 7892 4828 8264 4910
<< metal3 >>
rect 7750 5602 8782 5633
rect 7750 5516 7850 5602
rect 8686 5516 8782 5602
rect 7750 5493 8782 5516
rect 7950 5206 8020 5208
rect 8398 5206 8468 5211
rect 7950 5203 8403 5206
rect 7950 5143 7955 5203
rect 8015 5146 8403 5203
rect 8463 5203 8468 5206
rect 8463 5146 8474 5203
rect 8015 5143 8474 5146
rect 7950 5138 8020 5143
rect 8398 5141 8468 5143
rect 7750 4910 8782 4943
rect 7750 4828 7892 4910
rect 8264 4828 8782 4910
rect 7750 4803 8782 4828
use sky130_fd_pr__nfet_g5v0d10v5_NQZZCX  sky130_fd_pr__nfet_g5v0d10v5_NQZZCX_0
timestamp 1690460607
transform 1 0 8271 0 1 5044
box -108 -68 108 68
use sky130_fd_pr__nfet_g5v0d10v5_NQZZCX  sky130_fd_pr__nfet_g5v0d10v5_NQZZCX_1
timestamp 1690460607
transform 1 0 7983 0 1 5044
box -108 -68 108 68
use sky130_fd_pr__nfet_g5v0d10v5_NQZZCX  sky130_fd_pr__nfet_g5v0d10v5_NQZZCX_2
timestamp 1690460607
transform 1 0 8559 0 1 5054
box -108 -68 108 68
use sky130_fd_pr__pfet_g5v0d10v5_AWMFT3  sky130_fd_pr__pfet_g5v0d10v5_AWMFT3_0
timestamp 1690460607
transform 1 0 7983 0 1 5327
box -174 -150 174 150
use sky130_fd_pr__pfet_g5v0d10v5_AWMFT3  sky130_fd_pr__pfet_g5v0d10v5_AWMFT3_2
timestamp 1690460607
transform 1 0 8559 0 1 5327
box -174 -150 174 150
use sky130_fd_pr__pfet_g5v0d10v5_AWMFT3  sky130_fd_pr__pfet_g5v0d10v5_AWMFT3_3
timestamp 1690460607
transform 1 0 8271 0 1 5327
box -174 -150 174 150
<< labels >>
flabel metal3 s 7769 5567 7769 5567 0 FreeSans 320 0 0 0 VCC
flabel metal3 s 7791 4855 7791 4855 0 FreeSans 320 0 0 0 VSS
flabel metal2 s 8756 5314 8756 5314 0 FreeSans 320 0 0 0 OUT
flabel metal2 s 7888 5170 7888 5170 0 FreeSans 320 0 0 0 SEL
flabel metal2 s 7786 5316 7786 5316 0 FreeSans 320 0 0 0 A
flabel metal2 s 7775 5044 7775 5044 0 FreeSans 320 0 0 0 B
<< end >>
