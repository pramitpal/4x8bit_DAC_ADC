magic
tech sky130A
magscale 1 2
timestamp 1685680497
<< nwell >>
rect -6382 196 -5754 204
rect -6382 -316 -5062 196
<< pwell >>
rect -5682 -362 -5106 -360
rect -6342 -512 -5106 -362
rect -6342 -514 -5766 -512
rect -6342 -518 -5776 -514
rect -6368 -710 -5776 -518
<< mvnmos >>
rect -6258 -488 -6158 -388
rect -5950 -488 -5850 -388
rect -5598 -486 -5498 -386
rect -5290 -486 -5190 -386
<< mvpmos >>
rect -6258 -250 -6158 -50
rect -5950 -250 -5850 -50
rect -5598 -250 -5498 -50
rect -5290 -250 -5190 -50
<< mvndiff >>
rect -6316 -421 -6258 -388
rect -6316 -455 -6304 -421
rect -6270 -455 -6258 -421
rect -6316 -488 -6258 -455
rect -6158 -421 -6100 -388
rect -6158 -455 -6146 -421
rect -6112 -455 -6100 -421
rect -6158 -488 -6100 -455
rect -6008 -421 -5950 -388
rect -6008 -455 -5996 -421
rect -5962 -455 -5950 -421
rect -6008 -488 -5950 -455
rect -5850 -421 -5792 -388
rect -5850 -455 -5838 -421
rect -5804 -455 -5792 -421
rect -5850 -488 -5792 -455
rect -5656 -419 -5598 -386
rect -5656 -453 -5644 -419
rect -5610 -453 -5598 -419
rect -5656 -486 -5598 -453
rect -5498 -419 -5440 -386
rect -5498 -453 -5486 -419
rect -5452 -453 -5440 -419
rect -5498 -486 -5440 -453
rect -5348 -419 -5290 -386
rect -5348 -453 -5336 -419
rect -5302 -453 -5290 -419
rect -5348 -486 -5290 -453
rect -5190 -419 -5132 -386
rect -5190 -453 -5178 -419
rect -5144 -453 -5132 -419
rect -5190 -486 -5132 -453
<< mvpdiff >>
rect -6316 -65 -6258 -50
rect -6316 -99 -6304 -65
rect -6270 -99 -6258 -65
rect -6316 -133 -6258 -99
rect -6316 -167 -6304 -133
rect -6270 -167 -6258 -133
rect -6316 -201 -6258 -167
rect -6316 -235 -6304 -201
rect -6270 -235 -6258 -201
rect -6316 -250 -6258 -235
rect -6158 -65 -6100 -50
rect -6158 -99 -6146 -65
rect -6112 -99 -6100 -65
rect -6158 -133 -6100 -99
rect -6158 -167 -6146 -133
rect -6112 -167 -6100 -133
rect -6158 -201 -6100 -167
rect -6158 -235 -6146 -201
rect -6112 -235 -6100 -201
rect -6158 -250 -6100 -235
rect -6008 -65 -5950 -50
rect -6008 -99 -5996 -65
rect -5962 -99 -5950 -65
rect -6008 -133 -5950 -99
rect -6008 -167 -5996 -133
rect -5962 -167 -5950 -133
rect -6008 -201 -5950 -167
rect -6008 -235 -5996 -201
rect -5962 -235 -5950 -201
rect -6008 -250 -5950 -235
rect -5850 -65 -5792 -50
rect -5850 -99 -5838 -65
rect -5804 -99 -5792 -65
rect -5850 -133 -5792 -99
rect -5850 -167 -5838 -133
rect -5804 -167 -5792 -133
rect -5850 -201 -5792 -167
rect -5850 -235 -5838 -201
rect -5804 -235 -5792 -201
rect -5850 -250 -5792 -235
rect -5656 -65 -5598 -50
rect -5656 -99 -5644 -65
rect -5610 -99 -5598 -65
rect -5656 -133 -5598 -99
rect -5656 -167 -5644 -133
rect -5610 -167 -5598 -133
rect -5656 -201 -5598 -167
rect -5656 -235 -5644 -201
rect -5610 -235 -5598 -201
rect -5656 -250 -5598 -235
rect -5498 -65 -5440 -50
rect -5498 -99 -5486 -65
rect -5452 -99 -5440 -65
rect -5498 -133 -5440 -99
rect -5498 -167 -5486 -133
rect -5452 -167 -5440 -133
rect -5498 -201 -5440 -167
rect -5498 -235 -5486 -201
rect -5452 -235 -5440 -201
rect -5498 -250 -5440 -235
rect -5348 -65 -5290 -50
rect -5348 -99 -5336 -65
rect -5302 -99 -5290 -65
rect -5348 -133 -5290 -99
rect -5348 -167 -5336 -133
rect -5302 -167 -5290 -133
rect -5348 -201 -5290 -167
rect -5348 -235 -5336 -201
rect -5302 -235 -5290 -201
rect -5348 -250 -5290 -235
rect -5190 -65 -5132 -50
rect -5190 -99 -5178 -65
rect -5144 -99 -5132 -65
rect -5190 -133 -5132 -99
rect -5190 -167 -5178 -133
rect -5144 -167 -5132 -133
rect -5190 -201 -5132 -167
rect -5190 -235 -5178 -201
rect -5144 -235 -5132 -201
rect -5190 -250 -5132 -235
<< mvndiffc >>
rect -6304 -455 -6270 -421
rect -6146 -455 -6112 -421
rect -5996 -455 -5962 -421
rect -5838 -455 -5804 -421
rect -5644 -453 -5610 -419
rect -5486 -453 -5452 -419
rect -5336 -453 -5302 -419
rect -5178 -453 -5144 -419
<< mvpdiffc >>
rect -6304 -99 -6270 -65
rect -6304 -167 -6270 -133
rect -6304 -235 -6270 -201
rect -6146 -99 -6112 -65
rect -6146 -167 -6112 -133
rect -6146 -235 -6112 -201
rect -5996 -99 -5962 -65
rect -5996 -167 -5962 -133
rect -5996 -235 -5962 -201
rect -5838 -99 -5804 -65
rect -5838 -167 -5804 -133
rect -5838 -235 -5804 -201
rect -5644 -99 -5610 -65
rect -5644 -167 -5610 -133
rect -5644 -235 -5610 -201
rect -5486 -99 -5452 -65
rect -5486 -167 -5452 -133
rect -5486 -235 -5452 -201
rect -5336 -99 -5302 -65
rect -5336 -167 -5302 -133
rect -5336 -235 -5302 -201
rect -5178 -99 -5144 -65
rect -5178 -167 -5144 -133
rect -5178 -235 -5144 -201
<< psubdiff >>
rect -6342 -597 -5802 -544
rect -6342 -631 -6293 -597
rect -6259 -631 -6225 -597
rect -6191 -631 -6157 -597
rect -6123 -631 -6089 -597
rect -6055 -631 -6021 -597
rect -5987 -631 -5953 -597
rect -5919 -631 -5885 -597
rect -5851 -631 -5802 -597
rect -6342 -684 -5802 -631
<< mvnsubdiff >>
rect -6312 93 -5792 136
rect -6312 59 -6273 93
rect -6239 59 -6205 93
rect -6171 59 -6137 93
rect -6103 59 -6069 93
rect -6035 59 -6001 93
rect -5967 59 -5933 93
rect -5899 59 -5865 93
rect -5831 59 -5792 93
rect -6312 16 -5792 59
<< psubdiffcont >>
rect -6293 -631 -6259 -597
rect -6225 -631 -6191 -597
rect -6157 -631 -6123 -597
rect -6089 -631 -6055 -597
rect -6021 -631 -5987 -597
rect -5953 -631 -5919 -597
rect -5885 -631 -5851 -597
<< mvnsubdiffcont >>
rect -6273 59 -6239 93
rect -6205 59 -6171 93
rect -6137 59 -6103 93
rect -6069 59 -6035 93
rect -6001 59 -5967 93
rect -5933 59 -5899 93
rect -5865 59 -5831 93
<< poly >>
rect -6258 -50 -6158 -24
rect -5950 -50 -5850 -24
rect -5598 -50 -5498 -24
rect -5290 -50 -5190 -24
rect -6392 -291 -6326 -283
rect -6258 -291 -6158 -250
rect -6392 -293 -6158 -291
rect -6392 -327 -6376 -293
rect -6342 -327 -6158 -293
rect -6392 -330 -6158 -327
rect -6392 -337 -6326 -330
rect -6258 -388 -6158 -330
rect -6078 -300 -6012 -292
rect -5950 -300 -5850 -250
rect -6078 -302 -5850 -300
rect -6078 -336 -6062 -302
rect -6028 -336 -5850 -302
rect -6078 -339 -5850 -336
rect -6078 -346 -6012 -339
rect -5950 -388 -5850 -339
rect -5756 -308 -5690 -298
rect -5598 -308 -5498 -250
rect -5756 -342 -5740 -308
rect -5706 -342 -5498 -308
rect -5419 -290 -5365 -274
rect -5419 -324 -5409 -290
rect -5375 -292 -5365 -290
rect -5290 -292 -5190 -250
rect -5375 -323 -5190 -292
rect -5375 -324 -5365 -323
rect -5419 -340 -5365 -324
rect -5756 -343 -5498 -342
rect -5756 -352 -5690 -343
rect -5598 -386 -5498 -343
rect -5290 -386 -5190 -323
rect -6258 -514 -6158 -488
rect -5950 -514 -5850 -488
rect -5598 -512 -5498 -486
rect -5290 -512 -5190 -486
<< polycont >>
rect -6376 -327 -6342 -293
rect -6062 -336 -6028 -302
rect -5740 -342 -5706 -308
rect -5409 -324 -5375 -290
<< locali >>
rect -6322 93 -5782 146
rect -6322 59 -6273 93
rect -6215 59 -6205 93
rect -6143 59 -6137 93
rect -6071 59 -6069 93
rect -6035 59 -6033 93
rect -5967 59 -5961 93
rect -5899 59 -5889 93
rect -5831 59 -5782 93
rect -6322 6 -5782 59
rect -6304 -65 -6270 -46
rect -6304 -133 -6270 -131
rect -6304 -169 -6270 -167
rect -6304 -254 -6270 -235
rect -6146 -65 -6112 -46
rect -6146 -133 -6112 -131
rect -6146 -169 -6112 -167
rect -6146 -254 -6112 -235
rect -5996 -65 -5962 -46
rect -5996 -133 -5962 -131
rect -5996 -169 -5962 -167
rect -5996 -254 -5962 -235
rect -5838 -65 -5804 -46
rect -5838 -133 -5804 -131
rect -5838 -169 -5804 -167
rect -5838 -254 -5804 -235
rect -5644 -65 -5610 -46
rect -5644 -133 -5610 -131
rect -5644 -169 -5610 -167
rect -5644 -254 -5610 -235
rect -5486 -65 -5452 -46
rect -5486 -133 -5452 -131
rect -5486 -169 -5452 -167
rect -5486 -254 -5452 -235
rect -5336 -65 -5302 -46
rect -5336 -133 -5302 -131
rect -5336 -169 -5302 -167
rect -5336 -254 -5302 -235
rect -5178 -65 -5144 -46
rect -5178 -133 -5144 -131
rect -5178 -169 -5144 -167
rect -5178 -254 -5144 -235
rect -6376 -290 -6342 -277
rect -6378 -293 -6339 -290
rect -6378 -327 -6376 -293
rect -6342 -327 -6339 -293
rect -6062 -299 -6028 -286
rect -6378 -329 -6339 -327
rect -6064 -302 -6025 -299
rect -6376 -343 -6342 -329
rect -6064 -336 -6062 -302
rect -6028 -336 -6025 -302
rect -6064 -338 -6025 -336
rect -5740 -307 -5706 -292
rect -5740 -308 -5705 -307
rect -6062 -352 -6028 -338
rect -5706 -342 -5705 -308
rect -5425 -324 -5409 -290
rect -5375 -324 -5359 -290
rect -5740 -358 -5706 -342
rect -6304 -421 -6270 -384
rect -6304 -492 -6270 -455
rect -6146 -421 -6112 -384
rect -6146 -492 -6112 -455
rect -5996 -421 -5962 -384
rect -5996 -492 -5962 -455
rect -5838 -421 -5804 -384
rect -5838 -492 -5804 -455
rect -5644 -419 -5610 -382
rect -5644 -490 -5610 -453
rect -5486 -419 -5452 -382
rect -5486 -490 -5452 -453
rect -5336 -419 -5302 -382
rect -5336 -490 -5302 -453
rect -5178 -419 -5144 -382
rect -5178 -490 -5144 -453
rect -6342 -597 -5802 -544
rect -6342 -631 -6305 -597
rect -6259 -631 -6233 -597
rect -6191 -631 -6161 -597
rect -6123 -631 -6089 -597
rect -6055 -631 -6021 -597
rect -5983 -631 -5953 -597
rect -5911 -631 -5885 -597
rect -5839 -631 -5802 -597
rect -6342 -684 -5802 -631
<< viali >>
rect -6249 59 -6239 93
rect -6239 59 -6215 93
rect -6177 59 -6171 93
rect -6171 59 -6143 93
rect -6105 59 -6103 93
rect -6103 59 -6071 93
rect -6033 59 -6001 93
rect -6001 59 -5999 93
rect -5961 59 -5933 93
rect -5933 59 -5927 93
rect -5889 59 -5865 93
rect -5865 59 -5855 93
rect -6304 -99 -6270 -97
rect -6304 -131 -6270 -99
rect -6304 -201 -6270 -169
rect -6304 -203 -6270 -201
rect -6146 -99 -6112 -97
rect -6146 -131 -6112 -99
rect -6146 -201 -6112 -169
rect -6146 -203 -6112 -201
rect -5996 -99 -5962 -97
rect -5996 -131 -5962 -99
rect -5996 -201 -5962 -169
rect -5996 -203 -5962 -201
rect -5838 -99 -5804 -97
rect -5838 -131 -5804 -99
rect -5838 -201 -5804 -169
rect -5838 -203 -5804 -201
rect -5644 -99 -5610 -97
rect -5644 -131 -5610 -99
rect -5644 -201 -5610 -169
rect -5644 -203 -5610 -201
rect -5486 -99 -5452 -97
rect -5486 -131 -5452 -99
rect -5486 -201 -5452 -169
rect -5486 -203 -5452 -201
rect -5336 -99 -5302 -97
rect -5336 -131 -5302 -99
rect -5336 -201 -5302 -169
rect -5336 -203 -5302 -201
rect -5178 -99 -5144 -97
rect -5178 -131 -5144 -99
rect -5178 -201 -5144 -169
rect -5178 -203 -5144 -201
rect -6376 -327 -6342 -293
rect -6062 -336 -6028 -302
rect -5740 -342 -5706 -308
rect -5409 -324 -5375 -290
rect -6304 -455 -6270 -421
rect -6146 -455 -6112 -421
rect -5996 -455 -5962 -421
rect -5838 -455 -5804 -421
rect -5644 -453 -5610 -419
rect -5486 -453 -5452 -419
rect -5336 -453 -5302 -419
rect -5178 -453 -5144 -419
rect -6305 -631 -6293 -597
rect -6293 -631 -6271 -597
rect -6233 -631 -6225 -597
rect -6225 -631 -6199 -597
rect -6161 -631 -6157 -597
rect -6157 -631 -6127 -597
rect -6089 -631 -6055 -597
rect -6017 -631 -5987 -597
rect -5987 -631 -5983 -597
rect -5945 -631 -5919 -597
rect -5919 -631 -5911 -597
rect -5873 -631 -5851 -597
rect -5851 -631 -5839 -597
<< metal1 >>
rect -6322 102 -5782 146
rect -6322 50 -6270 102
rect -6218 93 -6206 102
rect -6154 93 -6142 102
rect -6090 93 -6078 102
rect -6026 93 -6014 102
rect -5962 93 -5950 102
rect -5898 93 -5886 102
rect -6215 59 -6206 93
rect -6143 59 -6142 93
rect -5962 59 -5961 93
rect -5898 59 -5889 93
rect -6218 50 -6206 59
rect -6154 50 -6142 59
rect -6090 50 -6078 59
rect -6026 50 -6014 59
rect -5962 50 -5950 59
rect -5898 50 -5886 59
rect -5834 50 -5782 102
rect -6322 6 -5782 50
rect -6305 -50 -6259 6
rect -6310 -51 -6259 -50
rect -6310 -97 -6264 -51
rect -6310 -131 -6304 -97
rect -6270 -131 -6264 -97
rect -6310 -169 -6264 -131
rect -6310 -203 -6304 -169
rect -6270 -203 -6264 -169
rect -6310 -250 -6264 -203
rect -6152 -97 -6106 -50
rect -6152 -131 -6146 -97
rect -6112 -131 -6106 -97
rect -6152 -169 -6106 -131
rect -6152 -203 -6146 -169
rect -6112 -203 -6106 -169
rect -6152 -250 -6106 -203
rect -6002 -97 -5956 6
rect -5488 -50 -5449 195
rect -5171 -50 -5142 207
rect -6002 -131 -5996 -97
rect -5962 -131 -5956 -97
rect -6002 -169 -5956 -131
rect -6002 -203 -5996 -169
rect -5962 -203 -5956 -169
rect -6002 -250 -5956 -203
rect -5844 -97 -5798 -50
rect -5844 -131 -5838 -97
rect -5804 -131 -5798 -97
rect -5650 -97 -5604 -50
rect -5650 -123 -5644 -97
rect -5844 -169 -5798 -131
rect -5844 -203 -5838 -169
rect -5804 -203 -5798 -169
rect -5761 -125 -5644 -123
rect -5761 -177 -5754 -125
rect -5702 -131 -5644 -125
rect -5610 -131 -5604 -97
rect -5702 -169 -5604 -131
rect -5702 -177 -5644 -169
rect -5761 -178 -5644 -177
rect -5844 -250 -5798 -203
rect -5650 -203 -5644 -178
rect -5610 -203 -5604 -169
rect -5650 -250 -5604 -203
rect -5492 -97 -5446 -50
rect -5492 -131 -5486 -97
rect -5452 -130 -5446 -97
rect -5342 -97 -5296 -50
rect -5342 -130 -5336 -97
rect -5452 -131 -5336 -130
rect -5302 -131 -5296 -97
rect -5492 -169 -5296 -131
rect -5492 -203 -5486 -169
rect -5452 -196 -5336 -169
rect -5452 -203 -5446 -196
rect -5492 -250 -5446 -203
rect -5342 -203 -5336 -196
rect -5302 -203 -5296 -169
rect -5342 -250 -5296 -203
rect -5184 -97 -5138 -50
rect -5184 -131 -5178 -97
rect -5144 -131 -5138 -97
rect -5019 -126 -4989 -117
rect -5184 -169 -5138 -131
rect -5184 -203 -5178 -169
rect -5144 -203 -5138 -169
rect -5036 -178 -5030 -126
rect -4978 -178 -4972 -126
rect -5184 -250 -5138 -203
rect -5020 -219 -4989 -178
rect -6491 -335 -6485 -283
rect -6433 -290 -6427 -283
rect -6384 -290 -6333 -278
rect -6433 -293 -6333 -290
rect -6433 -327 -6376 -293
rect -6342 -327 -6333 -293
rect -6433 -329 -6333 -327
rect -6433 -335 -6427 -329
rect -6384 -341 -6333 -329
rect -6149 -299 -6110 -250
rect -6070 -292 -6019 -287
rect -6076 -299 -6070 -292
rect -6149 -338 -6070 -299
rect -6149 -388 -6110 -338
rect -6076 -344 -6070 -338
rect -6018 -344 -6012 -292
rect -5840 -306 -5801 -250
rect -5746 -306 -5699 -295
rect -5840 -308 -5699 -306
rect -5840 -341 -5740 -308
rect -6070 -350 -6019 -344
rect -5840 -388 -5801 -341
rect -5746 -342 -5740 -341
rect -5706 -342 -5699 -308
rect -5746 -354 -5699 -342
rect -6310 -421 -6264 -388
rect -6310 -455 -6304 -421
rect -6270 -455 -6264 -421
rect -6310 -488 -6264 -455
rect -6152 -421 -6106 -388
rect -6152 -455 -6146 -421
rect -6112 -455 -6106 -421
rect -6002 -421 -5956 -388
rect -6002 -450 -5996 -421
rect -6152 -488 -6106 -455
rect -6004 -455 -5996 -450
rect -5962 -455 -5956 -421
rect -6004 -488 -5956 -455
rect -5844 -421 -5798 -388
rect -5844 -455 -5838 -421
rect -5804 -455 -5798 -421
rect -5844 -488 -5798 -455
rect -6310 -544 -6266 -488
rect -6004 -544 -5957 -488
rect -6342 -588 -5802 -544
rect -6342 -597 -6290 -588
rect -6238 -597 -6226 -588
rect -6342 -631 -6305 -597
rect -6238 -631 -6233 -597
rect -6342 -640 -6290 -631
rect -6238 -640 -6226 -631
rect -6174 -640 -6162 -588
rect -6110 -640 -6098 -588
rect -6046 -640 -6034 -588
rect -5982 -640 -5970 -588
rect -5918 -597 -5906 -588
rect -5854 -597 -5802 -588
rect -5911 -631 -5906 -597
rect -5839 -631 -5802 -597
rect -5918 -640 -5906 -631
rect -5854 -640 -5802 -631
rect -6342 -684 -5802 -640
rect -6487 -789 -6481 -737
rect -6429 -744 -6423 -737
rect -5740 -744 -5701 -354
rect -5488 -386 -5449 -250
rect -5418 -281 -5366 -275
rect -5421 -330 -5418 -284
rect -5366 -330 -5363 -284
rect -5171 -326 -5142 -250
rect -5418 -339 -5366 -333
rect -5171 -354 -5066 -326
rect -5650 -419 -5604 -386
rect -5650 -453 -5644 -419
rect -5610 -453 -5604 -419
rect -5650 -486 -5604 -453
rect -5492 -406 -5446 -386
rect -5342 -406 -5296 -386
rect -5184 -406 -5138 -386
rect -5492 -419 -5296 -406
rect -5492 -453 -5486 -419
rect -5452 -453 -5336 -419
rect -5302 -453 -5296 -419
rect -5492 -472 -5296 -453
rect -5190 -458 -5184 -406
rect -5132 -458 -5126 -406
rect -5492 -486 -5446 -472
rect -5342 -486 -5296 -472
rect -5184 -486 -5138 -458
rect -5644 -636 -5616 -486
rect -5488 -531 -5449 -486
rect -5494 -537 -5442 -531
rect -5494 -595 -5442 -589
rect -5094 -636 -5066 -354
rect -5020 -404 -4990 -219
rect -5037 -456 -5031 -404
rect -4979 -456 -4973 -404
rect -5644 -664 -5066 -636
rect -6429 -783 -5701 -744
rect -5020 -775 -4990 -456
rect -6429 -789 -6423 -783
<< via1 >>
rect -6270 93 -6218 102
rect -6206 93 -6154 102
rect -6142 93 -6090 102
rect -6078 93 -6026 102
rect -6014 93 -5962 102
rect -5950 93 -5898 102
rect -5886 93 -5834 102
rect -6270 59 -6249 93
rect -6249 59 -6218 93
rect -6206 59 -6177 93
rect -6177 59 -6154 93
rect -6142 59 -6105 93
rect -6105 59 -6090 93
rect -6078 59 -6071 93
rect -6071 59 -6033 93
rect -6033 59 -6026 93
rect -6014 59 -5999 93
rect -5999 59 -5962 93
rect -5950 59 -5927 93
rect -5927 59 -5898 93
rect -5886 59 -5855 93
rect -5855 59 -5834 93
rect -6270 50 -6218 59
rect -6206 50 -6154 59
rect -6142 50 -6090 59
rect -6078 50 -6026 59
rect -6014 50 -5962 59
rect -5950 50 -5898 59
rect -5886 50 -5834 59
rect -5754 -177 -5702 -125
rect -5030 -178 -4978 -126
rect -6485 -335 -6433 -283
rect -6070 -302 -6018 -292
rect -6070 -336 -6062 -302
rect -6062 -336 -6028 -302
rect -6028 -336 -6018 -302
rect -6070 -344 -6018 -336
rect -6290 -597 -6238 -588
rect -6226 -597 -6174 -588
rect -6290 -631 -6271 -597
rect -6271 -631 -6238 -597
rect -6226 -631 -6199 -597
rect -6199 -631 -6174 -597
rect -6290 -640 -6238 -631
rect -6226 -640 -6174 -631
rect -6162 -597 -6110 -588
rect -6162 -631 -6161 -597
rect -6161 -631 -6127 -597
rect -6127 -631 -6110 -597
rect -6162 -640 -6110 -631
rect -6098 -597 -6046 -588
rect -6098 -631 -6089 -597
rect -6089 -631 -6055 -597
rect -6055 -631 -6046 -597
rect -6098 -640 -6046 -631
rect -6034 -597 -5982 -588
rect -6034 -631 -6017 -597
rect -6017 -631 -5983 -597
rect -5983 -631 -5982 -597
rect -6034 -640 -5982 -631
rect -5970 -597 -5918 -588
rect -5906 -597 -5854 -588
rect -5970 -631 -5945 -597
rect -5945 -631 -5918 -597
rect -5906 -631 -5873 -597
rect -5873 -631 -5854 -597
rect -5970 -640 -5918 -631
rect -5906 -640 -5854 -631
rect -6481 -789 -6429 -737
rect -5418 -290 -5366 -281
rect -5418 -324 -5409 -290
rect -5409 -324 -5375 -290
rect -5375 -324 -5366 -290
rect -5418 -333 -5366 -324
rect -5184 -419 -5132 -406
rect -5184 -453 -5178 -419
rect -5178 -453 -5144 -419
rect -5144 -453 -5132 -419
rect -5184 -458 -5132 -453
rect -5494 -589 -5442 -537
rect -5031 -456 -4979 -404
<< metal2 >>
rect -6482 -277 -6441 237
rect -6322 104 -5782 146
rect -6322 48 -6280 104
rect -6224 102 -6200 104
rect -6144 102 -6120 104
rect -6064 102 -6040 104
rect -5984 102 -5960 104
rect -5904 102 -5880 104
rect -6218 50 -6206 102
rect -6144 50 -6142 102
rect -5962 50 -5960 102
rect -5898 50 -5886 102
rect -6224 48 -6200 50
rect -6144 48 -6120 50
rect -6064 48 -6040 50
rect -5984 48 -5960 50
rect -5904 48 -5880 50
rect -5824 48 -5782 104
rect -6322 6 -5782 48
rect -5755 -123 -5700 -117
rect -5030 -123 -4978 -120
rect -5755 -125 -4962 -123
rect -5755 -177 -5754 -125
rect -5702 -126 -4962 -125
rect -5702 -177 -5030 -126
rect -5755 -178 -5030 -177
rect -4978 -178 -4962 -126
rect -5755 -184 -5700 -178
rect -5030 -184 -4978 -178
rect -6485 -283 -6433 -277
rect -6070 -292 -6018 -286
rect -6485 -341 -6433 -335
rect -6071 -341 -6070 -298
rect -6482 -380 -6441 -341
rect -5424 -333 -5418 -281
rect -5366 -333 -5360 -281
rect -6070 -350 -6018 -344
rect -6067 -397 -6028 -350
rect -5409 -397 -5375 -333
rect -6067 -436 -5373 -397
rect -5184 -406 -5132 -400
rect -5031 -404 -4979 -398
rect -5132 -446 -5031 -417
rect -6482 -731 -6441 -460
rect -5184 -464 -5132 -458
rect -5031 -462 -4979 -456
rect -6342 -586 -5802 -544
rect -6342 -642 -6300 -586
rect -6244 -588 -6220 -586
rect -6164 -588 -6140 -586
rect -6084 -588 -6060 -586
rect -6004 -588 -5980 -586
rect -5924 -588 -5900 -586
rect -6238 -640 -6226 -588
rect -6164 -640 -6162 -588
rect -5982 -640 -5980 -588
rect -5918 -640 -5906 -588
rect -6244 -642 -6220 -640
rect -6164 -642 -6140 -640
rect -6084 -642 -6060 -640
rect -6004 -642 -5980 -640
rect -5924 -642 -5900 -640
rect -5844 -642 -5802 -586
rect -5500 -589 -5494 -537
rect -5442 -589 -5436 -537
rect -6342 -684 -5802 -642
rect -6482 -737 -6429 -731
rect -6482 -789 -6481 -737
rect -5487 -753 -5448 -589
rect -6482 -795 -6429 -789
rect -6482 -860 -6441 -795
<< via2 >>
rect -6280 102 -6224 104
rect -6200 102 -6144 104
rect -6120 102 -6064 104
rect -6040 102 -5984 104
rect -5960 102 -5904 104
rect -5880 102 -5824 104
rect -6280 50 -6270 102
rect -6270 50 -6224 102
rect -6200 50 -6154 102
rect -6154 50 -6144 102
rect -6120 50 -6090 102
rect -6090 50 -6078 102
rect -6078 50 -6064 102
rect -6040 50 -6026 102
rect -6026 50 -6014 102
rect -6014 50 -5984 102
rect -5960 50 -5950 102
rect -5950 50 -5904 102
rect -5880 50 -5834 102
rect -5834 50 -5824 102
rect -6280 48 -6224 50
rect -6200 48 -6144 50
rect -6120 48 -6064 50
rect -6040 48 -5984 50
rect -5960 48 -5904 50
rect -5880 48 -5824 50
rect -6300 -588 -6244 -586
rect -6220 -588 -6164 -586
rect -6140 -588 -6084 -586
rect -6060 -588 -6004 -586
rect -5980 -588 -5924 -586
rect -5900 -588 -5844 -586
rect -6300 -640 -6290 -588
rect -6290 -640 -6244 -588
rect -6220 -640 -6174 -588
rect -6174 -640 -6164 -588
rect -6140 -640 -6110 -588
rect -6110 -640 -6098 -588
rect -6098 -640 -6084 -588
rect -6060 -640 -6046 -588
rect -6046 -640 -6034 -588
rect -6034 -640 -6004 -588
rect -5980 -640 -5970 -588
rect -5970 -640 -5924 -588
rect -5900 -640 -5854 -588
rect -5854 -640 -5844 -588
rect -6300 -642 -6244 -640
rect -6220 -642 -6164 -640
rect -6140 -642 -6084 -640
rect -6060 -642 -6004 -640
rect -5980 -642 -5924 -640
rect -5900 -642 -5844 -640
<< metal3 >>
rect -6614 104 -4922 146
rect -6614 48 -6280 104
rect -6224 48 -6200 104
rect -6144 48 -6120 104
rect -6064 48 -6040 104
rect -5984 48 -5960 104
rect -5904 48 -5880 104
rect -5824 48 -4922 104
rect -6614 6 -4922 48
rect -6614 -586 -4922 -544
rect -6614 -642 -6300 -586
rect -6244 -642 -6220 -586
rect -6164 -642 -6140 -586
rect -6084 -642 -6060 -586
rect -6004 -642 -5980 -586
rect -5924 -642 -5900 -586
rect -5844 -642 -4922 -586
rect -6614 -684 -4922 -642
<< labels >>
flabel metal1 s -6442 -329 -6422 -290 7 FreeSans 600 0 0 0 DX
flabel metal1 s -6471 -783 -6443 -744 7 FreeSans 600 0 0 0 DX_BUF
flabel metal3 s -4952 6 -4922 146 3 FreeSans 600 0 0 0 VCC
flabel metal3 s -4952 -684 -4922 -544 3 FreeSans 600 0 0 0 VSS
flabel metal1 s -5488 170 -5449 195 3 FreeSans 600 0 0 0 VOUT
flabel metal2 s -5487 -753 -5448 -729 7 FreeSans 600 0 0 0 VOUT
flabel metal1 s -6132 -354 -6132 -354 7 FreeSans 600 0 0 0 DX_
flabel metal3 s -6614 -684 -6584 -544 7 FreeSans 600 0 0 0 VSS
flabel metal3 s -6614 6 -6584 146 7 FreeSans 600 0 0 0 VCC
flabel metal1 s -5158 203 -5158 203 1 FreeSans 480 0 0 40 VREFH
flabel metal1 s -5005 -763 -5005 -763 5 FreeSans 480 0 0 -40 VREFL
<< end >>
