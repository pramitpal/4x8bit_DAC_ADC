* SPICE3 file created from 4_bit_dac.ext - technology: sky130A

.subckt x4_bit_dac D0 VREFL D0_BUF VREFH D1 D1_BUF D2 D3 D2_BUF D3_BUF VOUT VSS VCC
X0 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H D0_BUF.t2 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VCC.t63 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t34 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 3_bit_dac_0[0].D0 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X3 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_2862# 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L VCC.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X4 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_4090# 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH VCC.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X5 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_1634# 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH VCC.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X6 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[0].2_bit_dac_0[1].VOUT VSS.t60 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[0].D1 VSS.t77 VSS.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_4090# 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X10 3_bit_dac_0[0].switch_n_3v3_1.DX_ switch_n_3v3_0.D2 VCC.t16 VCC.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X11 3_bit_dac_0[1].switch_n_3v3_1.DX_ D2.t0 VCC.t39 VCC.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X12 3_bit_dac_0[0].VOUT D2_BUF.t2 3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X13 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[1].2_bit_dac_0[0].D1 VCC.t19 VCC.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X14 D3_BUF.t0 switch_n_3v3_0.DX_ VSS.t11 VSS.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X15 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 3_bit_dac_0[1].VREFH VSS.t35 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X16 3_bit_dac_0[1].2_bit_dac_0[0].D1 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS.t38 VSS.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X17 a_1556_1634# 3_bit_dac_0[0].D0 VCC.t67 VCC.t66 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X18 a_1556_4090# D0.t0 VCC.t21 VCC.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X19 a_1556_4090# D0.t1 VSS.t43 VSS.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X20 3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[0].2_bit_dac_0[0].D1 VSS.t74 VSS.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X21 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS.t8 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X22 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t3 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X23 3_bit_dac_0[0].2_bit_dac_0[0].D0 a_1556_1634# VCC.t28 VCC.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X24 3_bit_dac_0[1].2_bit_dac_0[0].D0 a_1556_4090# VCC.t53 VCC.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X25 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 3_bit_dac_0[0].2_bit_dac_0[0].D0 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X26 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_406# 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L VCC.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X27 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_2862# 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X28 3_bit_dac_0[1].2_bit_dac_0[0].D0 a_1556_4090# VSS.t54 VSS.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X29 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS.t8 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X30 3_bit_dac_0[1].2_bit_dac_0[0].VOUT 3_bit_dac_0[0].D1 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X31 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS.t8 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X32 3_bit_dac_0[1].VOUT switch_n_3v3_0.DX_ VOUT.t1 VSS.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X33 switch_n_3v3_0.DX_ D3.t0 VSS.t45 VSS.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X34 D0_BUF.t0 a_1556_406# VSS.t25 VSS.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X35 a_1556_406# 3_bit_dac_0[0].2_bit_dac_0[0].D0 VSS.t14 VSS.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X36 3_bit_dac_0[1].2_bit_dac_0[1].VREFH 3_bit_dac_0[0].D0 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X37 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[1].2_bit_dac_0[1].VOUT VSS.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X38 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ D1.t0 VSS.t40 VSS.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X39 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t34 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X40 3_bit_dac_0[0].2_bit_dac_0[0].D1 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VCC.t58 VCC.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X41 3_bit_dac_0[1].2_bit_dac_0[0].D1 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VCC.t37 VCC.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X42 3_bit_dac_0[0].2_bit_dac_0[1].VOUT 3_bit_dac_0[0].2_bit_dac_0[0].D1 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X43 3_bit_dac_0[1].2_bit_dac_0[1].VOUT 3_bit_dac_0[1].2_bit_dac_0[0].D1 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X44 3_bit_dac_0[1].VOUT switch_n_3v3_0.D2 3_bit_dac_0[1].2_bit_dac_0[0].VOUT VSS.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X45 D2_BUF.t0 3_bit_dac_0[0].switch_n_3v3_1.DX_ VSS.t63 VSS.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X46 3_bit_dac_0[0].2_bit_dac_0[0].VOUT 3_bit_dac_0[0].switch_n_3v3_1.DX_ 3_bit_dac_0[0].VOUT VCC.t61 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X47 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t35 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X48 3_bit_dac_0[1].2_bit_dac_0[0].VOUT 3_bit_dac_0[1].switch_n_3v3_1.DX_ 3_bit_dac_0[1].VOUT VCC.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X49 3_bit_dac_0[0].2_bit_dac_0[0].VOUT D1_BUF.t2 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X50 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 3_bit_dac_0[0].2_bit_dac_0[0].D0 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VCC.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X51 a_1556_2862# 3_bit_dac_0[1].2_bit_dac_0[0].D0 VSS.t7 VSS.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X52 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 3_bit_dac_0[1].2_bit_dac_0[0].D0 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VCC.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X53 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[1].2_bit_dac_0[0].VOUT VCC.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X54 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t3 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X55 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_406# 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH VCC.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X56 D3_BUF.t1 switch_n_3v3_0.DX_ VCC.t9 VCC.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X57 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_1634# 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L VCC.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X58 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_4090# 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L VCC.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X59 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3_bit_dac_0[1].2_bit_dac_0[0].D0 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X60 D1_BUF.t0 3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS.t47 VSS.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X61 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L D0_BUF.t3 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X62 VOUT.t3 D3_BUF.t2 3_bit_dac_0[1].VOUT VCC.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X63 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH D0_BUF.t4 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X64 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_4090# VREFL.t2 VSS.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X65 3_bit_dac_0[0].D0 a_1556_2862# VSS.t32 VSS.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X66 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_1634# 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X67 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH VREFH.t0 VSS.t35 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X68 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 3_bit_dac_0[1].VREFH VSS.t34 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X69 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L VREFL.t1 VSS.t34 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X70 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[0].D1 VCC.t73 VCC.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X71 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ D1.t1 VCC.t48 VCC.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X72 3_bit_dac_0[0].2_bit_dac_0[1].VOUT 3_bit_dac_0[0].2_bit_dac_0[0].D1 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X73 3_bit_dac_0[0].2_bit_dac_0[1].VOUT 3_bit_dac_0[0].switch_n_3v3_1.DX_ 3_bit_dac_0[0].VOUT VSS.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X74 3_bit_dac_0[0].switch_n_3v3_1.DX_ switch_n_3v3_0.D2 VSS.t17 VSS.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X75 3_bit_dac_0[0].2_bit_dac_0[0].VOUT D1_BUF.t3 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X76 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_2862# 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH VCC.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X77 3_bit_dac_0[0].D1 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS.t51 VSS.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X78 switch_n_3v3_0.DX_ D3.t1 VCC.t50 VCC.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X79 a_1556_1634# 3_bit_dac_0[0].D0 VSS.t68 VSS.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X80 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 3_bit_dac_0[0].D0 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X81 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t3 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X82 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t35 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X83 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_2862# 3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X84 switch_n_3v3_0.D2 3_bit_dac_0[1].switch_n_3v3_1.DX_ VSS.t2 VSS.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X85 3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[0].2_bit_dac_0[0].D1 VCC.t69 VCC.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X86 a_1556_2862# 3_bit_dac_0[1].2_bit_dac_0[0].D0 VCC.t5 VCC.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X87 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS.t8 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X88 3_bit_dac_0[0].2_bit_dac_0[0].D0 a_1556_1634# VSS.t28 VSS.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X89 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_406# 3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X90 3_bit_dac_0[1].VREFH 3_bit_dac_0[0].2_bit_dac_0[0].D0 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X91 VREFL.t0 3_bit_dac_0[1].2_bit_dac_0[0].D0 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X92 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[1].2_bit_dac_0[0].VOUT VSS.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X93 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[1].2_bit_dac_0[0].D1 VSS.t21 VSS.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X94 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 3_bit_dac_0[1].2_bit_dac_0[0].D0 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X95 3_bit_dac_0[0].D0 a_1556_2862# VCC.t32 VCC.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X96 D0_BUF.t1 a_1556_406# VCC.t23 VCC.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X97 a_1556_406# 3_bit_dac_0[0].2_bit_dac_0[0].D0 VCC.t11 VCC.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X98 VOUT.t2 D3_BUF.t3 3_bit_dac_0[0].VOUT VSS.t56 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X99 3_bit_dac_0[0].2_bit_dac_0[0].D1 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS.t59 VSS.t58 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X100 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[0].2_bit_dac_0[1].VOUT VCC.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X101 3_bit_dac_0[1].2_bit_dac_0[1].VOUT 3_bit_dac_0[1].2_bit_dac_0[0].D1 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X102 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[1].2_bit_dac_0[1].VOUT VCC.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X103 3_bit_dac_0[1].2_bit_dac_0[1].VOUT 3_bit_dac_0[1].switch_n_3v3_1.DX_ 3_bit_dac_0[1].VOUT VSS.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X104 3_bit_dac_0[1].switch_n_3v3_1.DX_ D2.t1 VSS.t71 VSS.t70 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X105 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[0].2_bit_dac_0[0].VOUT VCC.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X106 D2_BUF.t1 3_bit_dac_0[0].switch_n_3v3_1.DX_ VCC.t60 VCC.t59 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X107 switch_n_3v3_0.D2 3_bit_dac_0[1].switch_n_3v3_1.DX_ VCC.t1 VCC.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X108 3_bit_dac_0[0].VOUT D2_BUF.t3 3_bit_dac_0[0].2_bit_dac_0[1].VOUT VCC.t55 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X109 3_bit_dac_0[1].VOUT switch_n_3v3_0.D2 3_bit_dac_0[1].2_bit_dac_0[1].VOUT VCC.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X110 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3_bit_dac_0[0].2_bit_dac_0[0].D0 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X111 3_bit_dac_0[0].D1 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VCC.t45 VCC.t44 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X112 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_406# 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X113 3_bit_dac_0[1].2_bit_dac_0[0].VOUT 3_bit_dac_0[0].D1 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t71 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X114 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_1634# 3_bit_dac_0[1].VREFH VSS.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X115 3_bit_dac_0[0].VOUT switch_n_3v3_0.DX_ VOUT.t0 VCC.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X116 D1_BUF.t1 3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VCC.t41 VCC.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X117 3_bit_dac_0[0].2_bit_dac_0[1].VREFH D0_BUF.t5 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X118 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t3 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X119 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 3_bit_dac_0[0].D0 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VCC.t64 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
C0 VREFL 3_bit_dac_0[0].D0 4.97e-19
C1 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3_bit_dac_0[1].2_bit_dac_0[1].VREFH 0.0124f
C2 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.39f
C3 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 3_bit_dac_0[0].D0 1.9e-19
C4 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 3_bit_dac_0[0].2_bit_dac_0[0].D0 0.265f
C5 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3_bit_dac_0[0].D1 0.176f
C6 D1 VCC 0.459f
C7 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.00819f
C8 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.0172f
C9 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 1.46e-19
C10 switch_n_3v3_0.D7 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 4.71e-19
C11 D0_BUF 3_bit_dac_0[0].2_bit_dac_0[0].D1 0.0179f
C12 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.0923f
C13 3_bit_dac_0[1].2_bit_dac_0[1].VREFH 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.0579f
C14 switch_n_3v3_0.DX_ VCC 0.712f
C15 3_bit_dac_0[0].2_bit_dac_0[0].VOUT 3_bit_dac_0[0].2_bit_dac_0[0].D1 0.00692f
C16 3_bit_dac_0[0].switch_n_3v3_1.DX_ 3_bit_dac_0[1].VOUT 3.68e-19
C17 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0102f
C18 3_bit_dac_0[0].D0 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.472f
C19 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[1].2_bit_dac_0[0].D1 0.219f
C20 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.0018f
C21 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.0261f
C22 3_bit_dac_0[1].switch_n_3v3_1.DX_ 3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.125f
C23 VOUT switch_n_3v3_0.D6 2.29e-20
C24 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.805f
C25 VCC 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.836f
C26 3_bit_dac_0[0].D1 switch_n_3v3_0.D6 1.79e-20
C27 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 3_bit_dac_0[0].2_bit_dac_0[1].VREFH 0.482f
C28 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3_bit_dac_0[0].2_bit_dac_0[0].D0 0.00349f
C29 a_1556_4090# D0 0.0975f
C30 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH a_1556_406# 0.175f
C31 VCC 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.312f
C32 switch_n_3v3_0.D2 3_bit_dac_0[1].VOUT 0.0744f
C33 3_bit_dac_0[0].2_bit_dac_0[0].VOUT D0_BUF 2.29e-20
C34 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.236f
C35 D1_BUF 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.176f
C36 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0172f
C37 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.0035f
C38 D1_BUF 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 4.15e-19
C39 3_bit_dac_0[1].switch_n_3v3_1.DX_ switch_n_3v3_0.D4 1.33e-19
C40 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.68e-19
C41 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D4 2.51e-19
C42 D3 3_bit_dac_0[1].VOUT 2.78e-19
C43 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0927f
C44 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3_bit_dac_0[0].2_bit_dac_0[0].D1 1.85e-19
C45 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 4.25e-19
C46 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.579f
C47 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 1.68e-19
C48 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3_bit_dac_0[0].D0 0.00164f
C49 D2_BUF 3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.177f
C50 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.00819f
C51 a_1556_4090# D1 0.003f
C52 3_bit_dac_0[0].2_bit_dac_0[0].D0 3_bit_dac_0[1].2_bit_dac_0[1].VREFH 4.97e-19
C53 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00163f
C54 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.511f
C55 3_bit_dac_0[0].2_bit_dac_0[0].D0 3_bit_dac_0[0].2_bit_dac_0[1].VOUT 2.29e-20
C56 D3_BUF D2_BUF 0.307f
C57 switch_n_3v3_0.D2 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.129f
C58 switch_n_3v3_0.D5 3_bit_dac_0[1].VOUT 3.23e-20
C59 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VCC 0.714f
C60 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 7.75e-19
C61 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3.82e-19
C62 switch_n_3v3_0.D6 3_bit_dac_0[0].2_bit_dac_0[0].D1 1.79e-20
C63 3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[0].2_bit_dac_0[0].D1 0.111f
C64 3_bit_dac_0[1].2_bit_dac_0[1].VOUT D1 0.0057f
C65 3_bit_dac_0[0].D0 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5.84e-19
C66 switch_n_3v3_0.D2 3_bit_dac_0[1].2_bit_dac_0[0].D1 0.0155f
C67 3_bit_dac_0[1].2_bit_dac_0[1].VOUT switch_n_3v3_0.DX_ 3.68e-19
C68 3_bit_dac_0[0].VOUT 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 2.49e-22
C69 a_1556_4090# 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.175f
C70 3_bit_dac_0[0].switch_n_3v3_1.DX_ 3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.125f
C71 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL D3 0.017f
C72 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 3.82e-19
C73 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3_bit_dac_0[1].2_bit_dac_0[0].D0 2.38e-19
C74 D3_BUF 3_bit_dac_0[0].switch_n_3v3_1.DX_ 3.74e-19
C75 VCC D2_BUF 0.337f
C76 3_bit_dac_0[1].2_bit_dac_0[0].D1 D3 3.11e-20
C77 3_bit_dac_0[1].2_bit_dac_0[1].VOUT 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 2.34e-21
C78 3_bit_dac_0[1].2_bit_dac_0[0].D0 3_bit_dac_0[1].2_bit_dac_0[0].D1 0.00262f
C79 a_1556_1634# 3_bit_dac_0[0].2_bit_dac_0[0].D0 0.325f
C80 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.39f
C81 a_1556_4090# 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.397f
C82 3_bit_dac_0[0].2_bit_dac_0[0].D0 VCC 1.17f
C83 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_2862# 0.0892f
C84 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.322f
C85 3_bit_dac_0[0].D0 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2.38e-19
C86 VOUT 3_bit_dac_0[1].VOUT 0.505f
C87 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH switch_n_3v3_0.D7 4.71e-19
C88 3_bit_dac_0[1].2_bit_dac_0[1].VOUT 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 3.62e-20
C89 D0_BUF 3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5.84e-19
C90 3_bit_dac_0[0].2_bit_dac_0[0].VOUT 3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.229f
C91 3_bit_dac_0[0].2_bit_dac_0[0].VOUT switch_n_3v3_0.D6 0.0199f
C92 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL switch_n_3v3_0.D5 0.00306f
C93 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 3_bit_dac_0[1].2_bit_dac_0[1].VREFH 0.005f
C94 VCC 3_bit_dac_0[0].switch_n_3v3_1.DX_ 0.698f
C95 VREFL D0 0.77f
C96 switch_n_3v3_0.D2 3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.613f
C97 D1 switch_n_3v3_0.D4 1.41e-21
C98 switch_n_3v3_0.D2 3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.14f
C99 3_bit_dac_0[1].2_bit_dac_0[0].D1 switch_n_3v3_0.D5 2.05e-20
C100 a_1556_406# D1_BUF 6.04e-19
C101 switch_n_3v3_0.DX_ switch_n_3v3_0.D4 1.33e-19
C102 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 8.92e-19
C103 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D7 1.45e-19
C104 3_bit_dac_0[0].D0 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.24f
C105 switch_n_3v3_0.D2 D3_BUF 0.631f
C106 3_bit_dac_0[0].2_bit_dac_0[1].VREFH a_1556_1634# 2.68e-20
C107 VREFH 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 7.62e-19
C108 3_bit_dac_0[0].2_bit_dac_0[1].VREFH VCC 0.132f
C109 D3 3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.0607f
C110 D3 3_bit_dac_0[0].2_bit_dac_0[1].VOUT 2.69e-19
C111 3_bit_dac_0[1].2_bit_dac_0[0].D0 3_bit_dac_0[1].2_bit_dac_0[1].VREFH 1.06f
C112 D0 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 1.9e-19
C113 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 3_bit_dac_0[0].D0 0.00349f
C114 a_1556_406# 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0892f
C115 D3_BUF D3 0.0618f
C116 a_1556_4090# 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 1.21e-20
C117 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 3_bit_dac_0[1].VREFH 0.005f
C118 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L a_1556_1634# 0.403f
C119 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L VCC 0.291f
C120 a_1556_406# 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00538f
C121 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH switch_n_3v3_0.D7 2.94e-20
C122 switch_n_3v3_0.D2 VCC 0.776f
C123 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3_bit_dac_0[0].D1 0.635f
C124 3_bit_dac_0[1].2_bit_dac_0[0].D0 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.315f
C125 switch_n_3v3_0.D7 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00143f
C126 3_bit_dac_0[1].2_bit_dac_0[1].VOUT 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.229f
C127 VREFL D1 1.7e-19
C128 3_bit_dac_0[1].2_bit_dac_0[0].D1 3_bit_dac_0[0].D1 0.044f
C129 D2 switch_n_3v3_0.D6 0.0325f
C130 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.189f
C131 switch_n_3v3_0.D5 3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.0259f
C132 switch_n_3v3_0.D5 3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.027f
C133 3_bit_dac_0[1].switch_n_3v3_1.DX_ 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 9.82e-21
C134 3_bit_dac_0[1].2_bit_dac_0[0].D1 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.00319f
C135 D3 VCC 0.331f
C136 3_bit_dac_0[1].2_bit_dac_0[0].D0 VCC 1.18f
C137 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 3_bit_dac_0[0].2_bit_dac_0[0].D0 0.24f
C138 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH switch_n_3v3_0.D6 6.67e-19
C139 D3_BUF switch_n_3v3_0.D5 0.0301f
C140 VREFL 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.201f
C141 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3_bit_dac_0[1].VREFH 3.38e-20
C142 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 3_bit_dac_0[0].2_bit_dac_0[0].D1 0.00319f
C143 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.0104f
C144 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ D1_BUF 6.11e-19
C145 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL switch_n_3v3_0.D7 0.00143f
C146 VREFL 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.138f
C147 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5.55e-20
C148 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H D1_BUF 0.00237f
C149 switch_n_3v3_0.D5 VCC 0.164f
C150 3_bit_dac_0[0].VOUT switch_n_3v3_0.D7 0.0133f
C151 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 3.82e-19
C152 VOUT 3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.00174f
C153 VOUT 3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.00583f
C154 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.322f
C155 D1_BUF 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.632f
C156 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D4 2.51e-19
C157 3_bit_dac_0[0].D1 3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.0757f
C158 3_bit_dac_0[0].D1 3_bit_dac_0[1].2_bit_dac_0[1].VREFH 3.54e-19
C159 3_bit_dac_0[0].D1 3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.0057f
C160 3_bit_dac_0[0].2_bit_dac_0[1].VREFH 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.0579f
C161 D3_BUF VOUT 0.0719f
C162 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.00143f
C163 D3_BUF 3_bit_dac_0[0].D1 4.43e-21
C164 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 3_bit_dac_0[1].2_bit_dac_0[1].VREFH 0.482f
C165 3_bit_dac_0[0].2_bit_dac_0[0].VOUT 3_bit_dac_0[1].VOUT 0.00117f
C166 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.128f
C167 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.00832f
C168 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3_bit_dac_0[0].2_bit_dac_0[0].D1 4.15e-19
C169 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.394f
C170 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.805f
C171 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.00832f
C172 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L D0_BUF 0.315f
C173 switch_n_3v3_0.D4 D2_BUF 0.0295f
C174 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 8.92e-19
C175 D2_BUF 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00476f
C176 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.579f
C177 3_bit_dac_0[1].2_bit_dac_0[1].VREFH 3_bit_dac_0[1].VREFH 0.0988f
C178 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0107f
C179 VOUT VCC 0.287f
C180 3_bit_dac_0[0].2_bit_dac_0[0].D0 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.347f
C181 3_bit_dac_0[0].D1 a_1556_1634# 0.003f
C182 3_bit_dac_0[0].D1 VCC 0.797f
C183 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3_bit_dac_0[0].D0 0.0824f
C184 switch_n_3v3_0.D2 3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.177f
C185 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH D1 0.0778f
C186 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L a_1556_1634# 1.29e-19
C187 a_1556_4090# 3_bit_dac_0[1].2_bit_dac_0[0].D0 0.325f
C188 3_bit_dac_0[1].2_bit_dac_0[0].D0 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.48e-19
C189 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L VCC 0.291f
C190 3_bit_dac_0[1].switch_n_3v3_1.DX_ 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00394f
C191 switch_n_3v3_0.D4 3_bit_dac_0[0].switch_n_3v3_1.DX_ 1.33e-19
C192 VREFH VCC 0.0022f
C193 3_bit_dac_0[0].switch_n_3v3_1.DX_ 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 9.82e-21
C194 3_bit_dac_0[1].2_bit_dac_0[1].VOUT D3 0.0236f
C195 3_bit_dac_0[1].2_bit_dac_0[1].VOUT 3_bit_dac_0[1].2_bit_dac_0[0].D0 2.29e-20
C196 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 3_bit_dac_0[0].D0 1.48e-19
C197 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.236f
C198 D2 3_bit_dac_0[1].VOUT 1.75e-20
C199 switch_n_3v3_0.DX_ 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 1.79e-20
C200 a_1556_1634# 3_bit_dac_0[1].VREFH 0.337f
C201 VCC 3_bit_dac_0[1].VREFH 0.14f
C202 3_bit_dac_0[0].2_bit_dac_0[0].D1 3_bit_dac_0[1].2_bit_dac_0[0].VOUT 1.81e-20
C203 3_bit_dac_0[0].2_bit_dac_0[0].D1 3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.0757f
C204 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_2862# 0.296f
C205 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 3_bit_dac_0[0].2_bit_dac_0[0].D0 0.0824f
C206 D0 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.48e-19
C207 D3_BUF 3_bit_dac_0[0].2_bit_dac_0[0].D1 2.79e-20
C208 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.394f
C209 3_bit_dac_0[1].2_bit_dac_0[0].D1 a_1556_2862# 0.003f
C210 a_1556_406# 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 9.57e-20
C211 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0018f
C212 3_bit_dac_0[1].2_bit_dac_0[1].VOUT switch_n_3v3_0.D5 0.0234f
C213 switch_n_3v3_0.D2 switch_n_3v3_0.D4 0.084f
C214 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL D0 8.97e-20
C215 switch_n_3v3_0.D2 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00872f
C216 3_bit_dac_0[0].2_bit_dac_0[0].D0 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.00105f
C217 switch_n_3v3_0.D6 3_bit_dac_0[1].VOUT 4.36e-20
C218 a_1556_1634# 3_bit_dac_0[0].2_bit_dac_0[0].D1 6.04e-19
C219 VCC 3_bit_dac_0[0].2_bit_dac_0[0].D1 0.793f
C220 3_bit_dac_0[1].switch_n_3v3_1.DX_ switch_n_3v3_0.D7 0.0268f
C221 D3 switch_n_3v3_0.D4 1.02f
C222 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D7 1.45e-19
C223 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 4.25e-19
C224 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H a_1556_406# 0.397f
C225 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 3_bit_dac_0[0].2_bit_dac_0[1].VREFH 0.205f
C226 3_bit_dac_0[0].2_bit_dac_0[0].VOUT 3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.349f
C227 3_bit_dac_0[1].2_bit_dac_0[0].D1 D2 0.0026f
C228 3_bit_dac_0[0].D1 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.037f
C229 a_1556_406# 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.296f
C230 3_bit_dac_0[0].2_bit_dac_0[0].VOUT D3_BUF 0.0201f
C231 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.579f
C232 3_bit_dac_0[1].2_bit_dac_0[1].VOUT VOUT 0.0157f
C233 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.00368f
C234 a_1556_2862# 3_bit_dac_0[1].2_bit_dac_0[1].VREFH 0.337f
C235 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3_bit_dac_0[1].2_bit_dac_0[0].D1 0.0801f
C236 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.00577f
C237 3_bit_dac_0[1].2_bit_dac_0[1].VOUT 3_bit_dac_0[0].D1 1.81e-20
C238 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.0927f
C239 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL D1 0.007f
C240 switch_n_3v3_0.D4 switch_n_3v3_0.D5 1.92f
C241 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.0018f
C242 switch_n_3v3_0.D5 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 8.21e-19
C243 switch_n_3v3_0.DX_ 3_bit_dac_0[0].VOUT 0.0858f
C244 a_1556_2862# 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 1.29e-19
C245 a_1556_1634# D0_BUF 0.00365f
C246 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 3_bit_dac_0[1].VREFH 0.138f
C247 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL switch_n_3v3_0.D6 0.00202f
C248 D0_BUF VCC 0.732f
C249 3_bit_dac_0[0].2_bit_dac_0[0].VOUT VCC 0.379f
C250 VREFL 3_bit_dac_0[1].2_bit_dac_0[0].D0 0.544f
C251 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.0104f
C252 3_bit_dac_0[1].2_bit_dac_0[0].D1 switch_n_3v3_0.D6 1.79e-20
C253 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.322f
C254 3_bit_dac_0[0].D0 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.00105f
C255 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.0261f
C256 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5.89e-20
C257 D2 3_bit_dac_0[1].2_bit_dac_0[0].VOUT 2.96e-19
C258 a_1556_2862# a_1556_1634# 0.00981f
C259 a_1556_2862# VCC 0.713f
C260 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.0018f
C261 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.115f
C262 3_bit_dac_0[0].D0 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.00379f
C263 3_bit_dac_0[1].2_bit_dac_0[0].D0 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0824f
C264 VOUT switch_n_3v3_0.D4 1.74e-20
C265 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.504f
C266 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.00114f
C267 3_bit_dac_0[0].D1 switch_n_3v3_0.D4 2.52e-20
C268 3_bit_dac_0[0].D1 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0801f
C269 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 3_bit_dac_0[0].2_bit_dac_0[0].D1 0.00237f
C270 D3_BUF 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 2.09e-21
C271 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.0172f
C272 switch_n_3v3_0.DX_ switch_n_3v3_0.D7 0.0268f
C273 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.115f
C274 switch_n_3v3_0.D6 3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.0258f
C275 D2 VCC 0.333f
C276 3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[0].2_bit_dac_0[1].VOUT 1.06e-19
C277 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH D2_BUF 1.98e-19
C278 switch_n_3v3_0.D6 3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.027f
C279 D2_BUF 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0668f
C280 3_bit_dac_0[0].2_bit_dac_0[0].D0 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3.36e-19
C281 3_bit_dac_0[0].2_bit_dac_0[0].D0 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.38f
C282 D3_BUF switch_n_3v3_0.D6 0.0299f
C283 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VCC 0.622f
C284 3_bit_dac_0[0].2_bit_dac_0[1].VREFH D1_BUF 3.54e-19
C285 switch_n_3v3_0.D2 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00476f
C286 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.128f
C287 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H D0_BUF 0.00379f
C288 VREFL 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.005f
C289 3_bit_dac_0[0].switch_n_3v3_1.DX_ 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00394f
C290 3_bit_dac_0[0].2_bit_dac_0[0].D0 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.00379f
C291 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH VREFH 0.0124f
C292 switch_n_3v3_0.D6 VCC 0.169f
C293 3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VCC 0.697f
C294 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH D3 0.00189f
C295 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3_bit_dac_0[1].2_bit_dac_0[0].D0 0.347f
C296 switch_n_3v3_0.D2 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.0211f
C297 3_bit_dac_0[0].D1 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.00375f
C298 a_1556_4090# a_1556_2862# 0.00981f
C299 a_1556_2862# 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 4.09e-19
C300 switch_n_3v3_0.D4 3_bit_dac_0[0].2_bit_dac_0[0].D1 2.38e-20
C301 3_bit_dac_0[0].VOUT D2_BUF 0.0719f
C302 3_bit_dac_0[0].2_bit_dac_0[1].VREFH 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 3.38e-20
C303 3_bit_dac_0[0].2_bit_dac_0[0].D1 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.176f
C304 3_bit_dac_0[0].D0 3_bit_dac_0[0].2_bit_dac_0[0].D0 0.132f
C305 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0923f
C306 3_bit_dac_0[1].switch_n_3v3_1.DX_ switch_n_3v3_0.DX_ 0.0104f
C307 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 3_bit_dac_0[1].VREFH 0.0551f
C308 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ D3 0.00594f
C309 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.189f
C310 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH switch_n_3v3_0.D5 8.21e-19
C311 switch_n_3v3_0.D2 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0701f
C312 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 3_bit_dac_0[1].VREFH 0.0124f
C313 3_bit_dac_0[0].VOUT 3_bit_dac_0[0].switch_n_3v3_1.DX_ 0.236f
C314 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D7 1.45e-19
C315 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D5 2.07e-19
C316 3_bit_dac_0[0].D0 3_bit_dac_0[0].2_bit_dac_0[1].VREFH 0.0104f
C317 3_bit_dac_0[0].2_bit_dac_0[0].VOUT switch_n_3v3_0.D4 0.02f
C318 D0_BUF 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00164f
C319 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.68e-19
C320 3_bit_dac_0[1].2_bit_dac_0[1].VOUT D2 0.134f
C321 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 3_bit_dac_0[0].2_bit_dac_0[0].D1 0.00491f
C322 3_bit_dac_0[0].2_bit_dac_0[0].VOUT 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00114f
C323 a_1556_406# 3_bit_dac_0[0].2_bit_dac_0[0].D0 0.0981f
C324 switch_n_3v3_0.D7 D2_BUF 0.0399f
C325 3_bit_dac_0[1].2_bit_dac_0[1].VOUT 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 6.14e-19
C326 3_bit_dac_0[0].D0 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.265f
C327 3_bit_dac_0[1].VOUT 3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.463f
C328 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3_bit_dac_0[1].2_bit_dac_0[0].D1 0.00805f
C329 switch_n_3v3_0.D2 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0668f
C330 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3_bit_dac_0[0].D1 1.85e-19
C331 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH D0 0.0572f
C332 3_bit_dac_0[0].2_bit_dac_0[1].VOUT 3_bit_dac_0[1].VOUT 0.0129f
C333 switch_n_3v3_0.D2 3_bit_dac_0[0].VOUT 1.85e-20
C334 3_bit_dac_0[1].2_bit_dac_0[0].D0 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.13f
C335 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH switch_n_3v3_0.D5 5.19e-20
C336 D3_BUF 3_bit_dac_0[1].VOUT 0.15f
C337 switch_n_3v3_0.D5 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00306f
C338 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL D3 0.0269f
C339 switch_n_3v3_0.D7 3_bit_dac_0[0].switch_n_3v3_1.DX_ 0.0268f
C340 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H D0 0.117f
C341 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[0].D1 0.219f
C342 3_bit_dac_0[1].2_bit_dac_0[1].VOUT switch_n_3v3_0.D6 0.0234f
C343 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 3_bit_dac_0[1].2_bit_dac_0[0].D0 0.38f
C344 3_bit_dac_0[1].2_bit_dac_0[0].D0 3_bit_dac_0[0].D0 0.132f
C345 3_bit_dac_0[0].VOUT D3 1.26e-20
C346 a_1556_406# 3_bit_dac_0[0].2_bit_dac_0[1].VREFH 0.337f
C347 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH D0_BUF 0.472f
C348 3_bit_dac_0[0].2_bit_dac_0[0].VOUT 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 2.34e-21
C349 3_bit_dac_0[1].switch_n_3v3_1.DX_ 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 1.79e-20
C350 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 4.25e-19
C351 D2 switch_n_3v3_0.D4 0.0322f
C352 VCC 3_bit_dac_0[1].VOUT 0.525f
C353 VREFL a_1556_2862# 1.97e-19
C354 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3_bit_dac_0[0].2_bit_dac_0[0].D0 0.472f
C355 a_1556_406# 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 1.29e-19
C356 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH switch_n_3v3_0.D4 0.00127f
C357 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L VCC 0.29f
C358 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.302f
C359 D1 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.00491f
C360 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00123f
C361 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3_bit_dac_0[1].2_bit_dac_0[1].VREFH 0.404f
C362 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.045f
C363 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL switch_n_3v3_0.D5 0.00306f
C364 3_bit_dac_0[0].D1 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3.53e-19
C365 3_bit_dac_0[1].2_bit_dac_0[0].D1 3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.00692f
C366 3_bit_dac_0[1].2_bit_dac_0[0].D1 3_bit_dac_0[1].2_bit_dac_0[1].VREFH 1.7e-19
C367 3_bit_dac_0[0].D1 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00805f
C368 3_bit_dac_0[0].VOUT switch_n_3v3_0.D5 3.8e-20
C369 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ D2_BUF 0.00132f
C370 D3_BUF 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.0204f
C371 switch_n_3v3_0.D2 switch_n_3v3_0.D7 0.0916f
C372 a_1556_2862# 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.175f
C373 3_bit_dac_0[0].2_bit_dac_0[0].D0 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5.84e-19
C374 D1 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.037f
C375 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 3_bit_dac_0[0].2_bit_dac_0[0].D0 0.13f
C376 3_bit_dac_0[1].2_bit_dac_0[0].D1 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 2.51e-20
C377 switch_n_3v3_0.D6 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 6.1e-19
C378 3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 1.46e-19
C379 D3 switch_n_3v3_0.D7 0.0518f
C380 3_bit_dac_0[0].D1 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.00237f
C381 3_bit_dac_0[0].2_bit_dac_0[0].D0 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 2.38e-19
C382 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_1634# 0.00538f
C383 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[0].switch_n_3v3_1.DX_ 1.79e-20
C384 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3_bit_dac_0[0].2_bit_dac_0[1].VREFH 0.0124f
C385 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 3_bit_dac_0[1].VREFH 0.404f
C386 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.39f
C387 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC 0.312f
C388 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.805f
C389 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[0].2_bit_dac_0[0].D1 6.11e-19
C390 3_bit_dac_0[1].2_bit_dac_0[0].D1 VCC 0.797f
C391 D1_BUF 3_bit_dac_0[0].2_bit_dac_0[0].D1 0.0392f
C392 VOUT 3_bit_dac_0[0].VOUT 0.301f
C393 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 3_bit_dac_0[0].D1 4.15e-19
C394 3_bit_dac_0[0].D0 3_bit_dac_0[0].D1 0.00262f
C395 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.0923f
C396 3_bit_dac_0[0].2_bit_dac_0[1].VOUT 3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.00805f
C397 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 3_bit_dac_0[0].D0 0.315f
C398 3_bit_dac_0[1].VREFH 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.0579f
C399 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 3_bit_dac_0[0].2_bit_dac_0[1].VREFH 0.138f
C400 D3_BUF 3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.00505f
C401 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.236f
C402 D3_BUF 3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.249f
C403 D1 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.111f
C404 3_bit_dac_0[0].2_bit_dac_0[1].VREFH 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.404f
C405 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 4.25e-19
C406 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5.89e-20
C407 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3_bit_dac_0[0].2_bit_dac_0[0].D1 0.0801f
C408 3_bit_dac_0[1].switch_n_3v3_1.DX_ switch_n_3v3_0.D2 0.219f
C409 3_bit_dac_0[1].2_bit_dac_0[1].VREFH 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.00183f
C410 switch_n_3v3_0.D2 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.0222f
C411 3_bit_dac_0[0].2_bit_dac_0[0].D1 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.635f
C412 3_bit_dac_0[0].D0 3_bit_dac_0[1].VREFH 1.06f
C413 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3_bit_dac_0[1].2_bit_dac_0[0].D0 1.9e-19
C414 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.00368f
C415 3_bit_dac_0[1].2_bit_dac_0[1].VOUT 3_bit_dac_0[1].VOUT 0.552f
C416 D0_BUF D1_BUF 0.00262f
C417 3_bit_dac_0[0].2_bit_dac_0[0].VOUT D1_BUF 0.0757f
C418 VCC 3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.529f
C419 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5.89e-20
C420 a_1556_1634# 3_bit_dac_0[1].2_bit_dac_0[1].VREFH 1.97e-19
C421 3_bit_dac_0[1].switch_n_3v3_1.DX_ D3 1.03e-19
C422 VCC 3_bit_dac_0[1].2_bit_dac_0[1].VREFH 0.143f
C423 VCC 3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.77f
C424 switch_n_3v3_0.DX_ D2_BUF 6.07e-19
C425 VOUT switch_n_3v3_0.D7 0.00687f
C426 D3_BUF VCC 0.396f
C427 a_1556_2862# 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 1.21e-20
C428 3_bit_dac_0[0].D1 switch_n_3v3_0.D7 1.57e-20
C429 VREFH a_1556_406# 2.68e-20
C430 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.00819f
C431 VCC 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.291f
C432 D0_BUF 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.347f
C433 3_bit_dac_0[0].2_bit_dac_0[0].VOUT 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.504f
C434 D0_BUF 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00349f
C435 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_4090# 2.93e-19
C436 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 8.92e-19
C437 3_bit_dac_0[0].2_bit_dac_0[0].VOUT 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.051f
C438 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH D2 0.00872f
C439 switch_n_3v3_0.DX_ 3_bit_dac_0[0].switch_n_3v3_1.DX_ 0.0104f
C440 3_bit_dac_0[1].switch_n_3v3_1.DX_ switch_n_3v3_0.D5 1.8e-19
C441 a_1556_4090# 3_bit_dac_0[1].2_bit_dac_0[0].D1 6.04e-19
C442 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D5 2.07e-19
C443 a_1556_406# 3_bit_dac_0[1].VREFH 1.97e-19
C444 a_1556_1634# VCC 0.713f
C445 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.00123f
C446 3_bit_dac_0[1].2_bit_dac_0[1].VOUT 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00473f
C447 switch_n_3v3_0.D4 3_bit_dac_0[1].VOUT 2.38e-20
C448 a_1556_2862# 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2.93e-19
C449 3_bit_dac_0[1].2_bit_dac_0[0].D0 D0 0.0255f
C450 3_bit_dac_0[1].2_bit_dac_0[1].VOUT 3_bit_dac_0[1].2_bit_dac_0[0].D1 0.0757f
C451 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3_bit_dac_0[0].D1 0.00491f
C452 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.0927f
C453 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH switch_n_3v3_0.D6 6.1e-19
C454 switch_n_3v3_0.D2 D1 1.48e-19
C455 switch_n_3v3_0.D2 switch_n_3v3_0.DX_ 3.53e-19
C456 a_1556_2862# 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.397f
C457 3_bit_dac_0[1].switch_n_3v3_1.DX_ VOUT 5.16e-19
C458 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.00577f
C459 3_bit_dac_0[0].2_bit_dac_0[0].VOUT 3_bit_dac_0[0].VOUT 0.314f
C460 a_1556_406# 3_bit_dac_0[0].2_bit_dac_0[0].D1 0.003f
C461 3_bit_dac_0[0].D1 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.111f
C462 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 3_bit_dac_0[1].2_bit_dac_0[1].VREFH 3.7e-20
C463 a_1556_4090# 3_bit_dac_0[1].2_bit_dac_0[1].VREFH 2.68e-20
C464 switch_n_3v3_0.D7 3_bit_dac_0[0].2_bit_dac_0[0].D1 1.57e-20
C465 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 3_bit_dac_0[0].2_bit_dac_0[1].VOUT 3.62e-20
C466 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_2862# 0.00538f
C467 D1 D3 2.93e-21
C468 a_1556_2862# 3_bit_dac_0[0].D0 0.325f
C469 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D6 1.72e-19
C470 3_bit_dac_0[1].2_bit_dac_0[0].D0 D1 0.0179f
C471 3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ D1_BUF 0.219f
C472 switch_n_3v3_0.DX_ D3 0.0904f
C473 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL switch_n_3v3_0.D4 0.00517f
C474 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3_bit_dac_0[1].VREFH 0.205f
C475 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00163f
C476 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.511f
C477 3_bit_dac_0[1].2_bit_dac_0[1].VOUT 3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.349f
C478 3_bit_dac_0[1].2_bit_dac_0[0].D1 switch_n_3v3_0.D4 2.52e-20
C479 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.0923f
C480 VREFH 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.0579f
C481 3_bit_dac_0[1].2_bit_dac_0[0].D1 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3.53e-19
C482 a_1556_4090# 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.403f
C483 3_bit_dac_0[1].2_bit_dac_0[0].D0 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.472f
C484 3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0927f
C485 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH switch_n_3v3_0.D6 3.83e-20
C486 a_1556_406# D0_BUF 0.325f
C487 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 3_bit_dac_0[1].VREFH 3.7e-20
C488 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.394f
C489 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H a_1556_1634# 0.397f
C490 a_1556_4090# VCC 0.713f
C491 3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 7.75e-19
C492 switch_n_3v3_0.DX_ switch_n_3v3_0.D5 1.8e-19
C493 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H VCC 0.312f
C494 switch_n_3v3_0.D6 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00202f
C495 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL D2 0.0701f
C496 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L D0 9.68e-20
C497 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3_bit_dac_0[1].VREFH 2.66e-20
C498 3_bit_dac_0[0].2_bit_dac_0[0].VOUT switch_n_3v3_0.D7 0.0265f
C499 3_bit_dac_0[1].2_bit_dac_0[0].D0 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.24f
C500 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3_bit_dac_0[0].2_bit_dac_0[0].D1 0.00375f
C501 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.511f
C502 VREFL 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 2.66e-20
C503 3_bit_dac_0[1].2_bit_dac_0[1].VOUT VCC 0.771f
C504 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3_bit_dac_0[0].D0 0.347f
C505 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3_bit_dac_0[0].VOUT 2.78e-22
C506 VREFL 3_bit_dac_0[1].2_bit_dac_0[0].D1 3.54e-19
C507 3_bit_dac_0[0].switch_n_3v3_1.DX_ D2_BUF 0.219f
C508 switch_n_3v3_0.D4 3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.0259f
C509 switch_n_3v3_0.D4 3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.0271f
C510 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3_bit_dac_0[1].2_bit_dac_0[0].VOUT 6.14e-19
C511 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[0].2_bit_dac_0[0].D1 0.219f
C512 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.514f
C513 D3_BUF switch_n_3v3_0.D4 0.929f
C514 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.322f
C515 switch_n_3v3_0.DX_ VOUT 0.236f
C516 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 3_bit_dac_0[0].2_bit_dac_0[0].D1 0.037f
C517 D3_BUF 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00189f
C518 switch_n_3v3_0.D2 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.00132f
C519 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL switch_n_3v3_0.D6 0.00202f
C520 3_bit_dac_0[1].2_bit_dac_0[0].D1 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.00491f
C521 switch_n_3v3_0.DX_ 3_bit_dac_0[0].D1 1.34e-20
C522 3_bit_dac_0[0].2_bit_dac_0[1].VREFH 3_bit_dac_0[0].2_bit_dac_0[0].D0 1.06f
C523 3_bit_dac_0[0].VOUT switch_n_3v3_0.D6 4.32e-20
C524 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3_bit_dac_0[0].2_bit_dac_0[0].D1 0.00805f
C525 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH D0_BUF 0.00105f
C526 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ D3 0.00213f
C527 3_bit_dac_0[1].2_bit_dac_0[0].D0 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5.84e-19
C528 D2 switch_n_3v3_0.D7 0.0518f
C529 switch_n_3v3_0.D2 D2_BUF 0.0694f
C530 switch_n_3v3_0.D4 VCC 0.161f
C531 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 3_bit_dac_0[0].2_bit_dac_0[0].D0 0.315f
C532 a_1556_1634# 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0892f
C533 VCC 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.622f
C534 VREFL 3_bit_dac_0[1].2_bit_dac_0[1].VREFH 0.0988f
C535 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH a_1556_2862# 0.0331f
C536 3_bit_dac_0[0].2_bit_dac_0[0].VOUT 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.0035f
C537 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH switch_n_3v3_0.D7 5.14e-19
C538 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H D0_BUF 0.24f
C539 3_bit_dac_0[0].2_bit_dac_0[0].VOUT 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 3.62e-20
C540 VREFL 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.482f
C541 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D5 2.07e-19
C542 D0_BUF 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.38f
C543 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L D1_BUF 2.51e-20
C544 switch_n_3v3_0.D2 3_bit_dac_0[0].switch_n_3v3_1.DX_ 0.0904f
C545 a_1556_406# 3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 1.21e-20
C546 3_bit_dac_0[0].2_bit_dac_0[0].VOUT 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.302f
C547 3_bit_dac_0[1].2_bit_dac_0[0].VOUT 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 2.34e-21
C548 3_bit_dac_0[1].2_bit_dac_0[1].VREFH 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.205f
C549 switch_n_3v3_0.D6 switch_n_3v3_0.D7 1.92f
C550 3_bit_dac_0[0].2_bit_dac_0[1].VREFH 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.00183f
C551 VREFL VCC 0.144f
C552 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00163f
C553 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.00577f
C554 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH a_1556_1634# 0.0331f
C555 switch_n_3v3_0.D5 D2_BUF 0.0293f
C556 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH VCC 0.835f
C557 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3_bit_dac_0[1].2_bit_dac_0[0].D1 0.176f
C558 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0018f
C559 3_bit_dac_0[1].switch_n_3v3_1.DX_ D2 0.0904f
C560 a_1556_1634# 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 9.57e-20
C561 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.128f
C562 VCC 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.836f
C563 3_bit_dac_0[1].2_bit_dac_0[0].D1 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.111f
C564 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[0].D1 6.11e-19
C565 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 1.46e-19
C566 switch_n_3v3_0.D5 3_bit_dac_0[0].switch_n_3v3_1.DX_ 1.8e-19
C567 3_bit_dac_0[1].2_bit_dac_0[0].D0 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 9.68e-20
C568 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.394f
C569 switch_n_3v3_0.D2 D3 0.628f
C570 VOUT D2_BUF 1.79e-20
C571 3_bit_dac_0[0].D1 D2_BUF 1.48e-19
C572 3_bit_dac_0[0].VOUT 3_bit_dac_0[1].VOUT 0.359f
C573 3_bit_dac_0[1].2_bit_dac_0[1].VOUT switch_n_3v3_0.D4 0.0234f
C574 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.00114f
C575 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0102f
C576 3_bit_dac_0[1].switch_n_3v3_1.DX_ switch_n_3v3_0.D6 2.54e-19
C577 3_bit_dac_0[0].D1 3_bit_dac_0[0].2_bit_dac_0[0].D0 0.0179f
C578 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 3_bit_dac_0[0].D0 9.68e-20
C579 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D6 1.72e-19
C580 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.0104f
C581 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 3_bit_dac_0[0].2_bit_dac_0[0].D0 1.9e-19
C582 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.00819f
C583 VREFH 3_bit_dac_0[0].2_bit_dac_0[0].D0 0.0104f
C584 VOUT 3_bit_dac_0[0].switch_n_3v3_1.DX_ 1.05e-19
C585 switch_n_3v3_0.D2 switch_n_3v3_0.D5 0.0616f
C586 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.0018f
C587 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.229f
C588 3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.128f
C589 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.0035f
C590 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.115f
C591 D1_BUF 3_bit_dac_0[0].2_bit_dac_0[1].VOUT 1.81e-20
C592 VREFL a_1556_4090# 0.337f
C593 3_bit_dac_0[1].2_bit_dac_0[0].D1 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.037f
C594 3_bit_dac_0[0].2_bit_dac_0[0].D0 3_bit_dac_0[1].VREFH 0.544f
C595 D3_BUF 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 8.04e-20
C596 a_1556_2862# 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 9.57e-20
C597 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.00832f
C598 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VCC 0.622f
C599 D3 switch_n_3v3_0.D5 0.0324f
C600 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.0107f
C601 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3_bit_dac_0[0].D0 0.38f
C602 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 3_bit_dac_0[1].2_bit_dac_0[0].D1 0.635f
C603 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3_bit_dac_0[0].VOUT 3.47e-20
C604 3_bit_dac_0[1].2_bit_dac_0[0].D1 3_bit_dac_0[0].D0 0.0179f
C605 D1 D2 0.00881f
C606 a_1556_2862# 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 4.83e-19
C607 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L a_1556_406# 0.403f
C608 a_1556_4090# 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0331f
C609 switch_n_3v3_0.D7 3_bit_dac_0[1].VOUT 0.0191f
C610 switch_n_3v3_0.D4 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00116f
C611 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3_bit_dac_0[0].2_bit_dac_0[1].VOUT 6.14e-19
C612 VREFH 3_bit_dac_0[0].2_bit_dac_0[1].VREFH 0.0988f
C613 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0018f
C614 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.00473f
C615 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.303f
C616 3_bit_dac_0[1].2_bit_dac_0[1].VREFH 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2.66e-20
C617 switch_n_3v3_0.D2 VOUT 1.25e-20
C618 3_bit_dac_0[0].D1 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.00319f
C619 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VCC 0.714f
C620 D1_BUF VCC 0.317f
C621 D3_BUF 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 1.15e-19
C622 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH D1 3.53e-19
C623 switch_n_3v3_0.D2 3_bit_dac_0[0].D1 0.0189f
C624 switch_n_3v3_0.DX_ 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 9.82e-21
C625 D3_BUF 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0269f
C626 3_bit_dac_0[0].2_bit_dac_0[0].D1 D2_BUF 0.00779f
C627 3_bit_dac_0[0].2_bit_dac_0[1].VREFH 3_bit_dac_0[1].VREFH 0.0988f
C628 3_bit_dac_0[0].2_bit_dac_0[0].D0 3_bit_dac_0[0].2_bit_dac_0[0].D1 0.00262f
C629 VOUT D3 1.93e-20
C630 3_bit_dac_0[1].2_bit_dac_0[0].VOUT 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 3.62e-20
C631 3_bit_dac_0[1].2_bit_dac_0[1].VREFH 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.138f
C632 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5.55e-20
C633 3_bit_dac_0[0].D1 D3 4.81e-19
C634 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 3_bit_dac_0[1].VREFH 0.482f
C635 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VCC 0.603f
C636 switch_n_3v3_0.DX_ switch_n_3v3_0.D6 2.54e-19
C637 a_1556_1634# 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.296f
C638 VCC 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.312f
C639 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.051f
C640 3_bit_dac_0[0].2_bit_dac_0[0].D1 3_bit_dac_0[0].switch_n_3v3_1.DX_ 1.34e-20
C641 3_bit_dac_0[1].2_bit_dac_0[0].D0 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.265f
C642 3_bit_dac_0[0].D0 3_bit_dac_0[1].2_bit_dac_0[0].VOUT 2.29e-20
C643 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 3_bit_dac_0[1].2_bit_dac_0[1].VREFH 3.38e-20
C644 3_bit_dac_0[0].D0 3_bit_dac_0[1].2_bit_dac_0[1].VREFH 0.544f
C645 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.00368f
C646 3_bit_dac_0[0].VOUT 3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.00426f
C647 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL switch_n_3v3_0.D7 0.00143f
C648 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5.59e-19
C649 3_bit_dac_0[0].VOUT 3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.651f
C650 3_bit_dac_0[1].2_bit_dac_0[0].D1 switch_n_3v3_0.D7 1.57e-20
C651 VOUT switch_n_3v3_0.D5 1.99e-20
C652 D3_BUF 3_bit_dac_0[0].VOUT 0.177f
C653 3_bit_dac_0[0].2_bit_dac_0[0].VOUT D2_BUF 0.546f
C654 3_bit_dac_0[0].2_bit_dac_0[1].VREFH 3_bit_dac_0[0].2_bit_dac_0[0].D1 1.7e-19
C655 3_bit_dac_0[0].D1 switch_n_3v3_0.D5 2.05e-20
C656 3_bit_dac_0[1].switch_n_3v3_1.DX_ 3_bit_dac_0[1].VOUT 0.255f
C657 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.189f
C658 3_bit_dac_0[0].2_bit_dac_0[0].D0 D0_BUF 0.124f
C659 3_bit_dac_0[1].2_bit_dac_0[0].D0 3_bit_dac_0[1].VREFH 0.0104f
C660 3_bit_dac_0[0].D0 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 1.9e-19
C661 a_1556_1634# 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 4.83e-19
C662 VCC 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.312f
C663 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5.55e-20
C664 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_4090# 0.0892f
C665 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 3_bit_dac_0[0].2_bit_dac_0[0].D1 2.51e-20
C666 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC 0.312f
C667 a_1556_2862# 3_bit_dac_0[0].2_bit_dac_0[0].D0 0.00365f
C668 3_bit_dac_0[0].D0 a_1556_1634# 0.0981f
C669 switch_n_3v3_0.D2 3_bit_dac_0[0].2_bit_dac_0[0].D1 0.0026f
C670 3_bit_dac_0[0].D0 VCC 1.18f
C671 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.805f
C672 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.514f
C673 3_bit_dac_0[0].VOUT VCC 0.338f
C674 3_bit_dac_0[0].2_bit_dac_0[0].VOUT 3_bit_dac_0[0].switch_n_3v3_1.DX_ 0.088f
C675 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ D2 0.0222f
C676 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.189f
C677 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.0102f
C678 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.00143f
C679 3_bit_dac_0[0].2_bit_dac_0[1].VREFH D0_BUF 0.538f
C680 switch_n_3v3_0.D7 3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.0324f
C681 switch_n_3v3_0.D7 3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.0397f
C682 3_bit_dac_0[1].2_bit_dac_0[1].VOUT 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 1.06e-19
C683 VREFL 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0551f
C684 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 7.75e-19
C685 D3_BUF switch_n_3v3_0.D7 0.0405f
C686 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 3_bit_dac_0[0].D1 2.51e-20
C687 3_bit_dac_0[1].switch_n_3v3_1.DX_ 3_bit_dac_0[1].2_bit_dac_0[0].D1 1.34e-20
C688 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5.59e-19
C689 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L D0_BUF 1.9e-19
C690 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.115f
C691 3_bit_dac_0[0].2_bit_dac_0[0].VOUT switch_n_3v3_0.D2 2.96e-19
C692 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D6 1.72e-19
C693 a_1556_406# a_1556_1634# 0.00981f
C694 a_1556_406# VCC 0.706f
C695 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3_bit_dac_0[0].2_bit_dac_0[0].D0 0.00164f
C696 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH switch_n_3v3_0.D4 0.00116f
C697 switch_n_3v3_0.D5 3_bit_dac_0[0].2_bit_dac_0[0].D1 2.05e-20
C698 3_bit_dac_0[0].D1 3_bit_dac_0[1].VREFH 1.7e-19
C699 switch_n_3v3_0.D7 VCC 0.425f
C700 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 3_bit_dac_0[1].VREFH 0.00183f
C701 a_1556_4090# 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 4.09e-19
C702 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.0261f
C703 switch_n_3v3_0.DX_ 3_bit_dac_0[1].VOUT 0.125f
C704 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3_bit_dac_0[1].2_bit_dac_0[1].VREFH 0.0551f
C705 switch_n_3v3_0.D6 D2_BUF 0.0293f
C706 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3_bit_dac_0[0].2_bit_dac_0[1].VOUT 2.34e-21
C707 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D4 2.51e-19
C708 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00143f
C709 D1_BUF 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 1.85e-19
C710 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_4090# 0.296f
C711 a_1556_4090# 3_bit_dac_0[0].D0 0.00365f
C712 3_bit_dac_0[1].switch_n_3v3_1.DX_ 3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.088f
C713 3_bit_dac_0[1].2_bit_dac_0[0].D0 a_1556_2862# 0.0981f
C714 3_bit_dac_0[0].D0 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.13f
C715 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[1].2_bit_dac_0[0].VOUT 1.06e-19
C716 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.229f
C717 3_bit_dac_0[1].switch_n_3v3_1.DX_ D3_BUF 6.07e-19
C718 3_bit_dac_0[0].2_bit_dac_0[0].VOUT switch_n_3v3_0.D5 0.0199f
C719 3_bit_dac_0[0].D1 3_bit_dac_0[0].2_bit_dac_0[0].D1 0.044f
C720 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.303f
C721 D3_BUF 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.00213f
C722 switch_n_3v3_0.D6 3_bit_dac_0[0].switch_n_3v3_1.DX_ 2.54e-19
C723 switch_n_3v3_0.D2 D2 0.0694f
C724 3_bit_dac_0[1].2_bit_dac_0[1].VOUT 3_bit_dac_0[0].VOUT 0.00112f
C725 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH switch_n_3v3_0.D4 7.43e-20
C726 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH a_1556_1634# 0.175f
C727 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.00473f
C728 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00123f
C729 switch_n_3v3_0.D4 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00517f
C730 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH VCC 0.836f
C731 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.579f
C732 switch_n_3v3_0.D2 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0145f
C733 switch_n_3v3_0.DX_ 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00394f
C734 D2 D3 0.398f
C735 3_bit_dac_0[1].switch_n_3v3_1.DX_ VCC 0.712f
C736 D1 3_bit_dac_0[1].2_bit_dac_0[0].D1 0.0384f
C737 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH D1_BUF 0.00375f
C738 a_1556_1634# 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 1.21e-20
C739 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VCC 0.714f
C740 3_bit_dac_0[1].2_bit_dac_0[1].VREFH D0 0.00555f
C741 3_bit_dac_0[0].2_bit_dac_0[0].D1 3_bit_dac_0[1].VREFH 3.54e-19
C742 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH D3 0.00213f
C743 a_1556_406# 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 4.83e-19
C744 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H a_1556_1634# 4.09e-19
C745 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H VCC 0.307f
C746 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3_bit_dac_0[1].2_bit_dac_0[0].D0 3.36e-19
C747 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5.59e-19
C748 switch_n_3v3_0.D2 switch_n_3v3_0.D6 0.0618f
C749 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5.89e-20
C750 a_1556_1634# 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 2.93e-19
C751 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC 0.243f
C752 3_bit_dac_0[1].2_bit_dac_0[0].D1 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.00375f
C753 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L D0 0.253f
C754 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL switch_n_3v3_0.D4 0.00517f
C755 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.236f
C756 D2 switch_n_3v3_0.D5 0.0322f
C757 3_bit_dac_0[0].D0 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3.36e-19
C758 VREFH D0_BUF 0.281f
C759 3_bit_dac_0[0].VOUT switch_n_3v3_0.D4 2.45e-20
C760 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0102f
C761 a_1556_2862# 3_bit_dac_0[0].D1 6.04e-19
C762 3_bit_dac_0[1].2_bit_dac_0[1].VOUT switch_n_3v3_0.D7 0.036f
C763 D3 switch_n_3v3_0.D6 0.0326f
C764 3_bit_dac_0[1].2_bit_dac_0[0].D1 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.00237f
C765 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH switch_n_3v3_0.D5 8.97e-19
C766 VCC D0 0.407f
C767 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L a_1556_2862# 0.403f
C768 D0_BUF 3_bit_dac_0[1].VREFH 4.97e-19
C769 switch_n_3v3_0.DX_ 3_bit_dac_0[1].2_bit_dac_0[0].VOUT 7.51e-19
C770 switch_n_3v3_0.DX_ 3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.0199f
C771 VREFL 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 3.7e-20
C772 switch_n_3v3_0.DX_ D3_BUF 0.219f
C773 a_1556_2862# 3_bit_dac_0[1].VREFH 2.68e-20
C774 switch_n_3v3_0.D5 switch_n_3v3_0.D6 1.92f
C775 D1 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.00319f
C776 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VREFL 0.404f
C777 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.39f
R0 D0_BUF.n15 D0_BUF.n0 400.238
R1 D0_BUF.n3 D0_BUF.n2 292.5
R2 D0_BUF.n17 D0_BUF.n16 153.333
R3 D0_BUF D0_BUF.n17 105.805
R4 D0_BUF.n0 D0_BUF.t2 83.8685
R5 D0_BUF.n16 D0_BUF.t5 80.9765
R6 D0_BUF.n16 D0_BUF.t3 57.8405
R7 D0_BUF.n0 D0_BUF.t4 54.9485
R8 D0_BUF.n5 D0_BUF.t0 47.274
R9 D0_BUF.n2 D0_BUF.t1 27.6955
R10 D0_BUF.n17 D0_BUF.n15 23.9595
R11 D0_BUF.n11 D0_BUF.n3 13.177
R12 D0_BUF.n8 D0_BUF.n3 13.177
R13 D0_BUF.n11 D0_BUF.n10 9.3005
R14 D0_BUF.n9 D0_BUF.n8 9.3005
R15 D0_BUF.n6 D0_BUF.n5 9.3005
R16 D0_BUF.n7 D0_BUF.n4 9.3005
R17 D0_BUF.n12 D0_BUF.n1 9.3005
R18 D0_BUF.n14 D0_BUF.n13 9.3005
R19 D0_BUF.n13 D0_BUF.n2 9.02061
R20 D0_BUF.n6 D0_BUF.n2 9.0206
R21 D0_BUF.n13 D0_BUF.n12 6.02403
R22 D0_BUF.n7 D0_BUF.n6 6.02403
R23 D0_BUF.n15 D0_BUF 5.08342
R24 D0_BUF D0_BUF.n14 2.37139
R25 D0_BUF.n12 D0_BUF.n11 0.376971
R26 D0_BUF.n8 D0_BUF.n7 0.376971
R27 D0_BUF.n10 D0_BUF.n9 0.190717
R28 D0_BUF.n14 D0_BUF.n1 0.0439783
R29 D0_BUF.n5 D0_BUF.n4 0.0439783
R30 D0_BUF.n10 D0_BUF.n1 0.00321739
R31 D0_BUF.n9 D0_BUF.n4 0.00321739
R32 VCC.n792 VCC.t6 4282.54
R33 VCC.n1344 VCC.t64 4282.54
R34 VCC.n1902 VCC.t13 4282.54
R35 VCC.t63 VCC.n227 4282.54
R36 VCC.t54 VCC.t3 1149.1
R37 VCC.t33 VCC.t65 1149.1
R38 VCC.t29 VCC.t12 1149.1
R39 VCC.t62 VCC.t24 1149.1
R40 VCC.t6 VCC.t54 978.443
R41 VCC.t64 VCC.t33 978.443
R42 VCC.t13 VCC.t29 978.443
R43 VCC.t24 VCC.t63 978.443
R44 VCC.t3 VCC.t51 972.755
R45 VCC.t65 VCC.t34 972.755
R46 VCC.t12 VCC.t26 972.755
R47 VCC.t25 VCC.t62 972.755
R48 VCC.t51 VCC.n791 723.087
R49 VCC.t34 VCC.n1343 723.087
R50 VCC.t26 VCC.n1901 723.087
R51 VCC.n230 VCC.t25 723.087
R52 VCC.t14 VCC.t2 571.485
R53 VCC.t17 VCC.t35 571.485
R54 VCC.t30 VCC.t7 571.485
R55 VCC.t71 VCC.t46 571.485
R56 VCC.t70 VCC.t56 571.485
R57 VCC.t55 VCC.t61 571.485
R58 VCC.t43 VCC.t42 571.485
R59 VCC.n488 VCC.t17 544.823
R60 VCC.n1040 VCC.t71 544.823
R61 VCC.n1597 VCC.t70 544.823
R62 VCC.n27 VCC.t43 544.823
R63 VCC.n575 VCC.t14 542.996
R64 VCC.n1127 VCC.t30 542.996
R65 VCC.n1685 VCC.t55 542.996
R66 VCC.n575 VCC.n560 187.349
R67 VCC.n489 VCC.n488 187.349
R68 VCC.n792 VCC.n445 187.349
R69 VCC.n1127 VCC.n1112 187.349
R70 VCC.n1041 VCC.n1040 187.349
R71 VCC.n1344 VCC.n997 187.349
R72 VCC.n1598 VCC.n1597 187.349
R73 VCC.n1902 VCC.n1554 187.349
R74 VCC.n1685 VCC.n1670 187.349
R75 VCC.n597 VCC.n596 185
R76 VCC.n596 VCC.n595 185
R77 VCC.n636 VCC.n635 185
R78 VCC.n635 VCC.n634 185
R79 VCC.n652 VCC.n506 185
R80 VCC.n656 VCC.n506 185
R81 VCC.n658 VCC.n507 185
R82 VCC.n658 VCC.n657 185
R83 VCC.n637 VCC.n509 185
R84 VCC.n509 VCC.n508 185
R85 VCC.n576 VCC.n574 185
R86 VCC.n549 VCC.n548 185
R87 VCC.n548 VCC.n547 185
R88 VCC.n591 VCC.n590 185
R89 VCC.n592 VCC.n591 185
R90 VCC.n546 VCC.n544 185
R91 VCC.n594 VCC.n546 185
R92 VCC.n725 VCC.n724 185
R93 VCC.n726 VCC.n725 185
R94 VCC.n458 VCC.n457 185
R95 VCC.n761 VCC.n458 185
R96 VCC.n782 VCC.n781 185
R97 VCC.n783 VCC.n782 185
R98 VCC.n780 VCC.n446 185
R99 VCC.n784 VCC.n446 185
R100 VCC.n764 VCC.n763 185
R101 VCC.n763 VCC.n762 185
R102 VCC.n793 VCC.n447 185
R103 VCC.n487 VCC.n486 185
R104 VCC.n485 VCC.n484 185
R105 VCC.n702 VCC.n485 185
R106 VCC.n705 VCC.n704 185
R107 VCC.n704 VCC.n703 185
R108 VCC.n473 VCC.n472 185
R109 VCC.n727 VCC.n473 185
R110 VCC.n912 VCC.n911 185
R111 VCC.n913 VCC.n912 185
R112 VCC.n787 VCC.n422 185
R113 VCC.n785 VCC.n422 185
R114 VCC.n859 VCC.n405 185
R115 VCC.n860 VCC.n859 185
R116 VCC.n387 VCC.n386 185
R117 VCC.n892 VCC.n387 185
R118 VCC.n895 VCC.n894 185
R119 VCC.n894 VCC.n893 185
R120 VCC.n390 VCC.n389 185
R121 VCC.n389 VCC.n388 185
R122 VCC.n864 VCC.n863 185
R123 VCC.n863 VCC.n862 185
R124 VCC.n858 VCC.n857 185
R125 VCC.n858 VCC.n407 185
R126 VCC.n841 VCC.n840 185
R127 VCC.n840 VCC.n839 185
R128 VCC.n421 VCC.n420 185
R129 VCC.n837 VCC.n421 185
R130 VCC.n789 VCC.n788 185
R131 VCC.n789 VCC.n786 185
R132 VCC.n370 VCC.n369 185
R133 VCC.n1149 VCC.n1148 185
R134 VCC.n1148 VCC.n1147 185
R135 VCC.n1188 VCC.n1187 185
R136 VCC.n1187 VCC.n1186 185
R137 VCC.n1204 VCC.n1058 185
R138 VCC.n1208 VCC.n1058 185
R139 VCC.n1210 VCC.n1059 185
R140 VCC.n1210 VCC.n1209 185
R141 VCC.n1189 VCC.n1061 185
R142 VCC.n1061 VCC.n1060 185
R143 VCC.n1128 VCC.n1126 185
R144 VCC.n1101 VCC.n1100 185
R145 VCC.n1100 VCC.n1099 185
R146 VCC.n1143 VCC.n1142 185
R147 VCC.n1144 VCC.n1143 185
R148 VCC.n1098 VCC.n1096 185
R149 VCC.n1146 VCC.n1098 185
R150 VCC.n1277 VCC.n1276 185
R151 VCC.n1278 VCC.n1277 185
R152 VCC.n1010 VCC.n1009 185
R153 VCC.n1313 VCC.n1010 185
R154 VCC.n1334 VCC.n1333 185
R155 VCC.n1335 VCC.n1334 185
R156 VCC.n1332 VCC.n998 185
R157 VCC.n1336 VCC.n998 185
R158 VCC.n1316 VCC.n1315 185
R159 VCC.n1315 VCC.n1314 185
R160 VCC.n1345 VCC.n999 185
R161 VCC.n1039 VCC.n1038 185
R162 VCC.n1037 VCC.n1036 185
R163 VCC.n1254 VCC.n1037 185
R164 VCC.n1257 VCC.n1256 185
R165 VCC.n1256 VCC.n1255 185
R166 VCC.n1025 VCC.n1024 185
R167 VCC.n1279 VCC.n1025 185
R168 VCC.n1339 VCC.n974 185
R169 VCC.n1337 VCC.n974 185
R170 VCC.n973 VCC.n972 185
R171 VCC.n1389 VCC.n973 185
R172 VCC.n1410 VCC.n1409 185
R173 VCC.n1410 VCC.n959 185
R174 VCC.n942 VCC.n941 185
R175 VCC.n941 VCC.n940 185
R176 VCC.n1447 VCC.n1446 185
R177 VCC.n1446 VCC.n1445 185
R178 VCC.n1466 VCC.n1465 185
R179 VCC.n1467 VCC.n1466 185
R180 VCC.n1416 VCC.n1415 185
R181 VCC.n1415 VCC.n1414 185
R182 VCC.n1393 VCC.n1392 185
R183 VCC.n1392 VCC.n1391 185
R184 VCC.n1411 VCC.n957 185
R185 VCC.n1412 VCC.n1411 185
R186 VCC.n939 VCC.n938 185
R187 VCC.n1444 VCC.n939 185
R188 VCC.n924 VCC.n923 185
R189 VCC.n1341 VCC.n1340 185
R190 VCC.n1341 VCC.n1338 185
R191 VCC.n1897 VCC.n1896 185
R192 VCC.n1896 VCC.n1895 185
R193 VCC.n1945 VCC.n1944 185
R194 VCC.n1946 VCC.n1945 185
R195 VCC.n1528 VCC.n1526 185
R196 VCC.n1950 VCC.n1528 185
R197 VCC.n1508 VCC.n1501 185
R198 VCC.n1986 VCC.n1508 185
R199 VCC.n2016 VCC.n2015 185
R200 VCC.n2017 VCC.n2016 185
R201 VCC.n2020 VCC.n1478 185
R202 VCC.n2020 VCC.n2019 185
R203 VCC.n1482 VCC.n1481 185
R204 VCC.n1481 VCC.n1480 185
R205 VCC.n1984 VCC.n1983 185
R206 VCC.n1985 VCC.n1984 185
R207 VCC.n1948 VCC.n1511 185
R208 VCC.n1949 VCC.n1948 185
R209 VCC.n1527 VCC.n1525 185
R210 VCC.n1947 VCC.n1527 185
R211 VCC.n2022 VCC.n2021 185
R212 VCC.n1899 VCC.n1898 185
R213 VCC.n1899 VCC.n1894 185
R214 VCC.n1814 VCC.n1813 185
R215 VCC.n1813 VCC.n1812 185
R216 VCC.n1582 VCC.n1581 185
R217 VCC.n1836 VCC.n1582 185
R218 VCC.n1567 VCC.n1566 185
R219 VCC.n1870 VCC.n1567 185
R220 VCC.n1891 VCC.n1890 185
R221 VCC.n1892 VCC.n1891 185
R222 VCC.n1889 VCC.n1555 185
R223 VCC.n1893 VCC.n1555 185
R224 VCC.n1834 VCC.n1833 185
R225 VCC.n1835 VCC.n1834 185
R226 VCC.n1594 VCC.n1593 185
R227 VCC.n1811 VCC.n1594 185
R228 VCC.n1873 VCC.n1872 185
R229 VCC.n1872 VCC.n1871 185
R230 VCC.n1903 VCC.n1556 185
R231 VCC.n1596 VCC.n1595 185
R232 VCC.n1701 VCC.n1700 185
R233 VCC.n1702 VCC.n1701 185
R234 VCC.n1656 VCC.n1654 185
R235 VCC.n1704 VCC.n1656 185
R236 VCC.n1746 VCC.n1745 185
R237 VCC.n1745 VCC.n1744 185
R238 VCC.n1762 VCC.n1616 185
R239 VCC.n1766 VCC.n1616 185
R240 VCC.n1768 VCC.n1617 185
R241 VCC.n1768 VCC.n1767 185
R242 VCC.n1707 VCC.n1706 185
R243 VCC.n1706 VCC.n1705 185
R244 VCC.n1659 VCC.n1658 185
R245 VCC.n1658 VCC.n1657 185
R246 VCC.n1747 VCC.n1619 185
R247 VCC.n1619 VCC.n1618 185
R248 VCC.n1686 VCC.n1684 185
R249 VCC.n595 VCC.n593 96.8274
R250 VCC.n655 VCC.n508 96.8274
R251 VCC.n726 VCC.n474 96.8274
R252 VCC.n762 VCC.n448 96.8274
R253 VCC.n1147 VCC.n1145 96.8274
R254 VCC.n1207 VCC.n1060 96.8274
R255 VCC.n1278 VCC.n1026 96.8274
R256 VCC.n1314 VCC.n1000 96.8274
R257 VCC.n1835 VCC.n1583 96.8274
R258 VCC.n1871 VCC.n1557 96.8274
R259 VCC.n1705 VCC.n1703 96.8274
R260 VCC.n1765 VCC.n1618 96.8274
R261 VCC.n632 VCC.n519 95.0005
R262 VCC.n633 VCC.n632 95.0005
R263 VCC.n728 VCC.n459 95.0005
R264 VCC.n760 VCC.n459 95.0005
R265 VCC.n1184 VCC.n1071 95.0005
R266 VCC.n1185 VCC.n1184 95.0005
R267 VCC.n1280 VCC.n1011 95.0005
R268 VCC.n1312 VCC.n1011 95.0005
R269 VCC.n1837 VCC.n1568 95.0005
R270 VCC.n1869 VCC.n1568 95.0005
R271 VCC.n1742 VCC.n1629 95.0005
R272 VCC.n1743 VCC.n1742 95.0005
R273 VCC.n197 VCC.n194 95.0005
R274 VCC.n839 VCC.n838 93.2412
R275 VCC.n861 VCC.n860 93.2412
R276 VCC.n862 VCC.n861 93.2412
R277 VCC.n913 VCC.n371 93.2412
R278 VCC.n1391 VCC.n1390 93.2412
R279 VCC.n1413 VCC.n1412 93.2412
R280 VCC.n1414 VCC.n1413 93.2412
R281 VCC.n1467 VCC.n925 93.2412
R282 VCC.n1951 VCC.n1947 93.2412
R283 VCC.n1949 VCC.n1509 93.2412
R284 VCC.n1985 VCC.n1509 93.2412
R285 VCC.n2019 VCC.n2018 93.2412
R286 VCC.n579 VCC.n560 92.5398
R287 VCC.n699 VCC.n489 92.5398
R288 VCC.n796 VCC.n445 92.5398
R289 VCC.n1131 VCC.n1112 92.5398
R290 VCC.n1251 VCC.n1041 92.5398
R291 VCC.n1348 VCC.n997 92.5398
R292 VCC.n1808 VCC.n1598 92.5398
R293 VCC.n1906 VCC.n1554 92.5398
R294 VCC.n1689 VCC.n1670 92.5398
R295 VCC.n631 VCC.n630 92.5005
R296 VCC.n632 VCC.n631 92.5005
R297 VCC.n751 VCC.n460 92.5005
R298 VCC.n460 VCC.n459 92.5005
R299 VCC.n1183 VCC.n1182 92.5005
R300 VCC.n1184 VCC.n1183 92.5005
R301 VCC.n1303 VCC.n1012 92.5005
R302 VCC.n1012 VCC.n1011 92.5005
R303 VCC.n1860 VCC.n1569 92.5005
R304 VCC.n1569 VCC.n1568 92.5005
R305 VCC.n1741 VCC.n1740 92.5005
R306 VCC.n1742 VCC.n1741 92.5005
R307 VCC.n577 VCC.t0 74.9043
R308 VCC.n1129 VCC.t8 74.9043
R309 VCC.n1687 VCC.t59 74.9043
R310 VCC.t36 VCC.n701 73.0774
R311 VCC.t44 VCC.n1253 73.0774
R312 VCC.t57 VCC.n1810 73.0774
R313 VCC.n659 VCC.t38 72.544
R314 VCC.n1211 VCC.t49 72.544
R315 VCC.n1769 VCC.t15 72.544
R316 VCC.t20 VCC.n891 70.3709
R317 VCC.t4 VCC.n1443 70.3709
R318 VCC.n1987 VCC.t66 70.3709
R319 VCC.n836 VCC.t52 66.8524
R320 VCC.n1388 VCC.t31 66.8524
R321 VCC.t27 VCC.n1529 66.8524
R322 VCC.n794 VCC.t47 65.7697
R323 VCC.n1346 VCC.t18 65.7697
R324 VCC.n1904 VCC.t72 65.7697
R325 VCC.n225 VCC.t68 65.7697
R326 VCC.n659 VCC.n658 50.4194
R327 VCC.n1211 VCC.n1210 50.4194
R328 VCC.n1769 VCC.n1768 50.4194
R329 VCC.n578 VCC.n548 50.3505
R330 VCC.n596 VCC.n545 50.3505
R331 VCC.n654 VCC.n509 50.3505
R332 VCC.n700 VCC.n485 50.3505
R333 VCC.n725 VCC.n475 50.3505
R334 VCC.n763 VCC.n449 50.3505
R335 VCC.n795 VCC.n446 50.3505
R336 VCC.n1130 VCC.n1100 50.3505
R337 VCC.n1148 VCC.n1097 50.3505
R338 VCC.n1206 VCC.n1061 50.3505
R339 VCC.n1252 VCC.n1037 50.3505
R340 VCC.n1277 VCC.n1027 50.3505
R341 VCC.n1315 VCC.n1001 50.3505
R342 VCC.n1347 VCC.n998 50.3505
R343 VCC.n1809 VCC.n1594 50.3505
R344 VCC.n1834 VCC.n1584 50.3505
R345 VCC.n1872 VCC.n1558 50.3505
R346 VCC.n1905 VCC.n1555 50.3505
R347 VCC.n1688 VCC.n1658 50.3505
R348 VCC.n1706 VCC.n1655 50.3505
R349 VCC.n1764 VCC.n1619 50.3505
R350 VCC.n631 VCC.n520 49.4005
R351 VCC.n631 VCC.n518 49.4005
R352 VCC.n729 VCC.n460 49.4005
R353 VCC.n759 VCC.n460 49.4005
R354 VCC.n1183 VCC.n1072 49.4005
R355 VCC.n1183 VCC.n1070 49.4005
R356 VCC.n1281 VCC.n1012 49.4005
R357 VCC.n1311 VCC.n1012 49.4005
R358 VCC.n1838 VCC.n1569 49.4005
R359 VCC.n1868 VCC.n1569 49.4005
R360 VCC.n1741 VCC.n1630 49.4005
R361 VCC.n1741 VCC.n1628 49.4005
R362 VCC.n198 VCC.n191 49.4005
R363 VCC.n835 VCC.n422 43.1576
R364 VCC.n840 VCC.n408 43.1576
R365 VCC.n859 VCC.n406 43.1576
R366 VCC.n863 VCC.n406 43.1576
R367 VCC.n890 VCC.n387 43.1576
R368 VCC.n912 VCC.n372 43.1576
R369 VCC.n1387 VCC.n974 43.1576
R370 VCC.n1392 VCC.n960 43.1576
R371 VCC.n1411 VCC.n958 43.1576
R372 VCC.n1415 VCC.n958 43.1576
R373 VCC.n1442 VCC.n939 43.1576
R374 VCC.n1466 VCC.n926 43.1576
R375 VCC.n1896 VCC.n1530 43.1576
R376 VCC.n1952 VCC.n1527 43.1576
R377 VCC.n1948 VCC.n1510 43.1576
R378 VCC.n1984 VCC.n1510 43.1576
R379 VCC.n1988 VCC.n1481 43.1576
R380 VCC.n2020 VCC.n1479 43.1576
R381 VCC.n914 VCC.n913 36.8662
R382 VCC.n1468 VCC.n1467 36.8662
R383 VCC.n2019 VCC.n1477 36.8662
R384 VCC.n284 VCC.n283 36.8662
R385 VCC.n812 VCC.t48 35.5869
R386 VCC.n1364 VCC.t19 35.5869
R387 VCC.n1922 VCC.t73 35.5869
R388 VCC.n218 VCC.t69 35.5869
R389 VCC.n377 VCC.t21 34.994
R390 VCC.n1457 VCC.t5 34.994
R391 VCC.n2006 VCC.t67 34.994
R392 VCC.n289 VCC.t11 34.994
R393 VCC.n418 VCC.t53 34.9892
R394 VCC.n970 VCC.t32 34.9892
R395 VCC.n1523 VCC.t28 34.9892
R396 VCC.n254 VCC.t23 34.9892
R397 VCC.n677 VCC.t39 34.9619
R398 VCC.n1229 VCC.t50 34.9619
R399 VCC.n1787 VCC.t16 34.9619
R400 VCC.n478 VCC.t37 34.945
R401 VCC.n1030 VCC.t45 34.945
R402 VCC.n1587 VCC.t58 34.945
R403 VCC.n60 VCC.t41 34.945
R404 VCC.n603 VCC.t1 34.9423
R405 VCC.n1155 VCC.t9 34.9423
R406 VCC.n1713 VCC.t60 34.9423
R407 VCC.n657 VCC.t38 32.8851
R408 VCC.n1209 VCC.t49 32.8851
R409 VCC.n1767 VCC.t15 32.8851
R410 VCC.t47 VCC.n784 31.0582
R411 VCC.t18 VCC.n1336 31.0582
R412 VCC.t72 VCC.n1893 31.0582
R413 VCC.n594 VCC.n519 29.2313
R414 VCC.n634 VCC.n633 29.2313
R415 VCC.n728 VCC.n727 29.2313
R416 VCC.n761 VCC.n760 29.2313
R417 VCC.n1146 VCC.n1071 29.2313
R418 VCC.n1186 VCC.n1185 29.2313
R419 VCC.n1280 VCC.n1279 29.2313
R420 VCC.n1313 VCC.n1312 29.2313
R421 VCC.n1837 VCC.n1836 29.2313
R422 VCC.n1870 VCC.n1869 29.2313
R423 VCC.n1704 VCC.n1629 29.2313
R424 VCC.n1744 VCC.n1743 29.2313
R425 VCC.n71 VCC.n70 29.2313
R426 VCC.n197 VCC.n196 29.2313
R427 VCC.n785 VCC.t52 26.3894
R428 VCC.n860 VCC.n407 26.3894
R429 VCC.n862 VCC.n388 26.3894
R430 VCC.n1337 VCC.t31 26.3894
R431 VCC.n1412 VCC.n959 26.3894
R432 VCC.n1414 VCC.n940 26.3894
R433 VCC.n1895 VCC.t27 26.3894
R434 VCC.n1950 VCC.n1949 26.3894
R435 VCC.n1986 VCC.n1985 26.3894
R436 VCC.n228 VCC.t22 26.3894
R437 VCC.n264 VCC.n263 26.3894
R438 VCC.n320 VCC.n319 26.3894
R439 VCC.n593 VCC.n592 25.5774
R440 VCC.n656 VCC.n655 25.5774
R441 VCC.n703 VCC.n474 25.5774
R442 VCC.n783 VCC.n448 25.5774
R443 VCC.n1145 VCC.n1144 25.5774
R444 VCC.n1208 VCC.n1207 25.5774
R445 VCC.n1255 VCC.n1026 25.5774
R446 VCC.n1335 VCC.n1000 25.5774
R447 VCC.n1812 VCC.n1583 25.5774
R448 VCC.n1892 VCC.n1557 25.5774
R449 VCC.n1703 VCC.n1702 25.5774
R450 VCC.n1766 VCC.n1765 25.5774
R451 VCC.n50 VCC.n49 25.5774
R452 VCC.n16 VCC.n15 25.5774
R453 VCC.n702 VCC.t36 23.7505
R454 VCC.n1254 VCC.t44 23.7505
R455 VCC.n1811 VCC.t57 23.7505
R456 VCC.n48 VCC.t40 23.7505
R457 VCC.n839 VCC.n837 22.8709
R458 VCC.n892 VCC.t20 22.8709
R459 VCC.n893 VCC.n892 22.8709
R460 VCC.n1391 VCC.n1389 22.8709
R461 VCC.n1444 VCC.t4 22.8709
R462 VCC.n1445 VCC.n1444 22.8709
R463 VCC.n1947 VCC.n1946 22.8709
R464 VCC.t66 VCC.n1480 22.8709
R465 VCC.n2017 VCC.n1480 22.8709
R466 VCC.n244 VCC.n243 22.8709
R467 VCC.n299 VCC.t10 22.8709
R468 VCC.n300 VCC.n299 22.8709
R469 VCC.n577 VCC.n576 21.9236
R470 VCC.t0 VCC.n547 21.9236
R471 VCC.n701 VCC.n486 21.9236
R472 VCC.n794 VCC.n793 21.9236
R473 VCC.n1129 VCC.n1128 21.9236
R474 VCC.t8 VCC.n1099 21.9236
R475 VCC.n1253 VCC.n1038 21.9236
R476 VCC.n1346 VCC.n1345 21.9236
R477 VCC.n1810 VCC.n1595 21.9236
R478 VCC.n1904 VCC.n1903 21.9236
R479 VCC.n1687 VCC.n1686 21.9236
R480 VCC.t59 VCC.n1657 21.9236
R481 VCC.n29 VCC.n28 21.9236
R482 VCC.n226 VCC.n225 21.9236
R483 VCC.n786 VCC.n785 19.3524
R484 VCC.n1338 VCC.n1337 19.3524
R485 VCC.n1895 VCC.n1894 19.3524
R486 VCC.n229 VCC.n228 19.3524
R487 VCC.n546 VCC.n520 15.2005
R488 VCC.n635 VCC.n518 15.2005
R489 VCC.n729 VCC.n473 15.2005
R490 VCC.n759 VCC.n458 15.2005
R491 VCC.n1098 VCC.n1072 15.2005
R492 VCC.n1187 VCC.n1070 15.2005
R493 VCC.n1281 VCC.n1025 15.2005
R494 VCC.n1311 VCC.n1010 15.2005
R495 VCC.n1838 VCC.n1582 15.2005
R496 VCC.n1868 VCC.n1567 15.2005
R497 VCC.n1656 VCC.n1630 15.2005
R498 VCC.n1745 VCC.n1628 15.2005
R499 VCC.n72 VCC.n68 15.2005
R500 VCC.n198 VCC.n193 15.2005
R501 VCC.n591 VCC.n545 13.3005
R502 VCC.n654 VCC.n506 13.3005
R503 VCC.n704 VCC.n475 13.3005
R504 VCC.n782 VCC.n449 13.3005
R505 VCC.n1143 VCC.n1097 13.3005
R506 VCC.n1206 VCC.n1058 13.3005
R507 VCC.n1256 VCC.n1027 13.3005
R508 VCC.n1334 VCC.n1001 13.3005
R509 VCC.n1813 VCC.n1584 13.3005
R510 VCC.n1891 VCC.n1558 13.3005
R511 VCC.n1701 VCC.n1655 13.3005
R512 VCC.n1764 VCC.n1616 13.3005
R513 VCC.n51 VCC.n47 13.3005
R514 VCC.n17 VCC.n13 13.3005
R515 VCC.n859 VCC.n858 12.2148
R516 VCC.n863 VCC.n389 12.2148
R517 VCC.n1411 VCC.n1410 12.2148
R518 VCC.n1415 VCC.n941 12.2148
R519 VCC.n1948 VCC.n1528 12.2148
R520 VCC.n1984 VCC.n1508 12.2148
R521 VCC.n262 VCC.n261 12.2148
R522 VCC.n318 VCC.n317 12.2148
R523 VCC.n578 VCC.n574 11.4005
R524 VCC.n700 VCC.n487 11.4005
R525 VCC.n795 VCC.n447 11.4005
R526 VCC.n1130 VCC.n1126 11.4005
R527 VCC.n1252 VCC.n1039 11.4005
R528 VCC.n1347 VCC.n999 11.4005
R529 VCC.n1809 VCC.n1596 11.4005
R530 VCC.n1905 VCC.n1556 11.4005
R531 VCC.n1688 VCC.n1684 11.4005
R532 VCC.n30 VCC.n26 11.4005
R533 VCC.n224 VCC.n6 11.4005
R534 VCC.n840 VCC.n421 10.5862
R535 VCC.n894 VCC.n387 10.5862
R536 VCC.n1392 VCC.n973 10.5862
R537 VCC.n1446 VCC.n939 10.5862
R538 VCC.n1945 VCC.n1527 10.5862
R539 VCC.n2016 VCC.n1481 10.5862
R540 VCC.n242 VCC.n241 10.5862
R541 VCC.n298 VCC.n297 10.5862
R542 VCC.n791 VCC.n786 10.5561
R543 VCC.n1343 VCC.n1338 10.5561
R544 VCC.n1901 VCC.n1894 10.5561
R545 VCC.n230 VCC.n229 10.5561
R546 VCC.n915 VCC.n914 9.80483
R547 VCC.n1469 VCC.n1468 9.80483
R548 VCC.n2023 VCC.n1477 9.80483
R549 VCC.n285 VCC.n284 9.80483
R550 VCC.n790 VCC.n431 9.38146
R551 VCC.n1342 VCC.n983 9.38146
R552 VCC.n232 VCC.n231 9.38146
R553 VCC.n1900 VCC.n1540 9.38145
R554 VCC.n599 VCC.n598 9.3005
R555 VCC.n568 VCC.n567 9.3005
R556 VCC.n664 VCC.n663 9.3005
R557 VCC.n639 VCC.n638 9.3005
R558 VCC.n527 VCC.n526 9.3005
R559 VCC.n528 VCC.n522 9.3005
R560 VCC.n517 VCC.n516 9.3005
R561 VCC.n518 VCC.n517 9.3005
R562 VCC.n633 VCC.n518 9.3005
R563 VCC.n511 VCC.n510 9.3005
R564 VCC.n653 VCC.n500 9.3005
R565 VCC.n654 VCC.n653 9.3005
R566 VCC.n655 VCC.n654 9.3005
R567 VCC.n505 VCC.n503 9.3005
R568 VCC.n661 VCC.n660 9.3005
R569 VCC.n543 VCC.n542 9.3005
R570 VCC.n580 VCC.n579 9.3005
R571 VCC.n579 VCC.n578 9.3005
R572 VCC.n578 VCC.n577 9.3005
R573 VCC.n562 VCC.n561 9.3005
R574 VCC.n589 VCC.n588 9.3005
R575 VCC.n589 VCC.n545 9.3005
R576 VCC.n593 VCC.n545 9.3005
R577 VCC.n536 VCC.n535 9.3005
R578 VCC.n535 VCC.n520 9.3005
R579 VCC.n520 VCC.n519 9.3005
R580 VCC.n614 VCC.n534 9.3005
R581 VCC.n616 VCC.n615 9.3005
R582 VCC.n723 VCC.n722 9.3005
R583 VCC.n693 VCC.n692 9.3005
R584 VCC.n799 VCC.n798 9.3005
R585 VCC.n766 VCC.n765 9.3005
R586 VCC.n755 VCC.n461 9.3005
R587 VCC.n754 VCC.n753 9.3005
R588 VCC.n451 VCC.n450 9.3005
R589 VCC.n444 VCC.n442 9.3005
R590 VCC.n477 VCC.n476 9.3005
R591 VCC.n691 VCC.n686 9.3005
R592 VCC.n731 VCC.n471 9.3005
R593 VCC.n464 VCC.n463 9.3005
R594 VCC.n758 VCC.n456 9.3005
R595 VCC.n759 VCC.n758 9.3005
R596 VCC.n760 VCC.n759 9.3005
R597 VCC.n779 VCC.n439 9.3005
R598 VCC.n779 VCC.n449 9.3005
R599 VCC.n449 VCC.n448 9.3005
R600 VCC.n796 VCC.n434 9.3005
R601 VCC.n796 VCC.n795 9.3005
R602 VCC.n795 VCC.n794 9.3005
R603 VCC.n699 VCC.n698 9.3005
R604 VCC.n700 VCC.n699 9.3005
R605 VCC.n701 VCC.n700 9.3005
R606 VCC.n708 VCC.n707 9.3005
R607 VCC.n707 VCC.n475 9.3005
R608 VCC.n475 VCC.n474 9.3005
R609 VCC.n730 VCC.n470 9.3005
R610 VCC.n730 VCC.n729 9.3005
R611 VCC.n729 VCC.n728 9.3005
R612 VCC.n843 VCC.n842 9.3005
R613 VCC.n889 VCC.n888 9.3005
R614 VCC.n890 VCC.n889 9.3005
R615 VCC.n891 VCC.n890 9.3005
R616 VCC.n374 VCC.n373 9.3005
R617 VCC.n882 VCC.n881 9.3005
R618 VCC.n910 VCC.n909 9.3005
R619 VCC.n898 VCC.n897 9.3005
R620 VCC.n897 VCC.n372 9.3005
R621 VCC.n372 VCC.n371 9.3005
R622 VCC.n856 VCC.n855 9.3005
R623 VCC.n856 VCC.n408 9.3005
R624 VCC.n838 VCC.n408 9.3005
R625 VCC.n835 VCC.n834 9.3005
R626 VCC.n836 VCC.n835 9.3005
R627 VCC.n791 VCC.n790 9.3005
R628 VCC.n1151 VCC.n1150 9.3005
R629 VCC.n1120 VCC.n1119 9.3005
R630 VCC.n1216 VCC.n1215 9.3005
R631 VCC.n1191 VCC.n1190 9.3005
R632 VCC.n1079 VCC.n1078 9.3005
R633 VCC.n1080 VCC.n1074 9.3005
R634 VCC.n1069 VCC.n1068 9.3005
R635 VCC.n1070 VCC.n1069 9.3005
R636 VCC.n1185 VCC.n1070 9.3005
R637 VCC.n1063 VCC.n1062 9.3005
R638 VCC.n1205 VCC.n1052 9.3005
R639 VCC.n1206 VCC.n1205 9.3005
R640 VCC.n1207 VCC.n1206 9.3005
R641 VCC.n1057 VCC.n1055 9.3005
R642 VCC.n1213 VCC.n1212 9.3005
R643 VCC.n1095 VCC.n1094 9.3005
R644 VCC.n1132 VCC.n1131 9.3005
R645 VCC.n1131 VCC.n1130 9.3005
R646 VCC.n1130 VCC.n1129 9.3005
R647 VCC.n1114 VCC.n1113 9.3005
R648 VCC.n1141 VCC.n1140 9.3005
R649 VCC.n1141 VCC.n1097 9.3005
R650 VCC.n1145 VCC.n1097 9.3005
R651 VCC.n1088 VCC.n1087 9.3005
R652 VCC.n1087 VCC.n1072 9.3005
R653 VCC.n1072 VCC.n1071 9.3005
R654 VCC.n1166 VCC.n1086 9.3005
R655 VCC.n1168 VCC.n1167 9.3005
R656 VCC.n1275 VCC.n1274 9.3005
R657 VCC.n1245 VCC.n1244 9.3005
R658 VCC.n1351 VCC.n1350 9.3005
R659 VCC.n1318 VCC.n1317 9.3005
R660 VCC.n1307 VCC.n1013 9.3005
R661 VCC.n1306 VCC.n1305 9.3005
R662 VCC.n1003 VCC.n1002 9.3005
R663 VCC.n996 VCC.n994 9.3005
R664 VCC.n1029 VCC.n1028 9.3005
R665 VCC.n1243 VCC.n1238 9.3005
R666 VCC.n1283 VCC.n1023 9.3005
R667 VCC.n1016 VCC.n1015 9.3005
R668 VCC.n1310 VCC.n1008 9.3005
R669 VCC.n1311 VCC.n1310 9.3005
R670 VCC.n1312 VCC.n1311 9.3005
R671 VCC.n1331 VCC.n991 9.3005
R672 VCC.n1331 VCC.n1001 9.3005
R673 VCC.n1001 VCC.n1000 9.3005
R674 VCC.n1348 VCC.n986 9.3005
R675 VCC.n1348 VCC.n1347 9.3005
R676 VCC.n1347 VCC.n1346 9.3005
R677 VCC.n1251 VCC.n1250 9.3005
R678 VCC.n1252 VCC.n1251 9.3005
R679 VCC.n1253 VCC.n1252 9.3005
R680 VCC.n1260 VCC.n1259 9.3005
R681 VCC.n1259 VCC.n1027 9.3005
R682 VCC.n1027 VCC.n1026 9.3005
R683 VCC.n1282 VCC.n1022 9.3005
R684 VCC.n1282 VCC.n1281 9.3005
R685 VCC.n1281 VCC.n1280 9.3005
R686 VCC.n1441 VCC.n1440 9.3005
R687 VCC.n1442 VCC.n1441 9.3005
R688 VCC.n1443 VCC.n1442 9.3005
R689 VCC.n1387 VCC.n1386 9.3005
R690 VCC.n1388 VCC.n1387 9.3005
R691 VCC.n1395 VCC.n1394 9.3005
R692 VCC.n1408 VCC.n1407 9.3005
R693 VCC.n1408 VCC.n960 9.3005
R694 VCC.n1390 VCC.n960 9.3005
R695 VCC.n1434 VCC.n1433 9.3005
R696 VCC.n1450 VCC.n1449 9.3005
R697 VCC.n1449 VCC.n926 9.3005
R698 VCC.n926 VCC.n925 9.3005
R699 VCC.n928 VCC.n927 9.3005
R700 VCC.n1464 VCC.n1463 9.3005
R701 VCC.n1343 VCC.n1342 9.3005
R702 VCC.n1506 VCC.n1505 9.3005
R703 VCC.n1491 VCC.n1490 9.3005
R704 VCC.n1489 VCC.n1488 9.3005
R705 VCC.n1961 VCC.n1960 9.3005
R706 VCC.n1954 VCC.n1953 9.3005
R707 VCC.n1953 VCC.n1952 9.3005
R708 VCC.n1952 VCC.n1951 9.3005
R709 VCC.n2014 VCC.n2013 9.3005
R710 VCC.n2014 VCC.n1479 9.3005
R711 VCC.n2018 VCC.n1479 9.3005
R712 VCC.n1990 VCC.n1989 9.3005
R713 VCC.n1989 VCC.n1988 9.3005
R714 VCC.n1988 VCC.n1987 9.3005
R715 VCC.n1943 VCC.n1530 9.3005
R716 VCC.n1530 VCC.n1529 9.3005
R717 VCC.n1901 VCC.n1900 9.3005
R718 VCC.n1909 VCC.n1908 9.3005
R719 VCC.n1875 VCC.n1874 9.3005
R720 VCC.n1864 VCC.n1570 9.3005
R721 VCC.n1573 VCC.n1572 9.3005
R722 VCC.n1817 VCC.n1816 9.3005
R723 VCC.n1816 VCC.n1584 9.3005
R724 VCC.n1584 VCC.n1583 9.3005
R725 VCC.n1586 VCC.n1585 9.3005
R726 VCC.n1832 VCC.n1831 9.3005
R727 VCC.n1839 VCC.n1579 9.3005
R728 VCC.n1839 VCC.n1838 9.3005
R729 VCC.n1838 VCC.n1837 9.3005
R730 VCC.n1840 VCC.n1580 9.3005
R731 VCC.n1863 VCC.n1862 9.3005
R732 VCC.n1867 VCC.n1565 9.3005
R733 VCC.n1868 VCC.n1867 9.3005
R734 VCC.n1869 VCC.n1868 9.3005
R735 VCC.n1560 VCC.n1559 9.3005
R736 VCC.n1888 VCC.n1548 9.3005
R737 VCC.n1888 VCC.n1558 9.3005
R738 VCC.n1558 VCC.n1557 9.3005
R739 VCC.n1553 VCC.n1551 9.3005
R740 VCC.n1906 VCC.n1543 9.3005
R741 VCC.n1906 VCC.n1905 9.3005
R742 VCC.n1905 VCC.n1904 9.3005
R743 VCC.n1808 VCC.n1807 9.3005
R744 VCC.n1809 VCC.n1808 9.3005
R745 VCC.n1810 VCC.n1809 9.3005
R746 VCC.n1800 VCC.n1796 9.3005
R747 VCC.n1802 VCC.n1801 9.3005
R748 VCC.n1774 VCC.n1773 9.3005
R749 VCC.n1749 VCC.n1748 9.3005
R750 VCC.n1637 VCC.n1636 9.3005
R751 VCC.n1726 VCC.n1725 9.3005
R752 VCC.n1699 VCC.n1698 9.3005
R753 VCC.n1699 VCC.n1655 9.3005
R754 VCC.n1703 VCC.n1655 9.3005
R755 VCC.n1653 VCC.n1652 9.3005
R756 VCC.n1709 VCC.n1708 9.3005
R757 VCC.n1646 VCC.n1645 9.3005
R758 VCC.n1645 VCC.n1630 9.3005
R759 VCC.n1630 VCC.n1629 9.3005
R760 VCC.n1724 VCC.n1644 9.3005
R761 VCC.n1638 VCC.n1632 9.3005
R762 VCC.n1627 VCC.n1626 9.3005
R763 VCC.n1628 VCC.n1627 9.3005
R764 VCC.n1743 VCC.n1628 9.3005
R765 VCC.n1621 VCC.n1620 9.3005
R766 VCC.n1763 VCC.n1610 9.3005
R767 VCC.n1764 VCC.n1763 9.3005
R768 VCC.n1765 VCC.n1764 9.3005
R769 VCC.n1615 VCC.n1613 9.3005
R770 VCC.n1771 VCC.n1770 9.3005
R771 VCC.n1690 VCC.n1689 9.3005
R772 VCC.n1689 VCC.n1688 9.3005
R773 VCC.n1688 VCC.n1687 9.3005
R774 VCC.n1672 VCC.n1671 9.3005
R775 VCC.n1678 VCC.n1677 9.3005
R776 VCC.n199 VCC.n198 9.3005
R777 VCC.n198 VCC.n197 9.3005
R778 VCC.n18 VCC.n17 9.3005
R779 VCC.n17 VCC.n16 9.3005
R780 VCC.n224 VCC.n223 9.3005
R781 VCC.n225 VCC.n224 9.3005
R782 VCC.n31 VCC.n30 9.3005
R783 VCC.n30 VCC.n29 9.3005
R784 VCC.n52 VCC.n51 9.3005
R785 VCC.n51 VCC.n50 9.3005
R786 VCC.n73 VCC.n72 9.3005
R787 VCC.n72 VCC.n71 9.3005
R788 VCC.n323 VCC.n322 9.3005
R789 VCC.n322 VCC.n321 9.3005
R790 VCC.n249 VCC.n246 9.3005
R791 VCC.n246 VCC.n245 9.3005
R792 VCC.n267 VCC.n266 9.3005
R793 VCC.n266 VCC.n265 9.3005
R794 VCC.n303 VCC.n302 9.3005
R795 VCC.n302 VCC.n301 9.3005
R796 VCC.n231 VCC.n230 9.3005
R797 VCC.n576 VCC.n575 9.13511
R798 VCC.n488 VCC.n486 9.13511
R799 VCC.n793 VCC.n792 9.13511
R800 VCC.n1128 VCC.n1127 9.13511
R801 VCC.n1040 VCC.n1038 9.13511
R802 VCC.n1345 VCC.n1344 9.13511
R803 VCC.n1597 VCC.n1595 9.13511
R804 VCC.n1903 VCC.n1902 9.13511
R805 VCC.n1686 VCC.n1685 9.13511
R806 VCC.n28 VCC.n27 9.13511
R807 VCC.n227 VCC.n226 9.13511
R808 VCC.n789 VCC.n422 8.95764
R809 VCC.n912 VCC.n370 8.95764
R810 VCC.n1341 VCC.n974 8.95764
R811 VCC.n1466 VCC.n924 8.95764
R812 VCC.n1899 VCC.n1896 8.95764
R813 VCC.n2021 VCC.n2020 8.95764
R814 VCC.n4 VCC.n3 8.95764
R815 VCC.n282 VCC.n281 8.95764
R816 VCC.n865 VCC.n406 8.85536
R817 VCC.n861 VCC.n406 8.85536
R818 VCC.n1417 VCC.n958 8.85536
R819 VCC.n1413 VCC.n958 8.85536
R820 VCC.n1982 VCC.n1510 8.85536
R821 VCC.n1510 VCC.n1509 8.85536
R822 VCC.n278 VCC.n277 8.85536
R823 VCC.n277 VCC.n276 8.85536
R824 VCC.n661 VCC.n659 8.47776
R825 VCC.n1213 VCC.n1211 8.47776
R826 VCC.n1771 VCC.n1769 8.47776
R827 VCC.n837 VCC.n836 7.03754
R828 VCC.n893 VCC.n371 7.03754
R829 VCC.n1389 VCC.n1388 7.03754
R830 VCC.n1445 VCC.n925 7.03754
R831 VCC.n1946 VCC.n1529 7.03754
R832 VCC.n2018 VCC.n2017 7.03754
R833 VCC.n245 VCC.n244 7.03754
R834 VCC.n301 VCC.n300 7.03754
R835 VCC.n592 VCC.n547 5.48127
R836 VCC.n657 VCC.n656 5.48127
R837 VCC.n703 VCC.n702 5.48127
R838 VCC.n784 VCC.n783 5.48127
R839 VCC.n1144 VCC.n1099 5.48127
R840 VCC.n1209 VCC.n1208 5.48127
R841 VCC.n1255 VCC.n1254 5.48127
R842 VCC.n1336 VCC.n1335 5.48127
R843 VCC.n1812 VCC.n1811 5.48127
R844 VCC.n1893 VCC.n1892 5.48127
R845 VCC.n1702 VCC.n1657 5.48127
R846 VCC.n1767 VCC.n1766 5.48127
R847 VCC.n49 VCC.n48 5.48127
R848 VCC.n15 VCC.n14 5.48127
R849 VCC.n790 VCC.n789 4.88621
R850 VCC.n1342 VCC.n1341 4.88621
R851 VCC.n1900 VCC.n1899 4.88621
R852 VCC.n231 VCC.n4 4.88621
R853 VCC.n865 VCC.n405 4.84621
R854 VCC.n865 VCC.n864 4.84621
R855 VCC.n1417 VCC.n957 4.84621
R856 VCC.n1417 VCC.n1416 4.84621
R857 VCC.n1982 VCC.n1511 4.84621
R858 VCC.n1983 VCC.n1982 4.84621
R859 VCC.n818 VCC.n423 4.6505
R860 VCC.n1370 VCC.n975 4.6505
R861 VCC.n1928 VCC.n1531 4.6505
R862 VCC.n581 VCC.n558 4.51211
R863 VCC.n1133 VCC.n1110 4.51211
R864 VCC.n1691 VCC.n1668 4.51211
R865 VCC.n680 VCC.n491 4.51121
R866 VCC.n1232 VCC.n1043 4.51121
R867 VCC.n1790 VCC.n1600 4.51121
R868 VCC.n667 VCC.n501 4.5005
R869 VCC.n666 VCC.n665 4.5005
R870 VCC.n570 VCC.n569 4.5005
R871 VCC.n566 VCC.n563 4.5005
R872 VCC.n602 VCC.n541 4.5005
R873 VCC.n612 VCC.n611 4.5005
R874 VCC.n613 VCC.n612 4.5005
R875 VCC.n565 VCC.n564 4.5005
R876 VCC.n587 VCC.n540 4.5005
R877 VCC.n587 VCC.n550 4.5005
R878 VCC.n572 VCC.n571 4.5005
R879 VCC.n573 VCC.n572 4.5005
R880 VCC.n617 VCC.n532 4.5005
R881 VCC.n617 VCC.n521 4.5005
R882 VCC.n678 VCC.n677 4.5005
R883 VCC.n642 VCC.n641 4.5005
R884 VCC.n640 VCC.n512 4.5005
R885 VCC.n620 VCC.n533 4.5005
R886 VCC.n628 VCC.n627 4.5005
R887 VCC.n629 VCC.n628 4.5005
R888 VCC.n524 VCC.n514 4.5005
R889 VCC.n525 VCC.n524 4.5005
R890 VCC.n650 VCC.n649 4.5005
R891 VCC.n651 VCC.n650 4.5005
R892 VCC.n669 VCC.n668 4.5005
R893 VCC.n504 VCC.n502 4.5005
R894 VCC.n662 VCC.n504 4.5005
R895 VCC.n605 VCC.n604 4.5005
R896 VCC.n802 VCC.n440 4.5005
R897 VCC.n801 VCC.n800 4.5005
R898 VCC.n695 VCC.n694 4.5005
R899 VCC.n690 VCC.n687 4.5005
R900 VCC.n719 VCC.n718 4.5005
R901 VCC.n689 VCC.n688 4.5005
R902 VCC.n813 VCC.n812 4.5005
R903 VCC.n769 VCC.n768 4.5005
R904 VCC.n767 VCC.n452 4.5005
R905 VCC.n804 VCC.n803 4.5005
R906 VCC.n721 VCC.n720 4.5005
R907 VCC.n734 VCC.n733 4.5005
R908 VCC.n733 VCC.n732 4.5005
R909 VCC.n483 VCC.n479 4.5005
R910 VCC.n706 VCC.n483 4.5005
R911 VCC.n697 VCC.n696 4.5005
R912 VCC.n697 VCC.n490 4.5005
R913 VCC.n749 VCC.n748 4.5005
R914 VCC.n750 VCC.n749 4.5005
R915 VCC.n741 VCC.n462 4.5005
R916 VCC.n752 VCC.n462 4.5005
R917 VCC.n756 VCC.n454 4.5005
R918 VCC.n757 VCC.n756 4.5005
R919 VCC.n777 VCC.n776 4.5005
R920 VCC.n778 VCC.n777 4.5005
R921 VCC.n443 VCC.n441 4.5005
R922 VCC.n797 VCC.n443 4.5005
R923 VCC.n906 VCC.n375 4.5005
R924 VCC.n908 VCC.n907 4.5005
R925 VCC.n885 VCC.n393 4.5005
R926 VCC.n419 VCC.n417 4.5005
R927 VCC.n426 VCC.n424 4.5005
R928 VCC.n817 VCC.n816 4.5005
R929 VCC.n822 VCC.n821 4.5005
R930 VCC.n828 VCC.n416 4.5005
R931 VCC.n414 VCC.n413 4.5005
R932 VCC.n884 VCC.n883 4.5005
R933 VCC.n875 VCC.n397 4.5005
R934 VCC.n887 VCC.n886 4.5005
R935 VCC.n887 VCC.n391 4.5005
R936 VCC.n395 VCC.n382 4.5005
R937 VCC.n383 VCC.n376 4.5005
R938 VCC.n385 VCC.n384 4.5005
R939 VCC.n896 VCC.n385 4.5005
R940 VCC.n874 VCC.n873 4.5005
R941 VCC.n404 VCC.n402 4.5005
R942 VCC.n412 VCC.n410 4.5005
R943 VCC.n410 VCC.n409 4.5005
R944 VCC.n845 VCC.n844 4.5005
R945 VCC.n833 VCC.n832 4.5005
R946 VCC.n820 VCC.n819 4.5005
R947 VCC.n917 VCC.n916 4.5005
R948 VCC.n1219 VCC.n1053 4.5005
R949 VCC.n1218 VCC.n1217 4.5005
R950 VCC.n1122 VCC.n1121 4.5005
R951 VCC.n1118 VCC.n1115 4.5005
R952 VCC.n1154 VCC.n1093 4.5005
R953 VCC.n1164 VCC.n1163 4.5005
R954 VCC.n1165 VCC.n1164 4.5005
R955 VCC.n1117 VCC.n1116 4.5005
R956 VCC.n1139 VCC.n1092 4.5005
R957 VCC.n1139 VCC.n1102 4.5005
R958 VCC.n1124 VCC.n1123 4.5005
R959 VCC.n1125 VCC.n1124 4.5005
R960 VCC.n1169 VCC.n1084 4.5005
R961 VCC.n1169 VCC.n1073 4.5005
R962 VCC.n1230 VCC.n1229 4.5005
R963 VCC.n1194 VCC.n1193 4.5005
R964 VCC.n1192 VCC.n1064 4.5005
R965 VCC.n1172 VCC.n1085 4.5005
R966 VCC.n1180 VCC.n1179 4.5005
R967 VCC.n1181 VCC.n1180 4.5005
R968 VCC.n1076 VCC.n1066 4.5005
R969 VCC.n1077 VCC.n1076 4.5005
R970 VCC.n1202 VCC.n1201 4.5005
R971 VCC.n1203 VCC.n1202 4.5005
R972 VCC.n1221 VCC.n1220 4.5005
R973 VCC.n1056 VCC.n1054 4.5005
R974 VCC.n1214 VCC.n1056 4.5005
R975 VCC.n1157 VCC.n1156 4.5005
R976 VCC.n1354 VCC.n992 4.5005
R977 VCC.n1353 VCC.n1352 4.5005
R978 VCC.n1247 VCC.n1246 4.5005
R979 VCC.n1242 VCC.n1239 4.5005
R980 VCC.n1271 VCC.n1270 4.5005
R981 VCC.n1241 VCC.n1240 4.5005
R982 VCC.n1365 VCC.n1364 4.5005
R983 VCC.n1321 VCC.n1320 4.5005
R984 VCC.n1319 VCC.n1004 4.5005
R985 VCC.n1356 VCC.n1355 4.5005
R986 VCC.n1273 VCC.n1272 4.5005
R987 VCC.n1286 VCC.n1285 4.5005
R988 VCC.n1285 VCC.n1284 4.5005
R989 VCC.n1035 VCC.n1031 4.5005
R990 VCC.n1258 VCC.n1035 4.5005
R991 VCC.n1249 VCC.n1248 4.5005
R992 VCC.n1249 VCC.n1042 4.5005
R993 VCC.n1301 VCC.n1300 4.5005
R994 VCC.n1302 VCC.n1301 4.5005
R995 VCC.n1293 VCC.n1014 4.5005
R996 VCC.n1304 VCC.n1014 4.5005
R997 VCC.n1308 VCC.n1006 4.5005
R998 VCC.n1309 VCC.n1308 4.5005
R999 VCC.n1329 VCC.n1328 4.5005
R1000 VCC.n1330 VCC.n1329 4.5005
R1001 VCC.n995 VCC.n993 4.5005
R1002 VCC.n1349 VCC.n995 4.5005
R1003 VCC.n935 VCC.n930 4.5005
R1004 VCC.n1462 VCC.n1461 4.5005
R1005 VCC.n1372 VCC.n1371 4.5005
R1006 VCC.n978 VCC.n976 4.5005
R1007 VCC.n1397 VCC.n1396 4.5005
R1008 VCC.n964 VCC.n962 4.5005
R1009 VCC.n962 VCC.n961 4.5005
R1010 VCC.n966 VCC.n965 4.5005
R1011 VCC.n1380 VCC.n968 4.5005
R1012 VCC.n1385 VCC.n1384 4.5005
R1013 VCC.n1369 VCC.n1368 4.5005
R1014 VCC.n1374 VCC.n1373 4.5005
R1015 VCC.n937 VCC.n936 4.5005
R1016 VCC.n1448 VCC.n937 4.5005
R1017 VCC.n1436 VCC.n1435 4.5005
R1018 VCC.n947 VCC.n934 4.5005
R1019 VCC.n1426 VCC.n1425 4.5005
R1020 VCC.n956 VCC.n954 4.5005
R1021 VCC.n1427 VCC.n949 4.5005
R1022 VCC.n1437 VCC.n945 4.5005
R1023 VCC.n1439 VCC.n1438 4.5005
R1024 VCC.n1439 VCC.n943 4.5005
R1025 VCC.n1460 VCC.n929 4.5005
R1026 VCC.n1471 VCC.n1470 4.5005
R1027 VCC.n971 VCC.n969 4.5005
R1028 VCC.n1930 VCC.n1532 4.5005
R1029 VCC.n1933 VCC.n1932 4.5005
R1030 VCC.n2007 VCC.n1487 4.5005
R1031 VCC.n2009 VCC.n2008 4.5005
R1032 VCC.n1504 VCC.n1503 4.5005
R1033 VCC.n1524 VCC.n1522 4.5005
R1034 VCC.n1534 VCC.n1521 4.5005
R1035 VCC.n1963 VCC.n1962 4.5005
R1036 VCC.n1972 VCC.n1971 4.5005
R1037 VCC.n1515 VCC.n1514 4.5005
R1038 VCC.n1495 VCC.n1494 4.5005
R1039 VCC.n1998 VCC.n1997 4.5005
R1040 VCC.n2010 VCC.n1485 4.5005
R1041 VCC.n1499 VCC.n1497 4.5005
R1042 VCC.n1970 VCC.n1969 4.5005
R1043 VCC.n1931 VCC.n1929 4.5005
R1044 VCC.n1927 VCC.n1926 4.5005
R1045 VCC.n1942 VCC.n1533 4.5005
R1046 VCC.n2012 VCC.n2011 4.5005
R1047 VCC.n2012 VCC.n1483 4.5005
R1048 VCC.n1502 VCC.n1500 4.5005
R1049 VCC.n1507 VCC.n1500 4.5005
R1050 VCC.n1958 VCC.n1957 4.5005
R1051 VCC.n1959 VCC.n1958 4.5005
R1052 VCC.n2025 VCC.n2024 4.5005
R1053 VCC.n1912 VCC.n1549 4.5005
R1054 VCC.n1911 VCC.n1910 4.5005
R1055 VCC.n1876 VCC.n1561 4.5005
R1056 VCC.n1830 VCC.n1829 4.5005
R1057 VCC.n1804 VCC.n1803 4.5005
R1058 VCC.n1799 VCC.n1795 4.5005
R1059 VCC.n1805 VCC.n1601 4.5005
R1060 VCC.n1601 VCC.n1599 4.5005
R1061 VCC.n1923 VCC.n1922 4.5005
R1062 VCC.n1878 VCC.n1877 4.5005
R1063 VCC.n1798 VCC.n1797 4.5005
R1064 VCC.n1592 VCC.n1588 4.5005
R1065 VCC.n1815 VCC.n1592 4.5005
R1066 VCC.n1828 VCC.n1827 4.5005
R1067 VCC.n1843 VCC.n1842 4.5005
R1068 VCC.n1842 VCC.n1841 4.5005
R1069 VCC.n1858 VCC.n1857 4.5005
R1070 VCC.n1859 VCC.n1858 4.5005
R1071 VCC.n1850 VCC.n1571 4.5005
R1072 VCC.n1861 VCC.n1571 4.5005
R1073 VCC.n1865 VCC.n1563 4.5005
R1074 VCC.n1866 VCC.n1865 4.5005
R1075 VCC.n1886 VCC.n1885 4.5005
R1076 VCC.n1887 VCC.n1886 4.5005
R1077 VCC.n1914 VCC.n1913 4.5005
R1078 VCC.n1552 VCC.n1550 4.5005
R1079 VCC.n1907 VCC.n1552 4.5005
R1080 VCC.n1777 VCC.n1611 4.5005
R1081 VCC.n1776 VCC.n1775 4.5005
R1082 VCC.n1750 VCC.n1622 4.5005
R1083 VCC.n1715 VCC.n1714 4.5005
R1084 VCC.n1680 VCC.n1679 4.5005
R1085 VCC.n1676 VCC.n1673 4.5005
R1086 VCC.n1682 VCC.n1681 4.5005
R1087 VCC.n1683 VCC.n1682 4.5005
R1088 VCC.n1788 VCC.n1787 4.5005
R1089 VCC.n1752 VCC.n1751 4.5005
R1090 VCC.n1675 VCC.n1674 4.5005
R1091 VCC.n1697 VCC.n1650 4.5005
R1092 VCC.n1697 VCC.n1660 4.5005
R1093 VCC.n1712 VCC.n1651 4.5005
R1094 VCC.n1722 VCC.n1721 4.5005
R1095 VCC.n1723 VCC.n1722 4.5005
R1096 VCC.n1727 VCC.n1642 4.5005
R1097 VCC.n1727 VCC.n1631 4.5005
R1098 VCC.n1730 VCC.n1643 4.5005
R1099 VCC.n1738 VCC.n1737 4.5005
R1100 VCC.n1739 VCC.n1738 4.5005
R1101 VCC.n1634 VCC.n1624 4.5005
R1102 VCC.n1635 VCC.n1634 4.5005
R1103 VCC.n1760 VCC.n1759 4.5005
R1104 VCC.n1761 VCC.n1760 4.5005
R1105 VCC.n1779 VCC.n1778 4.5005
R1106 VCC.n1614 VCC.n1612 4.5005
R1107 VCC.n1772 VCC.n1614 4.5005
R1108 VCC.n76 VCC.n75 4.5005
R1109 VCC.n56 VCC.n55 4.5005
R1110 VCC.n35 VCC.n34 4.5005
R1111 VCC.n82 VCC.n81 4.5005
R1112 VCC.n187 VCC.n186 4.5005
R1113 VCC.n201 VCC.n200 4.5005
R1114 VCC.n222 VCC.n221 4.5005
R1115 VCC.n269 VCC.n268 4.5005
R1116 VCC.n307 VCC.n306 4.5005
R1117 VCC.n326 VCC.n325 4.5005
R1118 VCC.n914 VCC.n370 4.31039
R1119 VCC.n1468 VCC.n924 4.31039
R1120 VCC.n2021 VCC.n1477 4.31039
R1121 VCC.n284 VCC.n282 4.31039
R1122 VCC.n838 VCC.n407 3.51902
R1123 VCC.n891 VCC.n388 3.51902
R1124 VCC.n1390 VCC.n959 3.51902
R1125 VCC.n1443 VCC.n940 3.51902
R1126 VCC.n1951 VCC.n1950 3.51902
R1127 VCC.n1987 VCC.n1986 3.51902
R1128 VCC.n265 VCC.n264 3.51902
R1129 VCC.n321 VCC.n320 3.51902
R1130 VCC.n679 VCC.n678 3.42479
R1131 VCC.n681 VCC.n680 3.42479
R1132 VCC.n1231 VCC.n1230 3.42479
R1133 VCC.n1233 VCC.n1232 3.42479
R1134 VCC.n1791 VCC.n1790 3.42479
R1135 VCC.n1789 VCC.n1788 3.42479
R1136 VCC.n558 VCC.n557 3.42389
R1137 VCC.n814 VCC.n813 3.42389
R1138 VCC.n816 VCC.n815 3.42389
R1139 VCC.n1110 VCC.n1109 3.42389
R1140 VCC.n1366 VCC.n1365 3.42389
R1141 VCC.n1368 VCC.n1367 3.42389
R1142 VCC.n1926 VCC.n1925 3.42389
R1143 VCC.n1924 VCC.n1923 3.42389
R1144 VCC.n1668 VCC.n1667 3.42389
R1145 VCC.n918 VCC.n917 3.423
R1146 VCC.n1472 VCC.n1471 3.423
R1147 VCC.n2026 VCC.n2025 3.423
R1148 VCC.n880 VCC.n879 3.4105
R1149 VCC.n902 VCC.n901 3.4105
R1150 VCC.n901 VCC.n900 3.4105
R1151 VCC.n870 VCC.n399 3.4105
R1152 VCC.n399 VCC.n398 3.4105
R1153 VCC.n872 VCC.n871 3.4105
R1154 VCC.n878 VCC.n877 3.4105
R1155 VCC.n877 VCC.n876 3.4105
R1156 VCC.n852 VCC.n851 3.4105
R1157 VCC.n852 VCC.n411 3.4105
R1158 VCC.n848 VCC.n401 3.4105
R1159 VCC.n869 VCC.n868 3.4105
R1160 VCC.n868 VCC.n867 3.4105
R1161 VCC.n830 VCC.n827 3.4105
R1162 VCC.n830 VCC.n829 3.4105
R1163 VCC.n847 VCC.n846 3.4105
R1164 VCC.n810 VCC.n809 3.4105
R1165 VCC.n811 VCC.n810 3.4105
R1166 VCC.n775 VCC.n774 3.4105
R1167 VCC.n808 VCC.n807 3.4105
R1168 VCC.n807 VCC.n806 3.4105
R1169 VCC.n745 VCC.n744 3.4105
R1170 VCC.n744 VCC.n743 3.4105
R1171 VCC.n740 VCC.n738 3.4105
R1172 VCC.n773 VCC.n772 3.4105
R1173 VCC.n772 VCC.n771 3.4105
R1174 VCC.n469 VCC.n468 3.4105
R1175 VCC.n716 VCC.n469 3.4105
R1176 VCC.n737 VCC.n466 3.4105
R1177 VCC.n747 VCC.n746 3.4105
R1178 VCC.n747 VCC.n465 3.4105
R1179 VCC.n710 VCC.n480 3.4105
R1180 VCC.n710 VCC.n709 3.4105
R1181 VCC.n714 VCC.n713 3.4105
R1182 VCC.n684 VCC.n683 3.4105
R1183 VCC.n684 VCC.n491 3.4105
R1184 VCC.n675 VCC.n674 3.4105
R1185 VCC.n676 VCC.n675 3.4105
R1186 VCC.n648 VCC.n647 3.4105
R1187 VCC.n673 VCC.n672 3.4105
R1188 VCC.n672 VCC.n671 3.4105
R1189 VCC.n624 VCC.n529 3.4105
R1190 VCC.n529 VCC.n523 3.4105
R1191 VCC.n626 VCC.n625 3.4105
R1192 VCC.n646 VCC.n645 3.4105
R1193 VCC.n645 VCC.n644 3.4105
R1194 VCC.n608 VCC.n537 3.4105
R1195 VCC.n537 VCC.n536 3.4105
R1196 VCC.n538 VCC.n531 3.4105
R1197 VCC.n623 VCC.n622 3.4105
R1198 VCC.n622 VCC.n621 3.4105
R1199 VCC.n585 VCC.n584 3.4105
R1200 VCC.n586 VCC.n585 3.4105
R1201 VCC.n607 VCC.n606 3.4105
R1202 VCC.n583 VCC.n582 3.4105
R1203 VCC.n582 VCC.n581 3.4105
R1204 VCC.n826 VCC.n825 3.4105
R1205 VCC.n825 VCC.n824 3.4105
R1206 VCC.n904 VCC.n903 3.4105
R1207 VCC.n904 VCC.n368 3.4105
R1208 VCC.n1456 VCC.n1455 3.4105
R1209 VCC.n1456 VCC.n922 3.4105
R1210 VCC.n1432 VCC.n1431 3.4105
R1211 VCC.n1454 VCC.n1453 3.4105
R1212 VCC.n1453 VCC.n1452 3.4105
R1213 VCC.n1422 VCC.n951 3.4105
R1214 VCC.n951 VCC.n950 3.4105
R1215 VCC.n1424 VCC.n1423 3.4105
R1216 VCC.n1430 VCC.n1429 3.4105
R1217 VCC.n1429 VCC.n1428 3.4105
R1218 VCC.n1404 VCC.n1403 3.4105
R1219 VCC.n1404 VCC.n963 3.4105
R1220 VCC.n1400 VCC.n953 3.4105
R1221 VCC.n1421 VCC.n1420 3.4105
R1222 VCC.n1420 VCC.n1419 3.4105
R1223 VCC.n1382 VCC.n1379 3.4105
R1224 VCC.n1382 VCC.n1381 3.4105
R1225 VCC.n1399 VCC.n1398 3.4105
R1226 VCC.n1378 VCC.n1377 3.4105
R1227 VCC.n1377 VCC.n1376 3.4105
R1228 VCC.n1362 VCC.n1361 3.4105
R1229 VCC.n1363 VCC.n1362 3.4105
R1230 VCC.n1327 VCC.n1326 3.4105
R1231 VCC.n1360 VCC.n1359 3.4105
R1232 VCC.n1359 VCC.n1358 3.4105
R1233 VCC.n1297 VCC.n1296 3.4105
R1234 VCC.n1296 VCC.n1295 3.4105
R1235 VCC.n1292 VCC.n1290 3.4105
R1236 VCC.n1325 VCC.n1324 3.4105
R1237 VCC.n1324 VCC.n1323 3.4105
R1238 VCC.n1021 VCC.n1020 3.4105
R1239 VCC.n1268 VCC.n1021 3.4105
R1240 VCC.n1289 VCC.n1018 3.4105
R1241 VCC.n1299 VCC.n1298 3.4105
R1242 VCC.n1299 VCC.n1017 3.4105
R1243 VCC.n1262 VCC.n1032 3.4105
R1244 VCC.n1262 VCC.n1261 3.4105
R1245 VCC.n1266 VCC.n1265 3.4105
R1246 VCC.n1236 VCC.n1235 3.4105
R1247 VCC.n1236 VCC.n1043 3.4105
R1248 VCC.n1227 VCC.n1226 3.4105
R1249 VCC.n1228 VCC.n1227 3.4105
R1250 VCC.n1200 VCC.n1199 3.4105
R1251 VCC.n1225 VCC.n1224 3.4105
R1252 VCC.n1224 VCC.n1223 3.4105
R1253 VCC.n1176 VCC.n1081 3.4105
R1254 VCC.n1081 VCC.n1075 3.4105
R1255 VCC.n1178 VCC.n1177 3.4105
R1256 VCC.n1198 VCC.n1197 3.4105
R1257 VCC.n1197 VCC.n1196 3.4105
R1258 VCC.n1160 VCC.n1089 3.4105
R1259 VCC.n1089 VCC.n1088 3.4105
R1260 VCC.n1090 VCC.n1083 3.4105
R1261 VCC.n1175 VCC.n1174 3.4105
R1262 VCC.n1174 VCC.n1173 3.4105
R1263 VCC.n1137 VCC.n1136 3.4105
R1264 VCC.n1138 VCC.n1137 3.4105
R1265 VCC.n1159 VCC.n1158 3.4105
R1266 VCC.n1135 VCC.n1134 3.4105
R1267 VCC.n1134 VCC.n1133 3.4105
R1268 VCC.n1785 VCC.n1784 3.4105
R1269 VCC.n1786 VCC.n1785 3.4105
R1270 VCC.n1758 VCC.n1757 3.4105
R1271 VCC.n1783 VCC.n1782 3.4105
R1272 VCC.n1782 VCC.n1781 3.4105
R1273 VCC.n1734 VCC.n1639 3.4105
R1274 VCC.n1639 VCC.n1633 3.4105
R1275 VCC.n1736 VCC.n1735 3.4105
R1276 VCC.n1756 VCC.n1755 3.4105
R1277 VCC.n1755 VCC.n1754 3.4105
R1278 VCC.n1718 VCC.n1647 3.4105
R1279 VCC.n1647 VCC.n1646 3.4105
R1280 VCC.n1648 VCC.n1641 3.4105
R1281 VCC.n1733 VCC.n1732 3.4105
R1282 VCC.n1732 VCC.n1731 3.4105
R1283 VCC.n1695 VCC.n1694 3.4105
R1284 VCC.n1696 VCC.n1695 3.4105
R1285 VCC.n1717 VCC.n1716 3.4105
R1286 VCC.n1693 VCC.n1692 3.4105
R1287 VCC.n1692 VCC.n1691 3.4105
R1288 VCC.n1937 VCC.n1936 3.4105
R1289 VCC.n1936 VCC.n1935 3.4105
R1290 VCC.n1996 VCC.n1995 3.4105
R1291 VCC.n2001 VCC.n2000 3.4105
R1292 VCC.n2000 VCC.n1999 3.4105
R1293 VCC.n1979 VCC.n1978 3.4105
R1294 VCC.n1980 VCC.n1979 3.4105
R1295 VCC.n1977 VCC.n1976 3.4105
R1296 VCC.n1994 VCC.n1993 3.4105
R1297 VCC.n1993 VCC.n1992 3.4105
R1298 VCC.n1966 VCC.n1519 3.4105
R1299 VCC.n1519 VCC.n1518 3.4105
R1300 VCC.n1517 VCC.n1516 3.4105
R1301 VCC.n1974 VCC.n1973 3.4105
R1302 VCC.n1973 VCC.n1512 3.4105
R1303 VCC.n1939 VCC.n1938 3.4105
R1304 VCC.n1939 VCC.n1535 3.4105
R1305 VCC.n1965 VCC.n1964 3.4105
R1306 VCC.n2003 VCC.n2002 3.4105
R1307 VCC.n2003 VCC.n1476 3.4105
R1308 VCC.n1920 VCC.n1919 3.4105
R1309 VCC.n1921 VCC.n1920 3.4105
R1310 VCC.n1884 VCC.n1883 3.4105
R1311 VCC.n1918 VCC.n1917 3.4105
R1312 VCC.n1917 VCC.n1916 3.4105
R1313 VCC.n1854 VCC.n1853 3.4105
R1314 VCC.n1853 VCC.n1852 3.4105
R1315 VCC.n1849 VCC.n1847 3.4105
R1316 VCC.n1882 VCC.n1881 3.4105
R1317 VCC.n1881 VCC.n1880 3.4105
R1318 VCC.n1578 VCC.n1577 3.4105
R1319 VCC.n1825 VCC.n1578 3.4105
R1320 VCC.n1846 VCC.n1575 3.4105
R1321 VCC.n1856 VCC.n1855 3.4105
R1322 VCC.n1856 VCC.n1574 3.4105
R1323 VCC.n1819 VCC.n1589 3.4105
R1324 VCC.n1819 VCC.n1818 3.4105
R1325 VCC.n1823 VCC.n1822 3.4105
R1326 VCC.n1794 VCC.n1793 3.4105
R1327 VCC.n1794 VCC.n1600 3.4105
R1328 VCC.n787 VCC.n423 3.29193
R1329 VCC.n842 VCC.n841 3.29193
R1330 VCC.n881 VCC.n386 3.29193
R1331 VCC.n1339 VCC.n975 3.29193
R1332 VCC.n1394 VCC.n1393 3.29193
R1333 VCC.n1433 VCC.n938 3.29193
R1334 VCC.n1897 VCC.n1531 3.29193
R1335 VCC.n1960 VCC.n1525 3.29193
R1336 VCC.n1506 VCC.n1482 3.29193
R1337 VCC.n835 VCC.n421 3.25764
R1338 VCC.n894 VCC.n372 3.25764
R1339 VCC.n1387 VCC.n973 3.25764
R1340 VCC.n1446 VCC.n926 3.25764
R1341 VCC.n1945 VCC.n1530 3.25764
R1342 VCC.n2016 VCC.n1479 3.25764
R1343 VCC.n246 VCC.n242 3.25764
R1344 VCC.n302 VCC.n298 3.25764
R1345 VCC.n911 VCC.n910 3.2005
R1346 VCC.n1465 VCC.n1464 3.2005
R1347 VCC.n1490 VCC.n1478 3.2005
R1348 VCC.n866 VCC.n865 3.03311
R1349 VCC.n834 VCC.n833 3.03311
R1350 VCC.n1386 VCC.n1385 3.03311
R1351 VCC.n1418 VCC.n1417 3.03311
R1352 VCC.n1982 VCC.n1981 3.03311
R1353 VCC.n1943 VCC.n1942 3.03311
R1354 VCC.n250 VCC.n249 3.03311
R1355 VCC.n333 VCC.n278 3.03311
R1356 VCC.n591 VCC.n548 2.8505
R1357 VCC.n658 VCC.n506 2.8505
R1358 VCC.n704 VCC.n485 2.8505
R1359 VCC.n782 VCC.n446 2.8505
R1360 VCC.n1143 VCC.n1100 2.8505
R1361 VCC.n1210 VCC.n1058 2.8505
R1362 VCC.n1256 VCC.n1037 2.8505
R1363 VCC.n1334 VCC.n998 2.8505
R1364 VCC.n1813 VCC.n1594 2.8505
R1365 VCC.n1891 VCC.n1555 2.8505
R1366 VCC.n1701 VCC.n1658 2.8505
R1367 VCC.n1768 VCC.n1616 2.8505
R1368 VCC.n47 VCC.n46 2.8505
R1369 VCC.n13 VCC.n12 2.8505
R1370 VCC.n638 VCC.n637 2.5605
R1371 VCC.n765 VCC.n764 2.5605
R1372 VCC.n1190 VCC.n1189 2.5605
R1373 VCC.n1317 VCC.n1316 2.5605
R1374 VCC.n1874 VCC.n1873 2.5605
R1375 VCC.n1748 VCC.n1747 2.5605
R1376 VCC.n9 VCC.n8 2.5605
R1377 VCC.n598 VCC.n597 2.46907
R1378 VCC.n724 VCC.n723 2.46907
R1379 VCC.n1150 VCC.n1149 2.46907
R1380 VCC.n1276 VCC.n1275 2.46907
R1381 VCC.n1833 VCC.n1832 2.46907
R1382 VCC.n1708 VCC.n1707 2.46907
R1383 VCC.n507 VCC.n505 2.37764
R1384 VCC.n780 VCC.n444 2.37764
R1385 VCC.n1059 VCC.n1057 2.37764
R1386 VCC.n1332 VCC.n996 2.37764
R1387 VCC.n1889 VCC.n1553 2.37764
R1388 VCC.n1617 VCC.n1615 2.37764
R1389 VCC.n21 VCC.n20 2.37764
R1390 VCC.n574 VCC.n560 2.34304
R1391 VCC.n447 VCC.n445 2.34304
R1392 VCC.n489 VCC.n487 2.34304
R1393 VCC.n1126 VCC.n1112 2.34304
R1394 VCC.n999 VCC.n997 2.34304
R1395 VCC.n1041 VCC.n1039 2.34304
R1396 VCC.n1556 VCC.n1554 2.34304
R1397 VCC.n1598 VCC.n1596 2.34304
R1398 VCC.n1684 VCC.n1670 2.34304
R1399 VCC.n6 VCC.n5 2.34304
R1400 VCC.n26 VCC.n25 2.34304
R1401 VCC.n2028 VCC.n1473 2.29829
R1402 VCC.n567 VCC.n549 2.28621
R1403 VCC.n692 VCC.n484 2.28621
R1404 VCC.n1119 VCC.n1101 2.28621
R1405 VCC.n1244 VCC.n1036 2.28621
R1406 VCC.n1801 VCC.n1593 2.28621
R1407 VCC.n1677 VCC.n1659 2.28621
R1408 VCC.n496 VCC.n495 2.2505
R1409 VCC.n670 VCC.n499 2.2505
R1410 VCC.n643 VCC.n515 2.2505
R1411 VCC.n559 VCC.n556 2.2505
R1412 VCC.n552 VCC.n551 2.2505
R1413 VCC.n601 VCC.n600 2.2505
R1414 VCC.n435 VCC.n434 2.2505
R1415 VCC.n805 VCC.n438 2.2505
R1416 VCC.n770 VCC.n455 2.2505
R1417 VCC.n698 VCC.n685 2.2505
R1418 VCC.n482 VCC.n481 2.2505
R1419 VCC.n717 VCC.n715 2.2505
R1420 VCC.n905 VCC.n378 2.2505
R1421 VCC.n831 VCC.n425 2.2505
R1422 VCC.n854 VCC.n853 2.2505
R1423 VCC.n394 VCC.n392 2.2505
R1424 VCC.n899 VCC.n381 2.2505
R1425 VCC.n823 VCC.n430 2.2505
R1426 VCC.n1048 VCC.n1047 2.2505
R1427 VCC.n1222 VCC.n1051 2.2505
R1428 VCC.n1195 VCC.n1067 2.2505
R1429 VCC.n1111 VCC.n1108 2.2505
R1430 VCC.n1104 VCC.n1103 2.2505
R1431 VCC.n1153 VCC.n1152 2.2505
R1432 VCC.n987 VCC.n986 2.2505
R1433 VCC.n1357 VCC.n990 2.2505
R1434 VCC.n1322 VCC.n1007 2.2505
R1435 VCC.n1250 VCC.n1237 2.2505
R1436 VCC.n1034 VCC.n1033 2.2505
R1437 VCC.n1269 VCC.n1267 2.2505
R1438 VCC.n1459 VCC.n1458 2.2505
R1439 VCC.n1451 VCC.n933 2.2505
R1440 VCC.n946 VCC.n944 2.2505
R1441 VCC.n1375 VCC.n982 2.2505
R1442 VCC.n1383 VCC.n977 2.2505
R1443 VCC.n1406 VCC.n1405 2.2505
R1444 VCC.n2005 VCC.n2004 2.2505
R1445 VCC.n1956 VCC.n1955 2.2505
R1446 VCC.n1486 VCC.n1484 2.2505
R1447 VCC.n1991 VCC.n1498 2.2505
R1448 VCC.n1941 VCC.n1940 2.2505
R1449 VCC.n1934 VCC.n1539 2.2505
R1450 VCC.n1544 VCC.n1543 2.2505
R1451 VCC.n1915 VCC.n1547 2.2505
R1452 VCC.n1879 VCC.n1564 2.2505
R1453 VCC.n1826 VCC.n1824 2.2505
R1454 VCC.n1591 VCC.n1590 2.2505
R1455 VCC.n1807 VCC.n1806 2.2505
R1456 VCC.n1606 VCC.n1605 2.2505
R1457 VCC.n1780 VCC.n1609 2.2505
R1458 VCC.n1753 VCC.n1625 2.2505
R1459 VCC.n1711 VCC.n1710 2.2505
R1460 VCC.n1662 VCC.n1661 2.2505
R1461 VCC.n1669 VCC.n1666 2.2505
R1462 VCC VCC.n2028 2.24163
R1463 VCC.n630 VCC.n629 2.10336
R1464 VCC.n752 VCC.n751 2.10336
R1465 VCC.n1182 VCC.n1181 2.10336
R1466 VCC.n1304 VCC.n1303 2.10336
R1467 VCC.n1861 VCC.n1860 2.10336
R1468 VCC.n1740 VCC.n1739 2.10336
R1469 VCC.n630 VCC.n521 2.01193
R1470 VCC.n751 VCC.n750 2.01193
R1471 VCC.n1182 VCC.n1073 2.01193
R1472 VCC.n1303 VCC.n1302 2.01193
R1473 VCC.n1860 VCC.n1859 2.01193
R1474 VCC.n1740 VCC.n1631 2.01193
R1475 VCC.n81 VCC.n80 2.01193
R1476 VCC.n916 VCC.n915 2.00996
R1477 VCC.n1470 VCC.n1469 2.00996
R1478 VCC.n2024 VCC.n2023 2.00996
R1479 VCC.n286 VCC.n285 2.00996
R1480 VCC.n817 VCC.n431 1.98102
R1481 VCC.n1369 VCC.n983 1.98102
R1482 VCC.n233 VCC.n232 1.98102
R1483 VCC.n1927 VCC.n1540 1.98071
R1484 VCC.n1473 VCC 1.87918
R1485 VCC.n595 VCC.n594 1.82742
R1486 VCC.n634 VCC.n508 1.82742
R1487 VCC.n727 VCC.n726 1.82742
R1488 VCC.n762 VCC.n761 1.82742
R1489 VCC.n1147 VCC.n1146 1.82742
R1490 VCC.n1186 VCC.n1060 1.82742
R1491 VCC.n1279 VCC.n1278 1.82742
R1492 VCC.n1314 VCC.n1313 1.82742
R1493 VCC.n1836 VCC.n1835 1.82742
R1494 VCC.n1871 VCC.n1870 1.82742
R1495 VCC.n1705 VCC.n1704 1.82742
R1496 VCC.n1744 VCC.n1618 1.82742
R1497 VCC.n70 VCC.n69 1.82742
R1498 VCC.n196 VCC.n195 1.82742
R1499 VCC.n858 VCC.n408 1.62907
R1500 VCC.n890 VCC.n389 1.62907
R1501 VCC.n1410 VCC.n960 1.62907
R1502 VCC.n1442 VCC.n941 1.62907
R1503 VCC.n1952 VCC.n1528 1.62907
R1504 VCC.n1988 VCC.n1508 1.62907
R1505 VCC.n266 VCC.n262 1.62907
R1506 VCC.n322 VCC.n318 1.62907
R1507 VCC.n834 VCC.n423 1.55479
R1508 VCC.n1386 VCC.n975 1.55479
R1509 VCC.n1943 VCC.n1531 1.55479
R1510 VCC.n249 VCC.n240 1.55479
R1511 VCC.n619 VCC.n618 1.5005
R1512 VCC.n1171 VCC.n1170 1.5005
R1513 VCC.n1729 VCC.n1728 1.5005
R1514 VCC.n544 VCC.n535 1.46336
R1515 VCC.n636 VCC.n517 1.46336
R1516 VCC.n730 VCC.n472 1.46336
R1517 VCC.n758 VCC.n457 1.46336
R1518 VCC.n896 VCC.n373 1.46336
R1519 VCC.n1096 VCC.n1087 1.46336
R1520 VCC.n1188 VCC.n1069 1.46336
R1521 VCC.n1282 VCC.n1024 1.46336
R1522 VCC.n1310 VCC.n1009 1.46336
R1523 VCC.n1448 VCC.n927 1.46336
R1524 VCC.n1489 VCC.n1483 1.46336
R1525 VCC.n1839 VCC.n1581 1.46336
R1526 VCC.n1867 VCC.n1566 1.46336
R1527 VCC.n1654 VCC.n1645 1.46336
R1528 VCC.n1746 VCC.n1627 1.46336
R1529 VCC.n73 VCC.n66 1.46336
R1530 VCC.n306 VCC.n305 1.46336
R1531 VCC.n842 VCC.n409 1.37193
R1532 VCC.n857 VCC.n405 1.37193
R1533 VCC.n864 VCC.n390 1.37193
R1534 VCC.n881 VCC.n391 1.37193
R1535 VCC.n1394 VCC.n961 1.37193
R1536 VCC.n1409 VCC.n957 1.37193
R1537 VCC.n1416 VCC.n942 1.37193
R1538 VCC.n1433 VCC.n943 1.37193
R1539 VCC.n1960 VCC.n1959 1.37193
R1540 VCC.n1526 VCC.n1511 1.37193
R1541 VCC.n1983 VCC.n1501 1.37193
R1542 VCC.n1507 VCC.n1506 1.37193
R1543 VCC.n268 VCC.n258 1.37193
R1544 VCC.n260 VCC.n259 1.37193
R1545 VCC.n316 VCC.n315 1.37193
R1546 VCC.n325 VCC.n324 1.37193
R1547 VCC.n590 VCC.n589 1.2805
R1548 VCC.n653 VCC.n652 1.2805
R1549 VCC.n707 VCC.n705 1.2805
R1550 VCC.n781 VCC.n779 1.2805
R1551 VCC.n1142 VCC.n1141 1.2805
R1552 VCC.n1205 VCC.n1204 1.2805
R1553 VCC.n1259 VCC.n1257 1.2805
R1554 VCC.n1333 VCC.n1331 1.2805
R1555 VCC.n1816 VCC.n1814 1.2805
R1556 VCC.n1890 VCC.n1888 1.2805
R1557 VCC.n1700 VCC.n1699 1.2805
R1558 VCC.n1763 VCC.n1762 1.2805
R1559 VCC.n52 VCC.n45 1.2805
R1560 VCC.n19 VCC.n18 1.2805
R1561 VCC.n841 VCC.n420 1.18907
R1562 VCC.n895 VCC.n386 1.18907
R1563 VCC.n1393 VCC.n972 1.18907
R1564 VCC.n1447 VCC.n938 1.18907
R1565 VCC.n1944 VCC.n1525 1.18907
R1566 VCC.n2015 VCC.n1482 1.18907
R1567 VCC.n248 VCC.n247 1.18907
R1568 VCC.n296 VCC.n295 1.18907
R1569 VCC.n367 VCC.n366 1.13717
R1570 VCC.n555 VCC.n554 1.13717
R1571 VCC.n553 VCC.n539 1.13717
R1572 VCC.n610 VCC.n609 1.13717
R1573 VCC.n530 VCC.n513 1.13717
R1574 VCC.n498 VCC.n497 1.13717
R1575 VCC.n494 VCC.n493 1.13717
R1576 VCC.n682 VCC.n492 1.13717
R1577 VCC.n712 VCC.n711 1.13717
R1578 VCC.n736 VCC.n735 1.13717
R1579 VCC.n739 VCC.n453 1.13717
R1580 VCC.n437 VCC.n436 1.13717
R1581 VCC.n433 VCC.n432 1.13717
R1582 VCC.n429 VCC.n428 1.13717
R1583 VCC.n427 VCC.n415 1.13717
R1584 VCC.n850 VCC.n849 1.13717
R1585 VCC.n400 VCC.n396 1.13717
R1586 VCC.n380 VCC.n379 1.13717
R1587 VCC.n1107 VCC.n1106 1.13717
R1588 VCC.n1105 VCC.n1091 1.13717
R1589 VCC.n1162 VCC.n1161 1.13717
R1590 VCC.n1082 VCC.n1065 1.13717
R1591 VCC.n1050 VCC.n1049 1.13717
R1592 VCC.n1046 VCC.n1045 1.13717
R1593 VCC.n1234 VCC.n1044 1.13717
R1594 VCC.n1264 VCC.n1263 1.13717
R1595 VCC.n1288 VCC.n1287 1.13717
R1596 VCC.n1291 VCC.n1005 1.13717
R1597 VCC.n989 VCC.n988 1.13717
R1598 VCC.n985 VCC.n984 1.13717
R1599 VCC.n981 VCC.n980 1.13717
R1600 VCC.n979 VCC.n967 1.13717
R1601 VCC.n1402 VCC.n1401 1.13717
R1602 VCC.n952 VCC.n948 1.13717
R1603 VCC.n932 VCC.n931 1.13717
R1604 VCC.n921 VCC.n920 1.13717
R1605 VCC.n1665 VCC.n1664 1.13717
R1606 VCC.n1663 VCC.n1649 1.13717
R1607 VCC.n1720 VCC.n1719 1.13717
R1608 VCC.n1640 VCC.n1623 1.13717
R1609 VCC.n1608 VCC.n1607 1.13717
R1610 VCC.n1604 VCC.n1603 1.13717
R1611 VCC.n1792 VCC.n1602 1.13717
R1612 VCC.n1536 VCC.n1520 1.13717
R1613 VCC.n1968 VCC.n1967 1.13717
R1614 VCC.n1975 VCC.n1496 1.13717
R1615 VCC.n1493 VCC.n1492 1.13717
R1616 VCC.n1475 VCC.n1474 1.13717
R1617 VCC.n1538 VCC.n1537 1.13717
R1618 VCC.n1821 VCC.n1820 1.13717
R1619 VCC.n1845 VCC.n1844 1.13717
R1620 VCC.n1848 VCC.n1562 1.13717
R1621 VCC.n1546 VCC.n1545 1.13717
R1622 VCC.n1542 VCC.n1541 1.13717
R1623 VCC.n112 VCC.n111 1.13717
R1624 VCC.n178 VCC.n177 1.13717
R1625 VCC.n168 VCC.n167 1.13717
R1626 VCC.n160 VCC.n159 1.13717
R1627 VCC.n149 VCC.n148 1.13717
R1628 VCC.n342 VCC.n341 1.13717
R1629 VCC.n354 VCC.n353 1.13717
R1630 VCC.n364 VCC.n363 1.13717
R1631 VCC.n742 VCC.n467 1.1255
R1632 VCC.n866 VCC.n403 1.1255
R1633 VCC.n1294 VCC.n1019 1.1255
R1634 VCC.n1418 VCC.n955 1.1255
R1635 VCC.n1981 VCC.n1513 1.1255
R1636 VCC.n1851 VCC.n1576 1.1255
R1637 VCC.n183 VCC.n182 1.1255
R1638 VCC.n334 VCC.n333 1.1255
R1639 VCC.n579 VCC.n573 1.00621
R1640 VCC.n567 VCC.n561 1.00621
R1641 VCC.n526 VCC.n525 1.00621
R1642 VCC.n699 VCC.n490 1.00621
R1643 VCC.n692 VCC.n691 1.00621
R1644 VCC.n757 VCC.n461 1.00621
R1645 VCC.n788 VCC.n787 1.00621
R1646 VCC.n911 VCC.n369 1.00621
R1647 VCC.n1131 VCC.n1125 1.00621
R1648 VCC.n1119 VCC.n1113 1.00621
R1649 VCC.n1078 VCC.n1077 1.00621
R1650 VCC.n1251 VCC.n1042 1.00621
R1651 VCC.n1244 VCC.n1243 1.00621
R1652 VCC.n1309 VCC.n1013 1.00621
R1653 VCC.n1340 VCC.n1339 1.00621
R1654 VCC.n1465 VCC.n923 1.00621
R1655 VCC.n1898 VCC.n1897 1.00621
R1656 VCC.n2022 VCC.n1478 1.00621
R1657 VCC.n1808 VCC.n1599 1.00621
R1658 VCC.n1801 VCC.n1800 1.00621
R1659 VCC.n1866 VCC.n1570 1.00621
R1660 VCC.n1689 VCC.n1683 1.00621
R1661 VCC.n1677 VCC.n1671 1.00621
R1662 VCC.n1636 VCC.n1635 1.00621
R1663 VCC.n34 VCC.n31 1.00621
R1664 VCC.n33 VCC.n32 1.00621
R1665 VCC.n200 VCC.n190 1.00621
R1666 VCC.n2 VCC.n1 1.00621
R1667 VCC.n280 VCC.n279 1.00621
R1668 VCC.n596 VCC.n546 0.9505
R1669 VCC.n635 VCC.n509 0.9505
R1670 VCC.n725 VCC.n473 0.9505
R1671 VCC.n763 VCC.n458 0.9505
R1672 VCC.n1148 VCC.n1098 0.9505
R1673 VCC.n1187 VCC.n1061 0.9505
R1674 VCC.n1277 VCC.n1025 0.9505
R1675 VCC.n1315 VCC.n1010 0.9505
R1676 VCC.n1834 VCC.n1582 0.9505
R1677 VCC.n1872 VCC.n1567 0.9505
R1678 VCC.n1706 VCC.n1656 0.9505
R1679 VCC.n1745 VCC.n1619 0.9505
R1680 VCC.n68 VCC.n67 0.9505
R1681 VCC.n193 VCC.n192 0.9505
R1682 VCC.n614 VCC.n613 0.914786
R1683 VCC.n629 VCC.n522 0.914786
R1684 VCC.n663 VCC.n505 0.914786
R1685 VCC.n662 VCC.n661 0.914786
R1686 VCC.n732 VCC.n731 0.914786
R1687 VCC.n750 VCC.n463 0.914786
R1688 VCC.n798 VCC.n444 0.914786
R1689 VCC.n797 VCC.n796 0.914786
R1690 VCC.n1166 VCC.n1165 0.914786
R1691 VCC.n1181 VCC.n1074 0.914786
R1692 VCC.n1215 VCC.n1057 0.914786
R1693 VCC.n1214 VCC.n1213 0.914786
R1694 VCC.n1284 VCC.n1283 0.914786
R1695 VCC.n1302 VCC.n1015 0.914786
R1696 VCC.n1350 VCC.n996 0.914786
R1697 VCC.n1349 VCC.n1348 0.914786
R1698 VCC.n1841 VCC.n1840 0.914786
R1699 VCC.n1859 VCC.n1572 0.914786
R1700 VCC.n1908 VCC.n1553 0.914786
R1701 VCC.n1907 VCC.n1906 0.914786
R1702 VCC.n1724 VCC.n1723 0.914786
R1703 VCC.n1739 VCC.n1632 0.914786
R1704 VCC.n1773 VCC.n1615 0.914786
R1705 VCC.n1772 VCC.n1771 0.914786
R1706 VCC.n75 VCC.n74 0.914786
R1707 VCC.n81 VCC.n79 0.914786
R1708 VCC.n22 VCC.n21 0.914786
R1709 VCC.n223 VCC.n222 0.914786
R1710 VCC.n589 VCC.n550 0.823357
R1711 VCC.n598 VCC.n543 0.823357
R1712 VCC.n615 VCC.n521 0.823357
R1713 VCC.n651 VCC.n510 0.823357
R1714 VCC.n707 VCC.n706 0.823357
R1715 VCC.n723 VCC.n476 0.823357
R1716 VCC.n753 VCC.n752 0.823357
R1717 VCC.n778 VCC.n450 0.823357
R1718 VCC.n1141 VCC.n1102 0.823357
R1719 VCC.n1150 VCC.n1095 0.823357
R1720 VCC.n1167 VCC.n1073 0.823357
R1721 VCC.n1203 VCC.n1062 0.823357
R1722 VCC.n1259 VCC.n1258 0.823357
R1723 VCC.n1275 VCC.n1028 0.823357
R1724 VCC.n1305 VCC.n1304 0.823357
R1725 VCC.n1330 VCC.n1002 0.823357
R1726 VCC.n1816 VCC.n1815 0.823357
R1727 VCC.n1832 VCC.n1585 0.823357
R1728 VCC.n1862 VCC.n1861 0.823357
R1729 VCC.n1887 VCC.n1559 0.823357
R1730 VCC.n1699 VCC.n1660 0.823357
R1731 VCC.n1708 VCC.n1653 0.823357
R1732 VCC.n1725 VCC.n1631 0.823357
R1733 VCC.n1761 VCC.n1620 0.823357
R1734 VCC.n55 VCC.n52 0.823357
R1735 VCC.n54 VCC.n53 0.823357
R1736 VCC.n186 VCC.n185 0.823357
R1737 VCC.n11 VCC.n10 0.823357
R1738 VCC.n550 VCC.n543 0.731929
R1739 VCC.n638 VCC.n510 0.731929
R1740 VCC.n653 VCC.n651 0.731929
R1741 VCC.n706 VCC.n476 0.731929
R1742 VCC.n765 VCC.n450 0.731929
R1743 VCC.n779 VCC.n778 0.731929
R1744 VCC.n1102 VCC.n1095 0.731929
R1745 VCC.n1190 VCC.n1062 0.731929
R1746 VCC.n1205 VCC.n1203 0.731929
R1747 VCC.n1258 VCC.n1028 0.731929
R1748 VCC.n1317 VCC.n1002 0.731929
R1749 VCC.n1331 VCC.n1330 0.731929
R1750 VCC.n1815 VCC.n1585 0.731929
R1751 VCC.n1874 VCC.n1559 0.731929
R1752 VCC.n1888 VCC.n1887 0.731929
R1753 VCC.n1660 VCC.n1653 0.731929
R1754 VCC.n1748 VCC.n1620 0.731929
R1755 VCC.n1763 VCC.n1761 0.731929
R1756 VCC.n55 VCC.n54 0.731929
R1757 VCC.n10 VCC.n9 0.731929
R1758 VCC.n18 VCC.n11 0.731929
R1759 VCC.n613 VCC.n535 0.6405
R1760 VCC.n663 VCC.n662 0.6405
R1761 VCC.n732 VCC.n730 0.6405
R1762 VCC.n798 VCC.n797 0.6405
R1763 VCC.n1165 VCC.n1087 0.6405
R1764 VCC.n1215 VCC.n1214 0.6405
R1765 VCC.n1284 VCC.n1282 0.6405
R1766 VCC.n1350 VCC.n1349 0.6405
R1767 VCC.n1841 VCC.n1839 0.6405
R1768 VCC.n1908 VCC.n1907 0.6405
R1769 VCC.n1723 VCC.n1645 0.6405
R1770 VCC.n1773 VCC.n1772 0.6405
R1771 VCC.n75 VCC.n73 0.6405
R1772 VCC.n222 VCC.n22 0.6405
R1773 VCC.n573 VCC.n561 0.549071
R1774 VCC.n525 VCC.n517 0.549071
R1775 VCC.n691 VCC.n490 0.549071
R1776 VCC.n758 VCC.n757 0.549071
R1777 VCC.n1125 VCC.n1113 0.549071
R1778 VCC.n1077 VCC.n1069 0.549071
R1779 VCC.n1243 VCC.n1042 0.549071
R1780 VCC.n1310 VCC.n1309 0.549071
R1781 VCC.n1800 VCC.n1599 0.549071
R1782 VCC.n1867 VCC.n1866 0.549071
R1783 VCC.n1683 VCC.n1671 0.549071
R1784 VCC.n1635 VCC.n1627 0.549071
R1785 VCC.n34 VCC.n33 0.549071
R1786 VCC.n200 VCC.n199 0.549071
R1787 VCC.n815 VCC 0.535293
R1788 VCC.n1367 VCC 0.535293
R1789 VCC.n1925 VCC 0.535293
R1790 VCC VCC.n169 0.535293
R1791 VCC.n915 VCC.n369 0.507747
R1792 VCC.n1469 VCC.n923 0.507747
R1793 VCC.n2023 VCC.n2022 0.507747
R1794 VCC.n285 VCC.n280 0.507747
R1795 VCC.n1898 VCC.n1540 0.465127
R1796 VCC.n788 VCC.n431 0.465115
R1797 VCC.n1340 VCC.n983 0.465115
R1798 VCC.n232 VCC.n2 0.465115
R1799 VCC.n615 VCC.n614 0.366214
R1800 VCC.n834 VCC.n420 0.366214
R1801 VCC.n897 VCC.n895 0.366214
R1802 VCC.n1167 VCC.n1166 0.366214
R1803 VCC.n1386 VCC.n972 0.366214
R1804 VCC.n1449 VCC.n1447 0.366214
R1805 VCC.n1944 VCC.n1943 0.366214
R1806 VCC.n2015 VCC.n2014 0.366214
R1807 VCC.n1725 VCC.n1724 0.366214
R1808 VCC.n249 VCC.n248 0.366214
R1809 VCC.n303 VCC.n296 0.366214
R1810 VCC VCC.n919 0.338784
R1811 VCC VCC.n918 0.300964
R1812 VCC VCC.n1472 0.300964
R1813 VCC VCC.n2026 0.300964
R1814 VCC VCC.n365 0.300964
R1815 VCC.n557 VCC 0.294921
R1816 VCC.n1109 VCC 0.294921
R1817 VCC.n1667 VCC 0.294921
R1818 VCC.n102 VCC 0.294921
R1819 VCC.n681 VCC 0.287536
R1820 VCC.n1233 VCC 0.287536
R1821 VCC.n1791 VCC 0.287536
R1822 VCC.n590 VCC.n549 0.274786
R1823 VCC.n652 VCC.n507 0.274786
R1824 VCC.n705 VCC.n484 0.274786
R1825 VCC.n731 VCC.n463 0.274786
R1826 VCC.n753 VCC.n461 0.274786
R1827 VCC.n781 VCC.n780 0.274786
R1828 VCC.n1142 VCC.n1101 0.274786
R1829 VCC.n1204 VCC.n1059 0.274786
R1830 VCC.n1257 VCC.n1036 0.274786
R1831 VCC.n1283 VCC.n1015 0.274786
R1832 VCC.n1305 VCC.n1013 0.274786
R1833 VCC.n1333 VCC.n1332 0.274786
R1834 VCC.n1814 VCC.n1593 0.274786
R1835 VCC.n1840 VCC.n1572 0.274786
R1836 VCC.n1862 VCC.n1570 0.274786
R1837 VCC.n1890 VCC.n1889 0.274786
R1838 VCC.n1700 VCC.n1659 0.274786
R1839 VCC.n1762 VCC.n1617 0.274786
R1840 VCC.n45 VCC.n44 0.274786
R1841 VCC.n20 VCC.n19 0.274786
R1842 VCC VCC.n679 0.213679
R1843 VCC VCC.n1231 0.213679
R1844 VCC VCC.n1789 0.213679
R1845 VCC.n526 VCC.n522 0.183357
R1846 VCC.n856 VCC.n409 0.183357
R1847 VCC.n857 VCC.n856 0.183357
R1848 VCC.n889 VCC.n390 0.183357
R1849 VCC.n889 VCC.n391 0.183357
R1850 VCC.n1078 VCC.n1074 0.183357
R1851 VCC.n1408 VCC.n961 0.183357
R1852 VCC.n1409 VCC.n1408 0.183357
R1853 VCC.n1441 VCC.n942 0.183357
R1854 VCC.n1441 VCC.n943 0.183357
R1855 VCC.n1959 VCC.n1953 0.183357
R1856 VCC.n1953 VCC.n1526 0.183357
R1857 VCC.n1989 VCC.n1501 0.183357
R1858 VCC.n1989 VCC.n1507 0.183357
R1859 VCC.n1636 VCC.n1632 0.183357
R1860 VCC.n268 VCC.n267 0.183357
R1861 VCC.n267 VCC.n260 0.183357
R1862 VCC.n323 VCC.n316 0.183357
R1863 VCC.n325 VCC.n323 0.183357
R1864 VCC VCC.n814 0.114307
R1865 VCC VCC.n1366 0.114307
R1866 VCC VCC.n1924 0.114307
R1867 VCC.n170 VCC 0.114307
R1868 VCC.n597 VCC.n544 0.0919286
R1869 VCC.n637 VCC.n636 0.0919286
R1870 VCC.n724 VCC.n472 0.0919286
R1871 VCC.n764 VCC.n457 0.0919286
R1872 VCC.n897 VCC.n896 0.0919286
R1873 VCC.n910 VCC.n373 0.0919286
R1874 VCC.n1149 VCC.n1096 0.0919286
R1875 VCC.n1189 VCC.n1188 0.0919286
R1876 VCC.n1276 VCC.n1024 0.0919286
R1877 VCC.n1316 VCC.n1009 0.0919286
R1878 VCC.n1449 VCC.n1448 0.0919286
R1879 VCC.n1464 VCC.n927 0.0919286
R1880 VCC.n2014 VCC.n1483 0.0919286
R1881 VCC.n1490 VCC.n1489 0.0919286
R1882 VCC.n1833 VCC.n1581 0.0919286
R1883 VCC.n1873 VCC.n1566 0.0919286
R1884 VCC.n1707 VCC.n1654 0.0919286
R1885 VCC.n1747 VCC.n1746 0.0919286
R1886 VCC.n66 VCC.n65 0.0919286
R1887 VCC.n8 VCC.n7 0.0919286
R1888 VCC.n306 VCC.n303 0.0919286
R1889 VCC.n305 VCC.n304 0.0919286
R1890 VCC.n1473 VCC 0.0247197
R1891 VCC.n919 VCC 0.0246714
R1892 VCC.n2027 VCC 0.0246714
R1893 VCC.n584 VCC.n583 0.024
R1894 VCC.n674 VCC.n673 0.024
R1895 VCC.n683 VCC.n480 0.024
R1896 VCC.n809 VCC.n808 0.024
R1897 VCC.n827 VCC.n826 0.024
R1898 VCC.n903 VCC.n902 0.024
R1899 VCC.n1136 VCC.n1135 0.024
R1900 VCC.n1226 VCC.n1225 0.024
R1901 VCC.n1235 VCC.n1032 0.024
R1902 VCC.n1361 VCC.n1360 0.024
R1903 VCC.n1379 VCC.n1378 0.024
R1904 VCC.n1455 VCC.n1454 0.024
R1905 VCC.n1694 VCC.n1693 0.024
R1906 VCC.n1784 VCC.n1783 0.024
R1907 VCC.n1793 VCC.n1589 0.024
R1908 VCC.n1919 VCC.n1918 0.024
R1909 VCC.n1938 VCC.n1937 0.024
R1910 VCC.n2002 VCC.n2001 0.024
R1911 VCC.n105 VCC.n104 0.024
R1912 VCC.n173 VCC.n172 0.024
R1913 VCC.n162 VCC.n161 0.024
R1914 VCC.n356 VCC.n355 0.024
R1915 VCC.n413 VCC.n404 0.0228214
R1916 VCC.n875 VCC.n874 0.0228214
R1917 VCC.n883 VCC.n382 0.0228214
R1918 VCC.n965 VCC.n956 0.0228214
R1919 VCC.n1427 VCC.n1426 0.0228214
R1920 VCC.n1435 VCC.n934 0.0228214
R1921 VCC.n1971 VCC.n1970 0.0228214
R1922 VCC.n1514 VCC.n1499 0.0228214
R1923 VCC.n1998 VCC.n1494 0.0228214
R1924 VCC.n274 VCC.n273 0.0228214
R1925 VCC.n331 VCC.n330 0.0228214
R1926 VCC.n312 VCC.n311 0.0228214
R1927 VCC.n919 VCC 0.0199714
R1928 VCC.n2027 VCC 0.0199714
R1929 VCC.n619 VCC.n523 0.0174643
R1930 VCC.n618 VCC.n529 0.0174643
R1931 VCC.n742 VCC.n465 0.0174643
R1932 VCC.n743 VCC.n742 0.0174643
R1933 VCC.n747 VCC.n467 0.0174643
R1934 VCC.n744 VCC.n467 0.0174643
R1935 VCC.n867 VCC.n866 0.0174643
R1936 VCC.n866 VCC.n398 0.0174643
R1937 VCC.n868 VCC.n403 0.0174643
R1938 VCC.n403 VCC.n399 0.0174643
R1939 VCC.n1171 VCC.n1075 0.0174643
R1940 VCC.n1170 VCC.n1081 0.0174643
R1941 VCC.n1294 VCC.n1017 0.0174643
R1942 VCC.n1295 VCC.n1294 0.0174643
R1943 VCC.n1299 VCC.n1019 0.0174643
R1944 VCC.n1296 VCC.n1019 0.0174643
R1945 VCC.n1419 VCC.n1418 0.0174643
R1946 VCC.n1418 VCC.n950 0.0174643
R1947 VCC.n1420 VCC.n955 0.0174643
R1948 VCC.n955 VCC.n951 0.0174643
R1949 VCC.n1981 VCC.n1512 0.0174643
R1950 VCC.n1981 VCC.n1980 0.0174643
R1951 VCC.n1973 VCC.n1513 0.0174643
R1952 VCC.n1979 VCC.n1513 0.0174643
R1953 VCC.n1851 VCC.n1574 0.0174643
R1954 VCC.n1852 VCC.n1851 0.0174643
R1955 VCC.n1856 VCC.n1576 0.0174643
R1956 VCC.n1853 VCC.n1576 0.0174643
R1957 VCC.n1729 VCC.n1633 0.0174643
R1958 VCC.n1728 VCC.n1639 0.0174643
R1959 VCC.n183 VCC.n83 0.0174643
R1960 VCC.n184 VCC.n183 0.0174643
R1961 VCC.n182 VCC.n115 0.0174643
R1962 VCC.n182 VCC.n181 0.0174643
R1963 VCC.n333 VCC.n275 0.0174643
R1964 VCC.n333 VCC.n332 0.0174643
R1965 VCC.n335 VCC.n334 0.0174643
R1966 VCC.n604 VCC.n599 0.0165714
R1967 VCC.n621 VCC.n620 0.0165714
R1968 VCC.n570 VCC.n563 0.0165714
R1969 VCC.n606 VCC.n605 0.0165714
R1970 VCC.n622 VCC.n533 0.0165714
R1971 VCC.n648 VCC.n512 0.0165714
R1972 VCC.n667 VCC.n666 0.0165714
R1973 VCC.n767 VCC.n766 0.0165714
R1974 VCC.n695 VCC.n687 0.0165714
R1975 VCC.n720 VCC.n714 0.0165714
R1976 VCC.n775 VCC.n452 0.0165714
R1977 VCC.n802 VCC.n801 0.0165714
R1978 VCC.n820 VCC.n426 0.0165714
R1979 VCC.n880 VCC.n395 0.0165714
R1980 VCC.n907 VCC.n376 0.0165714
R1981 VCC.n1156 VCC.n1151 0.0165714
R1982 VCC.n1173 VCC.n1172 0.0165714
R1983 VCC.n1122 VCC.n1115 0.0165714
R1984 VCC.n1158 VCC.n1157 0.0165714
R1985 VCC.n1174 VCC.n1085 0.0165714
R1986 VCC.n1200 VCC.n1064 0.0165714
R1987 VCC.n1219 VCC.n1218 0.0165714
R1988 VCC.n1319 VCC.n1318 0.0165714
R1989 VCC.n1247 VCC.n1239 0.0165714
R1990 VCC.n1272 VCC.n1266 0.0165714
R1991 VCC.n1327 VCC.n1004 0.0165714
R1992 VCC.n1354 VCC.n1353 0.0165714
R1993 VCC.n1372 VCC.n978 0.0165714
R1994 VCC.n1432 VCC.n947 0.0165714
R1995 VCC.n1461 VCC.n930 0.0165714
R1996 VCC.n1931 VCC.n1930 0.0165714
R1997 VCC.n1997 VCC.n1996 0.0165714
R1998 VCC.n2010 VCC.n2009 0.0165714
R1999 VCC.n1876 VCC.n1875 0.0165714
R2000 VCC.n1804 VCC.n1795 0.0165714
R2001 VCC.n1829 VCC.n1823 0.0165714
R2002 VCC.n1884 VCC.n1561 0.0165714
R2003 VCC.n1912 VCC.n1911 0.0165714
R2004 VCC.n1714 VCC.n1709 0.0165714
R2005 VCC.n1731 VCC.n1730 0.0165714
R2006 VCC.n1680 VCC.n1673 0.0165714
R2007 VCC.n1716 VCC.n1715 0.0165714
R2008 VCC.n1732 VCC.n1643 0.0165714
R2009 VCC.n1758 VCC.n1622 0.0165714
R2010 VCC.n1777 VCC.n1776 0.0165714
R2011 VCC.n207 VCC.n206 0.0165714
R2012 VCC.n90 VCC.n89 0.0165714
R2013 VCC.n97 VCC.n96 0.0165714
R2014 VCC.n129 VCC.n128 0.0165714
R2015 VCC.n122 VCC.n121 0.0165714
R2016 VCC.n153 VCC.n152 0.0165714
R2017 VCC.n349 VCC.n348 0.0165714
R2018 VCC.n358 VCC.n357 0.0165714
R2019 VCC.n640 VCC.n639 0.0156786
R2020 VCC.n606 VCC.n540 0.0156786
R2021 VCC.n722 VCC.n721 0.0156786
R2022 VCC.n776 VCC.n775 0.0156786
R2023 VCC.n846 VCC.n416 0.0156786
R2024 VCC.n1192 VCC.n1191 0.0156786
R2025 VCC.n1158 VCC.n1092 0.0156786
R2026 VCC.n1274 VCC.n1273 0.0156786
R2027 VCC.n1328 VCC.n1327 0.0156786
R2028 VCC.n1398 VCC.n968 0.0156786
R2029 VCC.n1964 VCC.n1521 0.0156786
R2030 VCC.n1831 VCC.n1830 0.0156786
R2031 VCC.n1885 VCC.n1884 0.0156786
R2032 VCC.n1750 VCC.n1749 0.0156786
R2033 VCC.n1716 VCC.n1650 0.0156786
R2034 VCC.n59 VCC.n58 0.0156786
R2035 VCC.n128 VCC.n127 0.0156786
R2036 VCC.n158 VCC.n157 0.0156786
R2037 VCC.n608 VCC.n607 0.0152714
R2038 VCC.n647 VCC.n646 0.0152714
R2039 VCC.n713 VCC.n468 0.0152714
R2040 VCC.n774 VCC.n773 0.0152714
R2041 VCC.n851 VCC.n847 0.0152714
R2042 VCC.n879 VCC.n878 0.0152714
R2043 VCC.n1160 VCC.n1159 0.0152714
R2044 VCC.n1199 VCC.n1198 0.0152714
R2045 VCC.n1265 VCC.n1020 0.0152714
R2046 VCC.n1326 VCC.n1325 0.0152714
R2047 VCC.n1403 VCC.n1399 0.0152714
R2048 VCC.n1431 VCC.n1430 0.0152714
R2049 VCC.n1718 VCC.n1717 0.0152714
R2050 VCC.n1757 VCC.n1756 0.0152714
R2051 VCC.n1822 VCC.n1577 0.0152714
R2052 VCC.n1883 VCC.n1882 0.0152714
R2053 VCC.n1966 VCC.n1965 0.0152714
R2054 VCC.n1995 VCC.n1994 0.0152714
R2055 VCC.n108 VCC.n107 0.0152714
R2056 VCC.n176 VCC.n175 0.0152714
R2057 VCC.n151 VCC.n150 0.0152714
R2058 VCC.n344 VCC.n343 0.0152714
R2059 VCC.n649 VCC.n648 0.0147857
R2060 VCC.n714 VCC.n479 0.0147857
R2061 VCC.n828 VCC.n418 0.0147857
R2062 VCC.n1201 VCC.n1200 0.0147857
R2063 VCC.n1266 VCC.n1031 0.0147857
R2064 VCC.n1380 VCC.n970 0.0147857
R2065 VCC.n1534 VCC.n1523 0.0147857
R2066 VCC.n1823 VCC.n1588 0.0147857
R2067 VCC.n1759 VCC.n1758 0.0147857
R2068 VCC.n96 VCC.n95 0.0147857
R2069 VCC.n254 VCC.n253 0.0147857
R2070 VCC.n624 VCC.n623 0.0132571
R2071 VCC.n746 VCC.n745 0.0132571
R2072 VCC.n870 VCC.n869 0.0132571
R2073 VCC.n1176 VCC.n1175 0.0132571
R2074 VCC.n1298 VCC.n1297 0.0132571
R2075 VCC.n1422 VCC.n1421 0.0132571
R2076 VCC.n1734 VCC.n1733 0.0132571
R2077 VCC.n1855 VCC.n1854 0.0132571
R2078 VCC.n1978 VCC.n1974 0.0132571
R2079 VCC.n137 VCC.n136 0.0132571
R2080 VCC.n568 VCC.n566 0.013
R2081 VCC.n442 VCC.n440 0.013
R2082 VCC.n908 VCC.n375 0.013
R2083 VCC.n916 VCC.n368 0.013
R2084 VCC.n907 VCC.n906 0.013
R2085 VCC.n1120 VCC.n1118 0.013
R2086 VCC.n994 VCC.n992 0.013
R2087 VCC.n1462 VCC.n929 0.013
R2088 VCC.n1470 VCC.n922 0.013
R2089 VCC.n1461 VCC.n1460 0.013
R2090 VCC.n2008 VCC.n2007 0.013
R2091 VCC.n2024 VCC.n1476 0.013
R2092 VCC.n2009 VCC.n1487 0.013
R2093 VCC.n1551 VCC.n1549 0.013
R2094 VCC.n1678 VCC.n1676 0.013
R2095 VCC.n215 VCC.n214 0.013
R2096 VCC.n291 VCC.n290 0.013
R2097 VCC.n287 VCC.n286 0.013
R2098 VCC.n359 VCC.n358 0.013
R2099 VCC.n503 VCC.n501 0.0121071
R2100 VCC.n571 VCC.n570 0.0121071
R2101 VCC.n693 VCC.n690 0.0121071
R2102 VCC.n812 VCC.n811 0.0121071
R2103 VCC.n801 VCC.n441 0.0121071
R2104 VCC.n824 VCC.n817 0.0121071
R2105 VCC.n822 VCC.n819 0.0121071
R2106 VCC.n821 VCC.n820 0.0121071
R2107 VCC.n384 VCC.n381 0.0121071
R2108 VCC.n1055 VCC.n1053 0.0121071
R2109 VCC.n1123 VCC.n1122 0.0121071
R2110 VCC.n1245 VCC.n1242 0.0121071
R2111 VCC.n1364 VCC.n1363 0.0121071
R2112 VCC.n1353 VCC.n993 0.0121071
R2113 VCC.n1376 VCC.n1369 0.0121071
R2114 VCC.n1374 VCC.n1371 0.0121071
R2115 VCC.n1373 VCC.n1372 0.0121071
R2116 VCC.n936 VCC.n933 0.0121071
R2117 VCC.n1935 VCC.n1927 0.0121071
R2118 VCC.n1933 VCC.n1929 0.0121071
R2119 VCC.n1932 VCC.n1931 0.0121071
R2120 VCC.n2011 VCC.n1486 0.0121071
R2121 VCC.n1802 VCC.n1799 0.0121071
R2122 VCC.n1922 VCC.n1921 0.0121071
R2123 VCC.n1911 VCC.n1550 0.0121071
R2124 VCC.n1613 VCC.n1611 0.0121071
R2125 VCC.n1681 VCC.n1680 0.0121071
R2126 VCC.n39 VCC.n38 0.0121071
R2127 VCC.n219 VCC.n218 0.0121071
R2128 VCC.n121 VCC.n120 0.0121071
R2129 VCC.n234 VCC.n233 0.0121071
R2130 VCC.n237 VCC.n236 0.0121071
R2131 VCC.n351 VCC.n350 0.0121071
R2132 VCC.n565 VCC.n551 0.0112143
R2133 VCC.n669 VCC.n501 0.0112143
R2134 VCC.n677 VCC.n676 0.0112143
R2135 VCC.n564 VCC.n552 0.0112143
R2136 VCC.n668 VCC.n667 0.0112143
R2137 VCC.n666 VCC.n502 0.0112143
R2138 VCC.n690 VCC.n689 0.0112143
R2139 VCC.n805 VCC.n804 0.0112143
R2140 VCC.n696 VCC.n695 0.0112143
R2141 VCC.n688 VCC.n687 0.0112143
R2142 VCC.n803 VCC.n438 0.0112143
R2143 VCC.n819 VCC.n818 0.0112143
R2144 VCC.n833 VCC.n425 0.0112143
R2145 VCC.n899 VCC.n898 0.0112143
R2146 VCC.n832 VCC.n831 0.0112143
R2147 VCC.n1117 VCC.n1103 0.0112143
R2148 VCC.n1221 VCC.n1053 0.0112143
R2149 VCC.n1229 VCC.n1228 0.0112143
R2150 VCC.n1116 VCC.n1104 0.0112143
R2151 VCC.n1220 VCC.n1219 0.0112143
R2152 VCC.n1218 VCC.n1054 0.0112143
R2153 VCC.n1242 VCC.n1241 0.0112143
R2154 VCC.n1357 VCC.n1356 0.0112143
R2155 VCC.n1248 VCC.n1247 0.0112143
R2156 VCC.n1240 VCC.n1239 0.0112143
R2157 VCC.n1355 VCC.n990 0.0112143
R2158 VCC.n1371 VCC.n1370 0.0112143
R2159 VCC.n1385 VCC.n977 0.0112143
R2160 VCC.n1451 VCC.n1450 0.0112143
R2161 VCC.n1384 VCC.n1383 0.0112143
R2162 VCC.n1929 VCC.n1928 0.0112143
R2163 VCC.n1942 VCC.n1941 0.0112143
R2164 VCC.n2013 VCC.n1484 0.0112143
R2165 VCC.n1940 VCC.n1533 0.0112143
R2166 VCC.n1799 VCC.n1798 0.0112143
R2167 VCC.n1915 VCC.n1914 0.0112143
R2168 VCC.n1805 VCC.n1804 0.0112143
R2169 VCC.n1797 VCC.n1795 0.0112143
R2170 VCC.n1913 VCC.n1547 0.0112143
R2171 VCC.n1675 VCC.n1661 0.0112143
R2172 VCC.n1779 VCC.n1611 0.0112143
R2173 VCC.n1787 VCC.n1786 0.0112143
R2174 VCC.n1674 VCC.n1662 0.0112143
R2175 VCC.n1778 VCC.n1777 0.0112143
R2176 VCC.n1776 VCC.n1612 0.0112143
R2177 VCC.n40 VCC.n39 0.0112143
R2178 VCC.n213 VCC.n212 0.0112143
R2179 VCC.n89 VCC.n88 0.0112143
R2180 VCC.n91 VCC.n90 0.0112143
R2181 VCC.n124 VCC.n123 0.0112143
R2182 VCC.n238 VCC.n237 0.0112143
R2183 VCC.n251 VCC.n250 0.0112143
R2184 VCC.n309 VCC.n308 0.0112143
R2185 VCC.n155 VCC.n154 0.0112143
R2186 VCC.n566 VCC.n565 0.0103214
R2187 VCC.n601 VCC.n536 0.0103214
R2188 VCC.n527 VCC.n524 0.0103214
R2189 VCC.n644 VCC.n643 0.0103214
R2190 VCC.n670 VCC.n669 0.0103214
R2191 VCC.n564 VCC.n563 0.0103214
R2192 VCC.n600 VCC.n537 0.0103214
R2193 VCC.n645 VCC.n515 0.0103214
R2194 VCC.n668 VCC.n499 0.0103214
R2195 VCC.n502 VCC.n496 0.0103214
R2196 VCC.n698 VCC.n697 0.0103214
R2197 VCC.n689 VCC.n482 0.0103214
R2198 VCC.n717 VCC.n716 0.0103214
R2199 VCC.n756 VCC.n755 0.0103214
R2200 VCC.n771 VCC.n770 0.0103214
R2201 VCC.n804 VCC.n440 0.0103214
R2202 VCC.n696 VCC.n685 0.0103214
R2203 VCC.n688 VCC.n481 0.0103214
R2204 VCC.n715 VCC.n469 0.0103214
R2205 VCC.n772 VCC.n455 0.0103214
R2206 VCC.n803 VCC.n802 0.0103214
R2207 VCC.n833 VCC.n424 0.0103214
R2208 VCC.n829 VCC.n828 0.0103214
R2209 VCC.n854 VCC.n411 0.0103214
R2210 VCC.n876 VCC.n392 0.0103214
R2211 VCC.n909 VCC.n908 0.0103214
R2212 VCC.n832 VCC.n426 0.0103214
R2213 VCC.n853 VCC.n852 0.0103214
R2214 VCC.n848 VCC.n402 0.0103214
R2215 VCC.n877 VCC.n394 0.0103214
R2216 VCC.n885 VCC.n884 0.0103214
R2217 VCC.n1118 VCC.n1117 0.0103214
R2218 VCC.n1153 VCC.n1088 0.0103214
R2219 VCC.n1079 VCC.n1076 0.0103214
R2220 VCC.n1196 VCC.n1195 0.0103214
R2221 VCC.n1222 VCC.n1221 0.0103214
R2222 VCC.n1116 VCC.n1115 0.0103214
R2223 VCC.n1152 VCC.n1089 0.0103214
R2224 VCC.n1197 VCC.n1067 0.0103214
R2225 VCC.n1220 VCC.n1051 0.0103214
R2226 VCC.n1054 VCC.n1048 0.0103214
R2227 VCC.n1250 VCC.n1249 0.0103214
R2228 VCC.n1241 VCC.n1034 0.0103214
R2229 VCC.n1269 VCC.n1268 0.0103214
R2230 VCC.n1308 VCC.n1307 0.0103214
R2231 VCC.n1323 VCC.n1322 0.0103214
R2232 VCC.n1356 VCC.n992 0.0103214
R2233 VCC.n1248 VCC.n1237 0.0103214
R2234 VCC.n1240 VCC.n1033 0.0103214
R2235 VCC.n1267 VCC.n1021 0.0103214
R2236 VCC.n1324 VCC.n1007 0.0103214
R2237 VCC.n1355 VCC.n1354 0.0103214
R2238 VCC.n1385 VCC.n976 0.0103214
R2239 VCC.n1381 VCC.n1380 0.0103214
R2240 VCC.n1406 VCC.n963 0.0103214
R2241 VCC.n1428 VCC.n944 0.0103214
R2242 VCC.n1463 VCC.n1462 0.0103214
R2243 VCC.n1384 VCC.n978 0.0103214
R2244 VCC.n1405 VCC.n1404 0.0103214
R2245 VCC.n1400 VCC.n954 0.0103214
R2246 VCC.n1429 VCC.n946 0.0103214
R2247 VCC.n1437 VCC.n1436 0.0103214
R2248 VCC.n1942 VCC.n1532 0.0103214
R2249 VCC.n1535 VCC.n1534 0.0103214
R2250 VCC.n1955 VCC.n1518 0.0103214
R2251 VCC.n1992 VCC.n1991 0.0103214
R2252 VCC.n2008 VCC.n1491 0.0103214
R2253 VCC.n1930 VCC.n1533 0.0103214
R2254 VCC.n1956 VCC.n1519 0.0103214
R2255 VCC.n1972 VCC.n1517 0.0103214
R2256 VCC.n1993 VCC.n1498 0.0103214
R2257 VCC.n1503 VCC.n1495 0.0103214
R2258 VCC.n1807 VCC.n1601 0.0103214
R2259 VCC.n1798 VCC.n1591 0.0103214
R2260 VCC.n1826 VCC.n1825 0.0103214
R2261 VCC.n1865 VCC.n1864 0.0103214
R2262 VCC.n1880 VCC.n1879 0.0103214
R2263 VCC.n1914 VCC.n1549 0.0103214
R2264 VCC.n1806 VCC.n1805 0.0103214
R2265 VCC.n1797 VCC.n1590 0.0103214
R2266 VCC.n1824 VCC.n1578 0.0103214
R2267 VCC.n1881 VCC.n1564 0.0103214
R2268 VCC.n1913 VCC.n1912 0.0103214
R2269 VCC.n1676 VCC.n1675 0.0103214
R2270 VCC.n1711 VCC.n1646 0.0103214
R2271 VCC.n1637 VCC.n1634 0.0103214
R2272 VCC.n1754 VCC.n1753 0.0103214
R2273 VCC.n1780 VCC.n1779 0.0103214
R2274 VCC.n1674 VCC.n1673 0.0103214
R2275 VCC.n1710 VCC.n1647 0.0103214
R2276 VCC.n1755 VCC.n1625 0.0103214
R2277 VCC.n1778 VCC.n1609 0.0103214
R2278 VCC.n1612 VCC.n1606 0.0103214
R2279 VCC.n35 VCC.n24 0.0103214
R2280 VCC.n41 VCC.n40 0.0103214
R2281 VCC.n63 VCC.n62 0.0103214
R2282 VCC.n201 VCC.n189 0.0103214
R2283 VCC.n204 VCC.n203 0.0103214
R2284 VCC.n214 VCC.n213 0.0103214
R2285 VCC.n88 VCC.n87 0.0103214
R2286 VCC.n92 VCC.n91 0.0103214
R2287 VCC.n100 VCC.n99 0.0103214
R2288 VCC.n132 VCC.n131 0.0103214
R2289 VCC.n123 VCC.n122 0.0103214
R2290 VCC.n250 VCC.n239 0.0103214
R2291 VCC.n253 VCC.n252 0.0103214
R2292 VCC.n272 VCC.n271 0.0103214
R2293 VCC.n329 VCC.n328 0.0103214
R2294 VCC.n292 VCC.n291 0.0103214
R2295 VCC.n154 VCC.n153 0.0103214
R2296 VCC.n143 VCC.n142 0.0103214
R2297 VCC.n147 VCC.n146 0.0103214
R2298 VCC.n339 VCC.n338 0.0103214
R2299 VCC.n347 VCC.n346 0.0103214
R2300 VCC.n572 VCC.n559 0.00942857
R2301 VCC.n612 VCC.n534 0.00942857
R2302 VCC.n628 VCC.n528 0.00942857
R2303 VCC.n660 VCC.n504 0.00942857
R2304 VCC.n571 VCC.n556 0.00942857
R2305 VCC.n627 VCC.n626 0.00942857
R2306 VCC.n733 VCC.n471 0.00942857
R2307 VCC.n749 VCC.n464 0.00942857
R2308 VCC.n443 VCC.n434 0.00942857
R2309 VCC.n748 VCC.n466 0.00942857
R2310 VCC.n441 VCC.n435 0.00942857
R2311 VCC.n823 VCC.n822 0.00942857
R2312 VCC.n900 VCC.n382 0.00942857
R2313 VCC.n385 VCC.n383 0.00942857
R2314 VCC.n821 VCC.n430 0.00942857
R2315 VCC.n845 VCC.n417 0.00942857
R2316 VCC.n873 VCC.n872 0.00942857
R2317 VCC.n384 VCC.n376 0.00942857
R2318 VCC.n1124 VCC.n1111 0.00942857
R2319 VCC.n1164 VCC.n1086 0.00942857
R2320 VCC.n1180 VCC.n1080 0.00942857
R2321 VCC.n1212 VCC.n1056 0.00942857
R2322 VCC.n1123 VCC.n1108 0.00942857
R2323 VCC.n1179 VCC.n1178 0.00942857
R2324 VCC.n1285 VCC.n1023 0.00942857
R2325 VCC.n1301 VCC.n1016 0.00942857
R2326 VCC.n995 VCC.n986 0.00942857
R2327 VCC.n1300 VCC.n1018 0.00942857
R2328 VCC.n993 VCC.n987 0.00942857
R2329 VCC.n1375 VCC.n1374 0.00942857
R2330 VCC.n1452 VCC.n934 0.00942857
R2331 VCC.n937 VCC.n935 0.00942857
R2332 VCC.n1373 VCC.n982 0.00942857
R2333 VCC.n1397 VCC.n969 0.00942857
R2334 VCC.n1425 VCC.n1424 0.00942857
R2335 VCC.n936 VCC.n930 0.00942857
R2336 VCC.n1934 VCC.n1933 0.00942857
R2337 VCC.n1999 VCC.n1998 0.00942857
R2338 VCC.n2012 VCC.n1485 0.00942857
R2339 VCC.n1932 VCC.n1539 0.00942857
R2340 VCC.n1963 VCC.n1522 0.00942857
R2341 VCC.n1976 VCC.n1515 0.00942857
R2342 VCC.n2011 VCC.n2010 0.00942857
R2343 VCC.n1842 VCC.n1580 0.00942857
R2344 VCC.n1858 VCC.n1573 0.00942857
R2345 VCC.n1552 VCC.n1543 0.00942857
R2346 VCC.n1857 VCC.n1575 0.00942857
R2347 VCC.n1550 VCC.n1544 0.00942857
R2348 VCC.n1682 VCC.n1669 0.00942857
R2349 VCC.n1722 VCC.n1644 0.00942857
R2350 VCC.n1738 VCC.n1638 0.00942857
R2351 VCC.n1770 VCC.n1614 0.00942857
R2352 VCC.n1681 VCC.n1666 0.00942857
R2353 VCC.n1737 VCC.n1736 0.00942857
R2354 VCC.n77 VCC.n76 0.00942857
R2355 VCC.n82 VCC.n78 0.00942857
R2356 VCC.n221 VCC.n220 0.00942857
R2357 VCC.n114 VCC.n113 0.00942857
R2358 VCC.n120 VCC.n119 0.00942857
R2359 VCC.n236 VCC.n235 0.00942857
R2360 VCC.n311 VCC.n310 0.00942857
R2361 VCC.n307 VCC.n294 0.00942857
R2362 VCC.n165 VCC.n164 0.00942857
R2363 VCC.n140 VCC.n139 0.00942857
R2364 VCC.n337 VCC.n336 0.00942857
R2365 VCC.n588 VCC.n587 0.00853571
R2366 VCC.n599 VCC.n542 0.00853571
R2367 VCC.n617 VCC.n616 0.00853571
R2368 VCC.n650 VCC.n511 0.00853571
R2369 VCC.n538 VCC.n532 0.00853571
R2370 VCC.n708 VCC.n483 0.00853571
R2371 VCC.n722 VCC.n477 0.00853571
R2372 VCC.n754 VCC.n462 0.00853571
R2373 VCC.n777 VCC.n451 0.00853571
R2374 VCC.n741 VCC.n740 0.00853571
R2375 VCC.n844 VCC.n418 0.00853571
R2376 VCC.n906 VCC.n905 0.00853571
R2377 VCC.n917 VCC.n367 0.00853571
R2378 VCC.n1140 VCC.n1139 0.00853571
R2379 VCC.n1151 VCC.n1094 0.00853571
R2380 VCC.n1169 VCC.n1168 0.00853571
R2381 VCC.n1202 VCC.n1063 0.00853571
R2382 VCC.n1090 VCC.n1084 0.00853571
R2383 VCC.n1260 VCC.n1035 0.00853571
R2384 VCC.n1274 VCC.n1029 0.00853571
R2385 VCC.n1306 VCC.n1014 0.00853571
R2386 VCC.n1329 VCC.n1003 0.00853571
R2387 VCC.n1293 VCC.n1292 0.00853571
R2388 VCC.n1396 VCC.n970 0.00853571
R2389 VCC.n1460 VCC.n1459 0.00853571
R2390 VCC.n1471 VCC.n921 0.00853571
R2391 VCC.n1962 VCC.n1523 0.00853571
R2392 VCC.n2004 VCC.n1487 0.00853571
R2393 VCC.n2025 VCC.n1475 0.00853571
R2394 VCC.n1817 VCC.n1592 0.00853571
R2395 VCC.n1831 VCC.n1586 0.00853571
R2396 VCC.n1863 VCC.n1571 0.00853571
R2397 VCC.n1886 VCC.n1560 0.00853571
R2398 VCC.n1850 VCC.n1849 0.00853571
R2399 VCC.n1698 VCC.n1697 0.00853571
R2400 VCC.n1709 VCC.n1652 0.00853571
R2401 VCC.n1727 VCC.n1726 0.00853571
R2402 VCC.n1760 VCC.n1621 0.00853571
R2403 VCC.n1648 VCC.n1642 0.00853571
R2404 VCC.n56 VCC.n43 0.00853571
R2405 VCC.n58 VCC.n57 0.00853571
R2406 VCC.n188 VCC.n187 0.00853571
R2407 VCC.n209 VCC.n208 0.00853571
R2408 VCC.n180 VCC.n179 0.00853571
R2409 VCC.n255 VCC.n254 0.00853571
R2410 VCC.n360 VCC.n359 0.00853571
R2411 VCC.n363 VCC.n362 0.00853571
R2412 VCC.n557 VCC.n554 0.00822143
R2413 VCC.n607 VCC.n539 0.00822143
R2414 VCC.n647 VCC.n497 0.00822143
R2415 VCC.n679 VCC.n493 0.00822143
R2416 VCC.n682 VCC.n681 0.00822143
R2417 VCC.n713 VCC.n712 0.00822143
R2418 VCC.n774 VCC.n436 0.00822143
R2419 VCC.n814 VCC.n432 0.00822143
R2420 VCC.n815 VCC.n428 0.00822143
R2421 VCC.n847 VCC.n415 0.00822143
R2422 VCC.n879 VCC.n379 0.00822143
R2423 VCC.n918 VCC.n366 0.00822143
R2424 VCC.n1109 VCC.n1106 0.00822143
R2425 VCC.n1159 VCC.n1091 0.00822143
R2426 VCC.n1199 VCC.n1049 0.00822143
R2427 VCC.n1231 VCC.n1045 0.00822143
R2428 VCC.n1234 VCC.n1233 0.00822143
R2429 VCC.n1265 VCC.n1264 0.00822143
R2430 VCC.n1326 VCC.n988 0.00822143
R2431 VCC.n1366 VCC.n984 0.00822143
R2432 VCC.n1367 VCC.n980 0.00822143
R2433 VCC.n1399 VCC.n967 0.00822143
R2434 VCC.n1431 VCC.n931 0.00822143
R2435 VCC.n1472 VCC.n920 0.00822143
R2436 VCC.n1667 VCC.n1664 0.00822143
R2437 VCC.n1717 VCC.n1649 0.00822143
R2438 VCC.n1757 VCC.n1607 0.00822143
R2439 VCC.n1789 VCC.n1603 0.00822143
R2440 VCC.n1792 VCC.n1791 0.00822143
R2441 VCC.n1822 VCC.n1821 0.00822143
R2442 VCC.n1883 VCC.n1545 0.00822143
R2443 VCC.n1924 VCC.n1541 0.00822143
R2444 VCC.n1925 VCC.n1537 0.00822143
R2445 VCC.n1965 VCC.n1520 0.00822143
R2446 VCC.n1995 VCC.n1492 0.00822143
R2447 VCC.n2026 VCC.n1474 0.00822143
R2448 VCC.n103 VCC.n102 0.00822143
R2449 VCC.n107 VCC.n106 0.00822143
R2450 VCC.n175 VCC.n174 0.00822143
R2451 VCC.n171 VCC.n170 0.00822143
R2452 VCC.n169 VCC.n168 0.00822143
R2453 VCC.n160 VCC.n151 0.00822143
R2454 VCC.n354 VCC.n344 0.00822143
R2455 VCC.n365 VCC.n364 0.00822143
R2456 VCC.n587 VCC.n542 0.00764286
R2457 VCC.n602 VCC.n601 0.00764286
R2458 VCC.n642 VCC.n640 0.00764286
R2459 VCC.n639 VCC.n511 0.00764286
R2460 VCC.n650 VCC.n500 0.00764286
R2461 VCC.n558 VCC.n555 0.00764286
R2462 VCC.n600 VCC.n541 0.00764286
R2463 VCC.n610 VCC.n538 0.00764286
R2464 VCC.n626 VCC.n530 0.00764286
R2465 VCC.n645 VCC.n514 0.00764286
R2466 VCC.n641 VCC.n512 0.00764286
R2467 VCC.n483 VCC.n477 0.00764286
R2468 VCC.n770 VCC.n769 0.00764286
R2469 VCC.n766 VCC.n451 0.00764286
R2470 VCC.n777 VCC.n439 0.00764286
R2471 VCC.n720 VCC.n719 0.00764286
R2472 VCC.n734 VCC.n469 0.00764286
R2473 VCC.n735 VCC.n466 0.00764286
R2474 VCC.n740 VCC.n739 0.00764286
R2475 VCC.n768 VCC.n455 0.00764286
R2476 VCC.n813 VCC.n433 0.00764286
R2477 VCC.n843 VCC.n419 0.00764286
R2478 VCC.n882 VCC.n393 0.00764286
R2479 VCC.n816 VCC.n429 0.00764286
R2480 VCC.n846 VCC.n845 0.00764286
R2481 VCC.n853 VCC.n412 0.00764286
R2482 VCC.n849 VCC.n848 0.00764286
R2483 VCC.n872 VCC.n400 0.00764286
R2484 VCC.n886 VCC.n394 0.00764286
R2485 VCC.n1139 VCC.n1094 0.00764286
R2486 VCC.n1154 VCC.n1153 0.00764286
R2487 VCC.n1194 VCC.n1192 0.00764286
R2488 VCC.n1191 VCC.n1063 0.00764286
R2489 VCC.n1202 VCC.n1052 0.00764286
R2490 VCC.n1110 VCC.n1107 0.00764286
R2491 VCC.n1152 VCC.n1093 0.00764286
R2492 VCC.n1162 VCC.n1090 0.00764286
R2493 VCC.n1178 VCC.n1082 0.00764286
R2494 VCC.n1197 VCC.n1066 0.00764286
R2495 VCC.n1193 VCC.n1064 0.00764286
R2496 VCC.n1035 VCC.n1029 0.00764286
R2497 VCC.n1322 VCC.n1321 0.00764286
R2498 VCC.n1318 VCC.n1003 0.00764286
R2499 VCC.n1329 VCC.n991 0.00764286
R2500 VCC.n1272 VCC.n1271 0.00764286
R2501 VCC.n1286 VCC.n1021 0.00764286
R2502 VCC.n1287 VCC.n1018 0.00764286
R2503 VCC.n1292 VCC.n1291 0.00764286
R2504 VCC.n1320 VCC.n1007 0.00764286
R2505 VCC.n1365 VCC.n985 0.00764286
R2506 VCC.n1395 VCC.n971 0.00764286
R2507 VCC.n1434 VCC.n945 0.00764286
R2508 VCC.n1368 VCC.n981 0.00764286
R2509 VCC.n1398 VCC.n1397 0.00764286
R2510 VCC.n1405 VCC.n964 0.00764286
R2511 VCC.n1401 VCC.n1400 0.00764286
R2512 VCC.n1424 VCC.n952 0.00764286
R2513 VCC.n1438 VCC.n946 0.00764286
R2514 VCC.n1961 VCC.n1524 0.00764286
R2515 VCC.n1505 VCC.n1504 0.00764286
R2516 VCC.n1926 VCC.n1538 0.00764286
R2517 VCC.n1964 VCC.n1963 0.00764286
R2518 VCC.n1957 VCC.n1956 0.00764286
R2519 VCC.n1968 VCC.n1517 0.00764286
R2520 VCC.n1976 VCC.n1975 0.00764286
R2521 VCC.n1502 VCC.n1498 0.00764286
R2522 VCC.n1592 VCC.n1586 0.00764286
R2523 VCC.n1879 VCC.n1878 0.00764286
R2524 VCC.n1875 VCC.n1560 0.00764286
R2525 VCC.n1886 VCC.n1548 0.00764286
R2526 VCC.n1829 VCC.n1828 0.00764286
R2527 VCC.n1843 VCC.n1578 0.00764286
R2528 VCC.n1844 VCC.n1575 0.00764286
R2529 VCC.n1849 VCC.n1848 0.00764286
R2530 VCC.n1877 VCC.n1564 0.00764286
R2531 VCC.n1923 VCC.n1542 0.00764286
R2532 VCC.n1697 VCC.n1652 0.00764286
R2533 VCC.n1712 VCC.n1711 0.00764286
R2534 VCC.n1752 VCC.n1750 0.00764286
R2535 VCC.n1749 VCC.n1621 0.00764286
R2536 VCC.n1760 VCC.n1610 0.00764286
R2537 VCC.n1668 VCC.n1665 0.00764286
R2538 VCC.n1710 VCC.n1651 0.00764286
R2539 VCC.n1720 VCC.n1648 0.00764286
R2540 VCC.n1736 VCC.n1640 0.00764286
R2541 VCC.n1755 VCC.n1624 0.00764286
R2542 VCC.n1751 VCC.n1622 0.00764286
R2543 VCC.n57 VCC.n56 0.00764286
R2544 VCC.n205 VCC.n204 0.00764286
R2545 VCC.n208 VCC.n207 0.00764286
R2546 VCC.n210 VCC.n209 0.00764286
R2547 VCC.n98 VCC.n97 0.00764286
R2548 VCC.n101 VCC.n100 0.00764286
R2549 VCC.n113 VCC.n112 0.00764286
R2550 VCC.n179 VCC.n178 0.00764286
R2551 VCC.n131 VCC.n130 0.00764286
R2552 VCC.n117 VCC.n116 0.00764286
R2553 VCC.n257 VCC.n256 0.00764286
R2554 VCC.n314 VCC.n313 0.00764286
R2555 VCC.n167 VCC.n163 0.00764286
R2556 VCC.n142 VCC.n141 0.00764286
R2557 VCC.n148 VCC.n147 0.00764286
R2558 VCC.n341 VCC.n337 0.00764286
R2559 VCC.n569 VCC.n562 0.00675
R2560 VCC.n612 VCC.n536 0.00675
R2561 VCC.n643 VCC.n642 0.00675
R2562 VCC.n664 VCC.n504 0.00675
R2563 VCC.n605 VCC.n541 0.00675
R2564 VCC.n611 VCC.n537 0.00675
R2565 VCC.n641 VCC.n515 0.00675
R2566 VCC.n649 VCC.n498 0.00675
R2567 VCC.n678 VCC.n494 0.00675
R2568 VCC.n718 VCC.n717 0.00675
R2569 VCC.n733 VCC.n470 0.00675
R2570 VCC.n769 VCC.n767 0.00675
R2571 VCC.n799 VCC.n443 0.00675
R2572 VCC.n680 VCC.n492 0.00675
R2573 VCC.n711 VCC.n479 0.00675
R2574 VCC.n719 VCC.n715 0.00675
R2575 VCC.n772 VCC.n454 0.00675
R2576 VCC.n768 VCC.n452 0.00675
R2577 VCC.n419 VCC.n410 0.00675
R2578 VCC.n413 VCC.n411 0.00675
R2579 VCC.n887 VCC.n393 0.00675
R2580 VCC.n417 VCC.n412 0.00675
R2581 VCC.n852 VCC.n414 0.00675
R2582 VCC.n400 VCC.n397 0.00675
R2583 VCC.n886 VCC.n885 0.00675
R2584 VCC.n884 VCC.n880 0.00675
R2585 VCC.n1121 VCC.n1114 0.00675
R2586 VCC.n1164 VCC.n1088 0.00675
R2587 VCC.n1195 VCC.n1194 0.00675
R2588 VCC.n1216 VCC.n1056 0.00675
R2589 VCC.n1157 VCC.n1093 0.00675
R2590 VCC.n1163 VCC.n1089 0.00675
R2591 VCC.n1193 VCC.n1067 0.00675
R2592 VCC.n1201 VCC.n1050 0.00675
R2593 VCC.n1230 VCC.n1046 0.00675
R2594 VCC.n1270 VCC.n1269 0.00675
R2595 VCC.n1285 VCC.n1022 0.00675
R2596 VCC.n1321 VCC.n1319 0.00675
R2597 VCC.n1351 VCC.n995 0.00675
R2598 VCC.n1232 VCC.n1044 0.00675
R2599 VCC.n1263 VCC.n1031 0.00675
R2600 VCC.n1271 VCC.n1267 0.00675
R2601 VCC.n1324 VCC.n1006 0.00675
R2602 VCC.n1320 VCC.n1004 0.00675
R2603 VCC.n971 VCC.n962 0.00675
R2604 VCC.n965 VCC.n963 0.00675
R2605 VCC.n1439 VCC.n945 0.00675
R2606 VCC.n969 VCC.n964 0.00675
R2607 VCC.n1404 VCC.n966 0.00675
R2608 VCC.n952 VCC.n949 0.00675
R2609 VCC.n1438 VCC.n1437 0.00675
R2610 VCC.n1436 VCC.n1432 0.00675
R2611 VCC.n1958 VCC.n1524 0.00675
R2612 VCC.n1970 VCC.n1518 0.00675
R2613 VCC.n1504 VCC.n1500 0.00675
R2614 VCC.n1957 VCC.n1522 0.00675
R2615 VCC.n1969 VCC.n1519 0.00675
R2616 VCC.n1975 VCC.n1497 0.00675
R2617 VCC.n1503 VCC.n1502 0.00675
R2618 VCC.n1996 VCC.n1495 0.00675
R2619 VCC.n1827 VCC.n1826 0.00675
R2620 VCC.n1842 VCC.n1579 0.00675
R2621 VCC.n1878 VCC.n1876 0.00675
R2622 VCC.n1909 VCC.n1552 0.00675
R2623 VCC.n1790 VCC.n1602 0.00675
R2624 VCC.n1820 VCC.n1588 0.00675
R2625 VCC.n1828 VCC.n1824 0.00675
R2626 VCC.n1881 VCC.n1563 0.00675
R2627 VCC.n1877 VCC.n1561 0.00675
R2628 VCC.n1679 VCC.n1672 0.00675
R2629 VCC.n1722 VCC.n1646 0.00675
R2630 VCC.n1753 VCC.n1752 0.00675
R2631 VCC.n1774 VCC.n1614 0.00675
R2632 VCC.n1715 VCC.n1651 0.00675
R2633 VCC.n1721 VCC.n1647 0.00675
R2634 VCC.n1751 VCC.n1625 0.00675
R2635 VCC.n1759 VCC.n1608 0.00675
R2636 VCC.n1788 VCC.n1604 0.00675
R2637 VCC.n62 VCC.n61 0.00675
R2638 VCC.n76 VCC.n64 0.00675
R2639 VCC.n206 VCC.n205 0.00675
R2640 VCC.n221 VCC.n217 0.00675
R2641 VCC.n85 VCC.n84 0.00675
R2642 VCC.n95 VCC.n94 0.00675
R2643 VCC.n99 VCC.n98 0.00675
R2644 VCC.n133 VCC.n132 0.00675
R2645 VCC.n130 VCC.n129 0.00675
R2646 VCC.n269 VCC.n257 0.00675
R2647 VCC.n273 VCC.n272 0.00675
R2648 VCC.n326 VCC.n314 0.00675
R2649 VCC.n141 VCC.n140 0.00675
R2650 VCC.n144 VCC.n143 0.00675
R2651 VCC.n341 VCC.n340 0.00675
R2652 VCC.n346 VCC.n345 0.00675
R2653 VCC.n348 VCC.n347 0.00675
R2654 VCC.n572 VCC.n562 0.00585714
R2655 VCC.n604 VCC.n603 0.00585714
R2656 VCC.n524 VCC.n516 0.00585714
R2657 VCC.n553 VCC.n540 0.00585714
R2658 VCC.n611 VCC.n610 0.00585714
R2659 VCC.n697 VCC.n686 0.00585714
R2660 VCC.n694 VCC.n686 0.00585714
R2661 VCC.n721 VCC.n478 0.00585714
R2662 VCC.n756 VCC.n456 0.00585714
R2663 VCC.n800 VCC.n799 0.00585714
R2664 VCC.n739 VCC.n454 0.00585714
R2665 VCC.n776 VCC.n437 0.00585714
R2666 VCC.n818 VCC.n424 0.00585714
R2667 VCC.n855 VCC.n854 0.00585714
R2668 VCC.n876 VCC.n875 0.00585714
R2669 VCC.n888 VCC.n392 0.00585714
R2670 VCC.n383 VCC.n374 0.00585714
R2671 VCC.n377 VCC.n375 0.00585714
R2672 VCC.n427 VCC.n416 0.00585714
R2673 VCC.n849 VCC.n414 0.00585714
R2674 VCC.n877 VCC.n397 0.00585714
R2675 VCC.n1124 VCC.n1114 0.00585714
R2676 VCC.n1156 VCC.n1155 0.00585714
R2677 VCC.n1076 VCC.n1068 0.00585714
R2678 VCC.n1105 VCC.n1092 0.00585714
R2679 VCC.n1163 VCC.n1162 0.00585714
R2680 VCC.n1249 VCC.n1238 0.00585714
R2681 VCC.n1246 VCC.n1238 0.00585714
R2682 VCC.n1273 VCC.n1030 0.00585714
R2683 VCC.n1308 VCC.n1008 0.00585714
R2684 VCC.n1352 VCC.n1351 0.00585714
R2685 VCC.n1291 VCC.n1006 0.00585714
R2686 VCC.n1328 VCC.n989 0.00585714
R2687 VCC.n1370 VCC.n976 0.00585714
R2688 VCC.n1407 VCC.n1406 0.00585714
R2689 VCC.n1428 VCC.n1427 0.00585714
R2690 VCC.n1440 VCC.n944 0.00585714
R2691 VCC.n935 VCC.n928 0.00585714
R2692 VCC.n1457 VCC.n929 0.00585714
R2693 VCC.n979 VCC.n968 0.00585714
R2694 VCC.n1401 VCC.n966 0.00585714
R2695 VCC.n1429 VCC.n949 0.00585714
R2696 VCC.n1928 VCC.n1532 0.00585714
R2697 VCC.n1955 VCC.n1954 0.00585714
R2698 VCC.n1992 VCC.n1499 0.00585714
R2699 VCC.n1991 VCC.n1990 0.00585714
R2700 VCC.n1488 VCC.n1485 0.00585714
R2701 VCC.n2007 VCC.n2006 0.00585714
R2702 VCC.n1536 VCC.n1521 0.00585714
R2703 VCC.n1969 VCC.n1968 0.00585714
R2704 VCC.n1993 VCC.n1497 0.00585714
R2705 VCC.n1796 VCC.n1601 0.00585714
R2706 VCC.n1803 VCC.n1796 0.00585714
R2707 VCC.n1830 VCC.n1587 0.00585714
R2708 VCC.n1865 VCC.n1565 0.00585714
R2709 VCC.n1910 VCC.n1909 0.00585714
R2710 VCC.n1848 VCC.n1563 0.00585714
R2711 VCC.n1885 VCC.n1546 0.00585714
R2712 VCC.n1682 VCC.n1672 0.00585714
R2713 VCC.n1714 VCC.n1713 0.00585714
R2714 VCC.n1634 VCC.n1626 0.00585714
R2715 VCC.n1663 VCC.n1650 0.00585714
R2716 VCC.n1721 VCC.n1720 0.00585714
R2717 VCC.n36 VCC.n35 0.00585714
R2718 VCC.n37 VCC.n36 0.00585714
R2719 VCC.n60 VCC.n59 0.00585714
R2720 VCC.n202 VCC.n201 0.00585714
R2721 VCC.n217 VCC.n216 0.00585714
R2722 VCC.n178 VCC.n133 0.00585714
R2723 VCC.n127 VCC.n126 0.00585714
R2724 VCC.n239 VCC.n238 0.00585714
R2725 VCC.n271 VCC.n270 0.00585714
R2726 VCC.n330 VCC.n329 0.00585714
R2727 VCC.n328 VCC.n327 0.00585714
R2728 VCC.n294 VCC.n293 0.00585714
R2729 VCC.n290 VCC.n289 0.00585714
R2730 VCC.n159 VCC.n158 0.00585714
R2731 VCC.n148 VCC.n144 0.00585714
R2732 VCC.n340 VCC.n339 0.00585714
R2733 VCC.n665 VCC.n503 0.00496429
R2734 VCC.n665 VCC.n664 0.00496429
R2735 VCC.n582 VCC.n555 0.00496429
R2736 VCC.n585 VCC.n553 0.00496429
R2737 VCC.n530 VCC.n514 0.00496429
R2738 VCC.n672 VCC.n498 0.00496429
R2739 VCC.n675 VCC.n494 0.00496429
R2740 VCC.n694 VCC.n693 0.00496429
R2741 VCC.n684 VCC.n492 0.00496429
R2742 VCC.n711 VCC.n710 0.00496429
R2743 VCC.n735 VCC.n734 0.00496429
R2744 VCC.n807 VCC.n437 0.00496429
R2745 VCC.n810 VCC.n433 0.00496429
R2746 VCC.n825 VCC.n429 0.00496429
R2747 VCC.n830 VCC.n427 0.00496429
R2748 VCC.n395 VCC.n380 0.00496429
R2749 VCC.n901 VCC.n380 0.00496429
R2750 VCC.n904 VCC.n367 0.00496429
R2751 VCC.n1217 VCC.n1055 0.00496429
R2752 VCC.n1217 VCC.n1216 0.00496429
R2753 VCC.n1134 VCC.n1107 0.00496429
R2754 VCC.n1137 VCC.n1105 0.00496429
R2755 VCC.n1082 VCC.n1066 0.00496429
R2756 VCC.n1224 VCC.n1050 0.00496429
R2757 VCC.n1227 VCC.n1046 0.00496429
R2758 VCC.n1246 VCC.n1245 0.00496429
R2759 VCC.n1236 VCC.n1044 0.00496429
R2760 VCC.n1263 VCC.n1262 0.00496429
R2761 VCC.n1287 VCC.n1286 0.00496429
R2762 VCC.n1359 VCC.n989 0.00496429
R2763 VCC.n1362 VCC.n985 0.00496429
R2764 VCC.n1377 VCC.n981 0.00496429
R2765 VCC.n1382 VCC.n979 0.00496429
R2766 VCC.n947 VCC.n932 0.00496429
R2767 VCC.n1453 VCC.n932 0.00496429
R2768 VCC.n1456 VCC.n921 0.00496429
R2769 VCC.n1936 VCC.n1538 0.00496429
R2770 VCC.n1939 VCC.n1536 0.00496429
R2771 VCC.n1997 VCC.n1493 0.00496429
R2772 VCC.n2000 VCC.n1493 0.00496429
R2773 VCC.n2003 VCC.n1475 0.00496429
R2774 VCC.n1803 VCC.n1802 0.00496429
R2775 VCC.n1794 VCC.n1602 0.00496429
R2776 VCC.n1820 VCC.n1819 0.00496429
R2777 VCC.n1844 VCC.n1843 0.00496429
R2778 VCC.n1917 VCC.n1546 0.00496429
R2779 VCC.n1920 VCC.n1542 0.00496429
R2780 VCC.n1775 VCC.n1613 0.00496429
R2781 VCC.n1775 VCC.n1774 0.00496429
R2782 VCC.n1692 VCC.n1665 0.00496429
R2783 VCC.n1695 VCC.n1663 0.00496429
R2784 VCC.n1640 VCC.n1624 0.00496429
R2785 VCC.n1782 VCC.n1608 0.00496429
R2786 VCC.n1785 VCC.n1604 0.00496429
R2787 VCC.n38 VCC.n37 0.00496429
R2788 VCC.n86 VCC.n85 0.00496429
R2789 VCC.n94 VCC.n93 0.00496429
R2790 VCC.n112 VCC.n101 0.00496429
R2791 VCC.n126 VCC.n125 0.00496429
R2792 VCC.n118 VCC.n117 0.00496429
R2793 VCC.n167 VCC.n166 0.00496429
R2794 VCC.n159 VCC.n156 0.00496429
R2795 VCC.n353 VCC.n349 0.00496429
R2796 VCC.n353 VCC.n352 0.00496429
R2797 VCC.n363 VCC.n361 0.00496429
R2798 VCC.n609 VCC.n608 0.00486429
R2799 VCC.n623 VCC.n531 0.00486429
R2800 VCC.n625 VCC.n624 0.00486429
R2801 VCC.n646 VCC.n513 0.00486429
R2802 VCC.n736 VCC.n468 0.00486429
R2803 VCC.n746 VCC.n737 0.00486429
R2804 VCC.n745 VCC.n738 0.00486429
R2805 VCC.n773 VCC.n453 0.00486429
R2806 VCC.n851 VCC.n850 0.00486429
R2807 VCC.n869 VCC.n401 0.00486429
R2808 VCC.n871 VCC.n870 0.00486429
R2809 VCC.n878 VCC.n396 0.00486429
R2810 VCC.n1161 VCC.n1160 0.00486429
R2811 VCC.n1175 VCC.n1083 0.00486429
R2812 VCC.n1177 VCC.n1176 0.00486429
R2813 VCC.n1198 VCC.n1065 0.00486429
R2814 VCC.n1288 VCC.n1020 0.00486429
R2815 VCC.n1298 VCC.n1289 0.00486429
R2816 VCC.n1297 VCC.n1290 0.00486429
R2817 VCC.n1325 VCC.n1005 0.00486429
R2818 VCC.n1403 VCC.n1402 0.00486429
R2819 VCC.n1421 VCC.n953 0.00486429
R2820 VCC.n1423 VCC.n1422 0.00486429
R2821 VCC.n1430 VCC.n948 0.00486429
R2822 VCC.n1719 VCC.n1718 0.00486429
R2823 VCC.n1733 VCC.n1641 0.00486429
R2824 VCC.n1735 VCC.n1734 0.00486429
R2825 VCC.n1756 VCC.n1623 0.00486429
R2826 VCC.n1845 VCC.n1577 0.00486429
R2827 VCC.n1855 VCC.n1846 0.00486429
R2828 VCC.n1854 VCC.n1847 0.00486429
R2829 VCC.n1882 VCC.n1562 0.00486429
R2830 VCC.n1967 VCC.n1966 0.00486429
R2831 VCC.n1974 VCC.n1516 0.00486429
R2832 VCC.n1978 VCC.n1977 0.00486429
R2833 VCC.n1994 VCC.n1496 0.00486429
R2834 VCC.n111 VCC.n108 0.00486429
R2835 VCC.n110 VCC.n109 0.00486429
R2836 VCC.n135 VCC.n134 0.00486429
R2837 VCC.n177 VCC.n176 0.00486429
R2838 VCC.n150 VCC.n149 0.00486429
R2839 VCC.n138 VCC.n137 0.00486429
R2840 VCC.n136 VCC.n0 0.00486429
R2841 VCC.n343 VCC.n342 0.00486429
R2842 VCC.n569 VCC.n568 0.00407143
R2843 VCC.n616 VCC.n534 0.00407143
R2844 VCC.n621 VCC.n617 0.00407143
R2845 VCC.n671 VCC.n500 0.00407143
R2846 VCC.n622 VCC.n532 0.00407143
R2847 VCC.n743 VCC.n462 0.00407143
R2848 VCC.n800 VCC.n442 0.00407143
R2849 VCC.n744 VCC.n741 0.00407143
R2850 VCC.n1121 VCC.n1120 0.00407143
R2851 VCC.n1168 VCC.n1086 0.00407143
R2852 VCC.n1173 VCC.n1169 0.00407143
R2853 VCC.n1223 VCC.n1052 0.00407143
R2854 VCC.n1174 VCC.n1084 0.00407143
R2855 VCC.n1295 VCC.n1014 0.00407143
R2856 VCC.n1352 VCC.n994 0.00407143
R2857 VCC.n1296 VCC.n1293 0.00407143
R2858 VCC.n1852 VCC.n1571 0.00407143
R2859 VCC.n1910 VCC.n1551 0.00407143
R2860 VCC.n1853 VCC.n1850 0.00407143
R2861 VCC.n1679 VCC.n1678 0.00407143
R2862 VCC.n1726 VCC.n1644 0.00407143
R2863 VCC.n1731 VCC.n1727 0.00407143
R2864 VCC.n1781 VCC.n1610 0.00407143
R2865 VCC.n1732 VCC.n1642 0.00407143
R2866 VCC.n187 VCC.n184 0.00407143
R2867 VCC.n216 VCC.n215 0.00407143
R2868 VCC.n181 VCC.n180 0.00407143
R2869 VCC.n609 VCC.n531 0.00318571
R2870 VCC.n625 VCC.n513 0.00318571
R2871 VCC.n737 VCC.n736 0.00318571
R2872 VCC.n738 VCC.n453 0.00318571
R2873 VCC.n850 VCC.n401 0.00318571
R2874 VCC.n871 VCC.n396 0.00318571
R2875 VCC.n1161 VCC.n1083 0.00318571
R2876 VCC.n1177 VCC.n1065 0.00318571
R2877 VCC.n1289 VCC.n1288 0.00318571
R2878 VCC.n1290 VCC.n1005 0.00318571
R2879 VCC.n1402 VCC.n953 0.00318571
R2880 VCC.n1423 VCC.n948 0.00318571
R2881 VCC.n1719 VCC.n1641 0.00318571
R2882 VCC.n1735 VCC.n1623 0.00318571
R2883 VCC.n1846 VCC.n1845 0.00318571
R2884 VCC.n1847 VCC.n1562 0.00318571
R2885 VCC.n1967 VCC.n1516 0.00318571
R2886 VCC.n1977 VCC.n1496 0.00318571
R2887 VCC.n111 VCC.n110 0.00318571
R2888 VCC.n177 VCC.n135 0.00318571
R2889 VCC.n149 VCC.n138 0.00318571
R2890 VCC.n342 VCC.n0 0.00318571
R2891 VCC.n586 VCC.n551 0.00317857
R2892 VCC.n628 VCC.n523 0.00317857
R2893 VCC.n671 VCC.n670 0.00317857
R2894 VCC.n676 VCC.n495 0.00317857
R2895 VCC.n582 VCC.n556 0.00317857
R2896 VCC.n585 VCC.n552 0.00317857
R2897 VCC.n627 VCC.n529 0.00317857
R2898 VCC.n672 VCC.n499 0.00317857
R2899 VCC.n675 VCC.n496 0.00317857
R2900 VCC.n698 VCC.n491 0.00317857
R2901 VCC.n709 VCC.n482 0.00317857
R2902 VCC.n709 VCC.n708 0.00317857
R2903 VCC.n471 VCC.n464 0.00317857
R2904 VCC.n749 VCC.n465 0.00317857
R2905 VCC.n755 VCC.n754 0.00317857
R2906 VCC.n806 VCC.n439 0.00317857
R2907 VCC.n806 VCC.n805 0.00317857
R2908 VCC.n811 VCC.n434 0.00317857
R2909 VCC.n685 VCC.n684 0.00317857
R2910 VCC.n710 VCC.n481 0.00317857
R2911 VCC.n748 VCC.n747 0.00317857
R2912 VCC.n807 VCC.n438 0.00317857
R2913 VCC.n810 VCC.n435 0.00317857
R2914 VCC.n824 VCC.n823 0.00317857
R2915 VCC.n829 VCC.n425 0.00317857
R2916 VCC.n874 VCC.n398 0.00317857
R2917 VCC.n883 VCC.n882 0.00317857
R2918 VCC.n900 VCC.n899 0.00317857
R2919 VCC.n378 VCC.n377 0.00317857
R2920 VCC.n378 VCC.n368 0.00317857
R2921 VCC.n825 VCC.n430 0.00317857
R2922 VCC.n831 VCC.n830 0.00317857
R2923 VCC.n873 VCC.n399 0.00317857
R2924 VCC.n901 VCC.n381 0.00317857
R2925 VCC.n905 VCC.n904 0.00317857
R2926 VCC.n1138 VCC.n1103 0.00317857
R2927 VCC.n1180 VCC.n1075 0.00317857
R2928 VCC.n1223 VCC.n1222 0.00317857
R2929 VCC.n1228 VCC.n1047 0.00317857
R2930 VCC.n1134 VCC.n1108 0.00317857
R2931 VCC.n1137 VCC.n1104 0.00317857
R2932 VCC.n1179 VCC.n1081 0.00317857
R2933 VCC.n1224 VCC.n1051 0.00317857
R2934 VCC.n1227 VCC.n1048 0.00317857
R2935 VCC.n1250 VCC.n1043 0.00317857
R2936 VCC.n1261 VCC.n1034 0.00317857
R2937 VCC.n1261 VCC.n1260 0.00317857
R2938 VCC.n1023 VCC.n1016 0.00317857
R2939 VCC.n1301 VCC.n1017 0.00317857
R2940 VCC.n1307 VCC.n1306 0.00317857
R2941 VCC.n1358 VCC.n991 0.00317857
R2942 VCC.n1358 VCC.n1357 0.00317857
R2943 VCC.n1363 VCC.n986 0.00317857
R2944 VCC.n1237 VCC.n1236 0.00317857
R2945 VCC.n1262 VCC.n1033 0.00317857
R2946 VCC.n1300 VCC.n1299 0.00317857
R2947 VCC.n1359 VCC.n990 0.00317857
R2948 VCC.n1362 VCC.n987 0.00317857
R2949 VCC.n1376 VCC.n1375 0.00317857
R2950 VCC.n1381 VCC.n977 0.00317857
R2951 VCC.n1426 VCC.n950 0.00317857
R2952 VCC.n1435 VCC.n1434 0.00317857
R2953 VCC.n1452 VCC.n1451 0.00317857
R2954 VCC.n1458 VCC.n1457 0.00317857
R2955 VCC.n1458 VCC.n922 0.00317857
R2956 VCC.n1377 VCC.n982 0.00317857
R2957 VCC.n1383 VCC.n1382 0.00317857
R2958 VCC.n1425 VCC.n951 0.00317857
R2959 VCC.n1453 VCC.n933 0.00317857
R2960 VCC.n1459 VCC.n1456 0.00317857
R2961 VCC.n1935 VCC.n1934 0.00317857
R2962 VCC.n1941 VCC.n1535 0.00317857
R2963 VCC.n1980 VCC.n1514 0.00317857
R2964 VCC.n1505 VCC.n1494 0.00317857
R2965 VCC.n1999 VCC.n1484 0.00317857
R2966 VCC.n2006 VCC.n2005 0.00317857
R2967 VCC.n2005 VCC.n1476 0.00317857
R2968 VCC.n1936 VCC.n1539 0.00317857
R2969 VCC.n1940 VCC.n1939 0.00317857
R2970 VCC.n1979 VCC.n1515 0.00317857
R2971 VCC.n2000 VCC.n1486 0.00317857
R2972 VCC.n2004 VCC.n2003 0.00317857
R2973 VCC.n1807 VCC.n1600 0.00317857
R2974 VCC.n1818 VCC.n1591 0.00317857
R2975 VCC.n1818 VCC.n1817 0.00317857
R2976 VCC.n1580 VCC.n1573 0.00317857
R2977 VCC.n1858 VCC.n1574 0.00317857
R2978 VCC.n1864 VCC.n1863 0.00317857
R2979 VCC.n1916 VCC.n1548 0.00317857
R2980 VCC.n1916 VCC.n1915 0.00317857
R2981 VCC.n1921 VCC.n1543 0.00317857
R2982 VCC.n1806 VCC.n1794 0.00317857
R2983 VCC.n1819 VCC.n1590 0.00317857
R2984 VCC.n1857 VCC.n1856 0.00317857
R2985 VCC.n1917 VCC.n1547 0.00317857
R2986 VCC.n1920 VCC.n1544 0.00317857
R2987 VCC.n1696 VCC.n1661 0.00317857
R2988 VCC.n1738 VCC.n1633 0.00317857
R2989 VCC.n1781 VCC.n1780 0.00317857
R2990 VCC.n1786 VCC.n1605 0.00317857
R2991 VCC.n1692 VCC.n1666 0.00317857
R2992 VCC.n1695 VCC.n1662 0.00317857
R2993 VCC.n1737 VCC.n1639 0.00317857
R2994 VCC.n1782 VCC.n1609 0.00317857
R2995 VCC.n1785 VCC.n1606 0.00317857
R2996 VCC.n24 VCC.n23 0.00317857
R2997 VCC.n42 VCC.n41 0.00317857
R2998 VCC.n43 VCC.n42 0.00317857
R2999 VCC.n78 VCC.n77 0.00317857
R3000 VCC.n83 VCC.n82 0.00317857
R3001 VCC.n189 VCC.n188 0.00317857
R3002 VCC.n211 VCC.n210 0.00317857
R3003 VCC.n212 VCC.n211 0.00317857
R3004 VCC.n220 VCC.n219 0.00317857
R3005 VCC.n87 VCC.n86 0.00317857
R3006 VCC.n93 VCC.n92 0.00317857
R3007 VCC.n115 VCC.n114 0.00317857
R3008 VCC.n125 VCC.n124 0.00317857
R3009 VCC.n119 VCC.n118 0.00317857
R3010 VCC.n235 VCC.n234 0.00317857
R3011 VCC.n252 VCC.n251 0.00317857
R3012 VCC.n332 VCC.n331 0.00317857
R3013 VCC.n313 VCC.n312 0.00317857
R3014 VCC.n310 VCC.n309 0.00317857
R3015 VCC.n289 VCC.n288 0.00317857
R3016 VCC.n288 VCC.n287 0.00317857
R3017 VCC.n166 VCC.n165 0.00317857
R3018 VCC.n156 VCC.n155 0.00317857
R3019 VCC.n336 VCC.n335 0.00317857
R3020 VCC.n352 VCC.n351 0.00317857
R3021 VCC.n361 VCC.n360 0.00317857
R3022 VCC.n581 VCC.n580 0.00228571
R3023 VCC.n588 VCC.n586 0.00228571
R3024 VCC.n528 VCC.n527 0.00228571
R3025 VCC.n644 VCC.n516 0.00228571
R3026 VCC.n718 VCC.n478 0.00228571
R3027 VCC.n844 VCC.n843 0.00228571
R3028 VCC.n855 VCC.n410 0.00228571
R3029 VCC.n867 VCC.n404 0.00228571
R3030 VCC.n888 VCC.n887 0.00228571
R3031 VCC.n868 VCC.n402 0.00228571
R3032 VCC.n1133 VCC.n1132 0.00228571
R3033 VCC.n1140 VCC.n1138 0.00228571
R3034 VCC.n1080 VCC.n1079 0.00228571
R3035 VCC.n1196 VCC.n1068 0.00228571
R3036 VCC.n1270 VCC.n1030 0.00228571
R3037 VCC.n1396 VCC.n1395 0.00228571
R3038 VCC.n1407 VCC.n962 0.00228571
R3039 VCC.n1419 VCC.n956 0.00228571
R3040 VCC.n1440 VCC.n1439 0.00228571
R3041 VCC.n1420 VCC.n954 0.00228571
R3042 VCC.n1962 VCC.n1961 0.00228571
R3043 VCC.n1958 VCC.n1954 0.00228571
R3044 VCC.n1971 VCC.n1512 0.00228571
R3045 VCC.n1990 VCC.n1500 0.00228571
R3046 VCC.n1973 VCC.n1972 0.00228571
R3047 VCC.n1827 VCC.n1587 0.00228571
R3048 VCC.n1691 VCC.n1690 0.00228571
R3049 VCC.n1698 VCC.n1696 0.00228571
R3050 VCC.n1638 VCC.n1637 0.00228571
R3051 VCC.n1754 VCC.n1626 0.00228571
R3052 VCC.n61 VCC.n60 0.00228571
R3053 VCC.n256 VCC.n255 0.00228571
R3054 VCC.n270 VCC.n269 0.00228571
R3055 VCC.n275 VCC.n274 0.00228571
R3056 VCC.n327 VCC.n326 0.00228571
R3057 VCC.n146 VCC.n145 0.00228571
R3058 VCC.n583 VCC.n554 0.00217857
R3059 VCC.n584 VCC.n539 0.00217857
R3060 VCC.n673 VCC.n497 0.00217857
R3061 VCC.n674 VCC.n493 0.00217857
R3062 VCC.n683 VCC.n682 0.00217857
R3063 VCC.n712 VCC.n480 0.00217857
R3064 VCC.n808 VCC.n436 0.00217857
R3065 VCC.n809 VCC.n432 0.00217857
R3066 VCC.n826 VCC.n428 0.00217857
R3067 VCC.n827 VCC.n415 0.00217857
R3068 VCC.n902 VCC.n379 0.00217857
R3069 VCC.n903 VCC.n366 0.00217857
R3070 VCC.n1135 VCC.n1106 0.00217857
R3071 VCC.n1136 VCC.n1091 0.00217857
R3072 VCC.n1225 VCC.n1049 0.00217857
R3073 VCC.n1226 VCC.n1045 0.00217857
R3074 VCC.n1235 VCC.n1234 0.00217857
R3075 VCC.n1264 VCC.n1032 0.00217857
R3076 VCC.n1360 VCC.n988 0.00217857
R3077 VCC.n1361 VCC.n984 0.00217857
R3078 VCC.n1378 VCC.n980 0.00217857
R3079 VCC.n1379 VCC.n967 0.00217857
R3080 VCC.n1454 VCC.n931 0.00217857
R3081 VCC.n1455 VCC.n920 0.00217857
R3082 VCC.n1693 VCC.n1664 0.00217857
R3083 VCC.n1694 VCC.n1649 0.00217857
R3084 VCC.n1783 VCC.n1607 0.00217857
R3085 VCC.n1784 VCC.n1603 0.00217857
R3086 VCC.n1793 VCC.n1792 0.00217857
R3087 VCC.n1821 VCC.n1589 0.00217857
R3088 VCC.n1918 VCC.n1545 0.00217857
R3089 VCC.n1919 VCC.n1541 0.00217857
R3090 VCC.n1937 VCC.n1537 0.00217857
R3091 VCC.n1938 VCC.n1520 0.00217857
R3092 VCC.n2001 VCC.n1492 0.00217857
R3093 VCC.n2002 VCC.n1474 0.00217857
R3094 VCC.n104 VCC.n103 0.00217857
R3095 VCC.n106 VCC.n105 0.00217857
R3096 VCC.n174 VCC.n173 0.00217857
R3097 VCC.n172 VCC.n171 0.00217857
R3098 VCC.n168 VCC.n162 0.00217857
R3099 VCC.n161 VCC.n160 0.00217857
R3100 VCC.n355 VCC.n354 0.00217857
R3101 VCC.n364 VCC.n356 0.00217857
R3102 VCC.n580 VCC.n559 0.00139286
R3103 VCC.n603 VCC.n602 0.00139286
R3104 VCC.n620 VCC.n619 0.00139286
R3105 VCC.n660 VCC.n495 0.00139286
R3106 VCC.n618 VCC.n533 0.00139286
R3107 VCC.n716 VCC.n470 0.00139286
R3108 VCC.n771 VCC.n456 0.00139286
R3109 VCC.n898 VCC.n385 0.00139286
R3110 VCC.n909 VCC.n374 0.00139286
R3111 VCC.n1132 VCC.n1111 0.00139286
R3112 VCC.n1155 VCC.n1154 0.00139286
R3113 VCC.n1172 VCC.n1171 0.00139286
R3114 VCC.n1212 VCC.n1047 0.00139286
R3115 VCC.n1170 VCC.n1085 0.00139286
R3116 VCC.n1268 VCC.n1022 0.00139286
R3117 VCC.n1323 VCC.n1008 0.00139286
R3118 VCC.n1450 VCC.n937 0.00139286
R3119 VCC.n1463 VCC.n928 0.00139286
R3120 VCC.n2013 VCC.n2012 0.00139286
R3121 VCC.n1491 VCC.n1488 0.00139286
R3122 VCC.n1825 VCC.n1579 0.00139286
R3123 VCC.n1880 VCC.n1565 0.00139286
R3124 VCC.n1690 VCC.n1669 0.00139286
R3125 VCC.n1713 VCC.n1712 0.00139286
R3126 VCC.n1730 VCC.n1729 0.00139286
R3127 VCC.n1770 VCC.n1605 0.00139286
R3128 VCC.n1728 VCC.n1643 0.00139286
R3129 VCC.n64 VCC.n63 0.00139286
R3130 VCC.n203 VCC.n202 0.00139286
R3131 VCC.n308 VCC.n307 0.00139286
R3132 VCC.n293 VCC.n292 0.00139286
R3133 VCC.n2028 VCC.n2027 0.00054824
R3134 VSS.n2187 VSS.n12 106073
R3135 VSS.n1822 VSS.n12 54262.5
R3136 VSS.n2187 VSS.n10 12274.8
R3137 VSS.n2187 VSS.n11 12232.2
R3138 VSS.n2188 VSS.n2187 12232.2
R3139 VSS.n2187 VSS.n2186 12232.2
R3140 VSS.n1822 VSS.n1821 6909.46
R3141 VSS.n1821 VSS.t61 6273.77
R3142 VSS.n741 VSS.t66 4305.17
R3143 VSS.n1314 VSS.t12 4305.17
R3144 VSS.n2047 VSS.t5 4305.17
R3145 VSS.n1774 VSS.n12 3531.03
R3146 VSS.n1774 VSS.n1773 3531.03
R3147 VSS.t36 VSS.n12 3054.19
R3148 VSS.n1774 VSS.t49 3054.19
R3149 VSS.n1725 VSS.t64 2804.58
R3150 VSS.n1724 VSS.t65 2770.93
R3151 VSS.n1726 VSS.n1725 2671.38
R3152 VSS.t65 VSS.t23 2603.46
R3153 VSS.n1927 VSS.n12 2588.02
R3154 VSS.n1775 VSS.n1774 2588.02
R3155 VSS.n742 VSS.n741 2406.66
R3156 VSS.n1315 VSS.n1314 2406.66
R3157 VSS.n2048 VSS.n2047 2406.66
R3158 VSS.t57 VSS.n1771 2349.66
R3159 VSS.t48 VSS.t57 2304.76
R3160 VSS.t75 VSS.n787 1937.11
R3161 VSS.t72 VSS.n1360 1937.11
R3162 VSS.n167 VSS.t19 1937.11
R3163 VSS.n1823 VSS.t18 1930.89
R3164 VSS.t56 VSS.n1820 1930.89
R3165 VSS.n741 VSS.n740 1896.55
R3166 VSS.n1314 VSS.n1313 1896.55
R3167 VSS.n2047 VSS.n2046 1896.55
R3168 VSS.t60 VSS.t72 1892.74
R3169 VSS.t18 VSS.t0 1892.74
R3170 VSS.t19 VSS.t36 1892.74
R3171 VSS.t9 VSS.t56 1892.74
R3172 VSS.t49 VSS.t75 1892.74
R3173 VSS.n740 VSS.t69 1791.5
R3174 VSS.n1313 VSS.t15 1791.5
R3175 VSS.n2046 VSS.t4 1791.5
R3176 VSS.t69 VSS.t30 1683.22
R3177 VSS.t15 VSS.t26 1683.22
R3178 VSS.t4 VSS.t52 1683.22
R3179 VSS.t23 VSS.n1723 1560.55
R3180 VSS.n1772 VSS.t48 1331.97
R3181 VSS.n1772 VSS.t60 1093.85
R3182 VSS.t0 VSS.n1822 1093.85
R3183 VSS.n1821 VSS.t9 1093.85
R3184 VSS.t30 VSS.n739 1045.79
R3185 VSS.t26 VSS.n1312 1045.79
R3186 VSS.t52 VSS.n2045 1045.79
R3187 VSS.n1773 VSS.n788 1017.62
R3188 VSS.n1773 VSS.n1772 772.908
R3189 VSS.n868 VSS.t41 758.37
R3190 VSS.t41 VSS.t61 746.255
R3191 VSS.n739 VSS.n738 590.341
R3192 VSS.n639 VSS.n11 590.341
R3193 VSS.n1312 VSS.n1311 590.341
R3194 VSS.n2188 VSS.n6 590.341
R3195 VSS.n2045 VSS.n2044 590.341
R3196 VSS.n2186 VSS.n2185 590.341
R3197 VSS.n1723 VSS.n1722 590.341
R3198 VSS.n1628 VSS.n10 590.341
R3199 VSS.n441 VSS.n440 585
R3200 VSS.n440 VSS.n439 585
R3201 VSS.n464 VSS.n463 585
R3202 VSS.n465 VSS.n464 585
R3203 VSS.n470 VSS.n433 585
R3204 VSS.n433 VSS.n432 585
R3205 VSS.n478 VSS.n429 585
R3206 VSS.n429 VSS.n428 585
R3207 VSS.n493 VSS.n492 585
R3208 VSS.n492 VSS.t20 585
R3209 VSS.n505 VSS.n504 585
R3210 VSS.n506 VSS.n505 585
R3211 VSS.n477 VSS.n476 585
R3212 VSS.n476 VSS.n475 585
R3213 VSS.n472 VSS.n471 585
R3214 VSS.n473 VSS.n472 585
R3215 VSS.n462 VSS.n436 585
R3216 VSS.n466 VSS.n436 585
R3217 VSS.n427 VSS.n426 585
R3218 VSS.n491 VSS.n427 585
R3219 VSS.n418 VSS.n417 585
R3220 VSS.n507 VSS.n418 585
R3221 VSS.n377 VSS.n376 585
R3222 VSS.n376 VSS.n375 585
R3223 VSS.n515 VSS.n512 585
R3224 VSS.n734 VSS.n512 585
R3225 VSS.n569 VSS.n565 585
R3226 VSS.n573 VSS.n565 585
R3227 VSS.n584 VSS.n583 585
R3228 VSS.n585 VSS.n584 585
R3229 VSS.n696 VSS.n695 585
R3230 VSS.n697 VSS.n696 585
R3231 VSS.n645 VSS.n643 585
R3232 VSS.t6 VSS.n643 585
R3233 VSS.n659 VSS.n658 585
R3234 VSS.n660 VSS.n659 585
R3235 VSS.n657 VSS.n640 585
R3236 VSS.n661 VSS.n640 585
R3237 VSS.n655 VSS.n623 585
R3238 VSS.n655 VSS.n654 585
R3239 VSS.n694 VSS.n588 585
R3240 VSS.n588 VSS.n587 585
R3241 VSS.n571 VSS.n570 585
R3242 VSS.n572 VSS.n571 585
R3243 VSS.n576 VSS.n547 585
R3244 VSS.n576 VSS.n564 585
R3245 VSS.n662 VSS.n641 585
R3246 VSS.n509 VSS.n508 585
R3247 VSS.n732 VSS.n731 585
R3248 VSS.n733 VSS.n732 585
R3249 VSS.n1033 VSS.n1032 585
R3250 VSS.n1032 VSS.n1031 585
R3251 VSS.n1056 VSS.n1055 585
R3252 VSS.n1057 VSS.n1056 585
R3253 VSS.n1062 VSS.n1025 585
R3254 VSS.n1025 VSS.n1024 585
R3255 VSS.n1070 VSS.n1021 585
R3256 VSS.n1021 VSS.n1020 585
R3257 VSS.n1085 VSS.n1084 585
R3258 VSS.n1084 VSS.t76 585
R3259 VSS.n1097 VSS.n1096 585
R3260 VSS.n1098 VSS.n1097 585
R3261 VSS.n1069 VSS.n1068 585
R3262 VSS.n1068 VSS.n1067 585
R3263 VSS.n1064 VSS.n1063 585
R3264 VSS.n1065 VSS.n1064 585
R3265 VSS.n1054 VSS.n1028 585
R3266 VSS.n1058 VSS.n1028 585
R3267 VSS.n1019 VSS.n1018 585
R3268 VSS.n1083 VSS.n1019 585
R3269 VSS.n1010 VSS.n1009 585
R3270 VSS.n1099 VSS.n1010 585
R3271 VSS.n791 VSS.n790 585
R3272 VSS.n790 VSS.n789 585
R3273 VSS.n1107 VSS.n1104 585
R3274 VSS.n1307 VSS.n1104 585
R3275 VSS.n1161 VSS.n1157 585
R3276 VSS.n1165 VSS.n1157 585
R3277 VSS.n1176 VSS.n1175 585
R3278 VSS.n1177 VSS.n1176 585
R3279 VSS.n1269 VSS.n1268 585
R3280 VSS.n1270 VSS.n1269 585
R3281 VSS.n1230 VSS.n1229 585
R3282 VSS.t67 VSS.n1230 585
R3283 VSS.n1219 VSS.n1217 585
R3284 VSS.n1232 VSS.n1219 585
R3285 VSS.n1216 VSS.n7 585
R3286 VSS.n9 VSS.n7 585
R3287 VSS.n1218 VSS.n1215 585
R3288 VSS.n1231 VSS.n1218 585
R3289 VSS.n1267 VSS.n1180 585
R3290 VSS.n1180 VSS.n1179 585
R3291 VSS.n1163 VSS.n1162 585
R3292 VSS.n1164 VSS.n1163 585
R3293 VSS.n1168 VSS.n1139 585
R3294 VSS.n1168 VSS.n1156 585
R3295 VSS.n2189 VSS.n8 585
R3296 VSS.n1101 VSS.n1100 585
R3297 VSS.n1305 VSS.n1304 585
R3298 VSS.n1306 VSS.n1305 585
R3299 VSS.n166 VSS.n155 585
R3300 VSS.n168 VSS.n155 585
R3301 VSS.n154 VSS.n153 585
R3302 VSS.n1955 VSS.n154 585
R3303 VSS.n1975 VSS.n1974 585
R3304 VSS.n1976 VSS.n1975 585
R3305 VSS.n121 VSS.n120 585
R3306 VSS.n120 VSS.n119 585
R3307 VSS.n2010 VSS.n2009 585
R3308 VSS.n2009 VSS.t39 585
R3309 VSS.n2028 VSS.n2027 585
R3310 VSS.n2029 VSS.n2028 585
R3311 VSS.n139 VSS.n137 585
R3312 VSS.n1978 VSS.n139 585
R3313 VSS.n138 VSS.n136 585
R3314 VSS.n1977 VSS.n138 585
R3315 VSS.n1958 VSS.n1957 585
R3316 VSS.n1957 VSS.n1956 585
R3317 VSS.n118 VSS.n117 585
R3318 VSS.n2008 VSS.n118 585
R3319 VSS.n103 VSS.n102 585
R3320 VSS.n2030 VSS.n103 585
R3321 VSS.n171 VSS.n170 585
R3322 VSS.n170 VSS.n169 585
R3323 VSS.n2139 VSS.n2138 585
R3324 VSS.n2140 VSS.n2139 585
R3325 VSS.n2098 VSS.n2097 585
R3326 VSS.n2099 VSS.n2098 585
R3327 VSS.n72 VSS.n65 585
R3328 VSS.n2100 VSS.n72 585
R3329 VSS.n85 VSS.n84 585
R3330 VSS.n2076 VSS.n85 585
R3331 VSS.n2032 VSS.n2031 585
R3332 VSS.n2039 VSS.n2038 585
R3333 VSS.n2040 VSS.n2039 585
R3334 VSS.n88 VSS.n87 585
R3335 VSS.n87 VSS.n86 585
R3336 VSS.n2079 VSS.n2078 585
R3337 VSS.n2078 VSS.n2077 585
R3338 VSS.n2133 VSS.n44 585
R3339 VSS.n2137 VSS.n44 585
R3340 VSS.n2135 VSS.n2134 585
R3341 VSS.n2136 VSS.n2135 585
R3342 VSS.n45 VSS.n39 585
R3343 VSS.t42 VSS.n45 585
R3344 VSS.n2177 VSS.n17 585
R3345 VSS.n2181 VSS.n17 585
R3346 VSS.n2179 VSS.n2178 585
R3347 VSS.n2180 VSS.n2179 585
R3348 VSS.n14 VSS.n13 585
R3349 VSS.n241 VSS.n230 585
R3350 VSS.n1824 VSS.n230 585
R3351 VSS.n229 VSS.n228 585
R3352 VSS.n1850 VSS.n229 585
R3353 VSS.n1870 VSS.n1869 585
R3354 VSS.n1871 VSS.n1870 585
R3355 VSS.n196 VSS.n195 585
R3356 VSS.n195 VSS.n194 585
R3357 VSS.n1906 VSS.n1905 585
R3358 VSS.n1905 VSS.n1904 585
R3359 VSS.n1924 VSS.n1923 585
R3360 VSS.n1925 VSS.n1924 585
R3361 VSS.n216 VSS.n214 585
R3362 VSS.n1873 VSS.n216 585
R3363 VSS.n215 VSS.n213 585
R3364 VSS.n1872 VSS.n215 585
R3365 VSS.n1853 VSS.n1852 585
R3366 VSS.n1852 VSS.n1851 585
R3367 VSS.n193 VSS.n192 585
R3368 VSS.n1903 VSS.n193 585
R3369 VSS.n178 VSS.n177 585
R3370 VSS.n1926 VSS.n178 585
R3371 VSS.n1827 VSS.n1826 585
R3372 VSS.n1826 VSS.n1825 585
R3373 VSS.n309 VSS.n308 585
R3374 VSS.n308 VSS.n307 585
R3375 VSS.n330 VSS.n329 585
R3376 VSS.n331 VSS.n330 585
R3377 VSS.n336 VSS.n301 585
R3378 VSS.n301 VSS.n300 585
R3379 VSS.n344 VSS.n296 585
R3380 VSS.n296 VSS.n295 585
R3381 VSS.n360 VSS.n359 585
R3382 VSS.n359 VSS.n358 585
R3383 VSS.n372 VSS.n371 585
R3384 VSS.n373 VSS.n372 585
R3385 VSS.n343 VSS.n342 585
R3386 VSS.n342 VSS.n341 585
R3387 VSS.n338 VSS.n337 585
R3388 VSS.n339 VSS.n338 585
R3389 VSS.n328 VSS.n304 585
R3390 VSS.n332 VSS.n304 585
R3391 VSS.n294 VSS.n293 585
R3392 VSS.n357 VSS.n294 585
R3393 VSS.n285 VSS.n284 585
R3394 VSS.n374 VSS.n285 585
R3395 VSS.n244 VSS.n243 585
R3396 VSS.n243 VSS.n242 585
R3397 VSS.n867 VSS.n866 585
R3398 VSS.n869 VSS.n867 585
R3399 VSS.n895 VSS.n894 585
R3400 VSS.n896 VSS.n895 585
R3401 VSS.n852 VSS.n850 585
R3402 VSS.n900 VSS.n852 585
R3403 VSS.n822 VSS.n820 585
R3404 VSS.n931 VSS.n822 585
R3405 VSS.n800 VSS.n799 585
R3406 VSS.n932 VSS.n799 585
R3407 VSS.n808 VSS.n798 585
R3408 VSS.n963 VSS.n798 585
R3409 VSS.n929 VSS.n928 585
R3410 VSS.n930 VSS.n929 585
R3411 VSS.n898 VSS.n832 585
R3412 VSS.n899 VSS.n898 585
R3413 VSS.n893 VSS.n851 585
R3414 VSS.n897 VSS.n851 585
R3415 VSS.n829 VSS.n828 585
R3416 VSS.n933 VSS.n829 585
R3417 VSS.n965 VSS.n797 585
R3418 VSS.n965 VSS.n964 585
R3419 VSS.n872 VSS.n871 585
R3420 VSS.n871 VSS.n870 585
R3421 VSS.n1426 VSS.n1425 585
R3422 VSS.n1425 VSS.n1424 585
R3423 VSS.n1449 VSS.n1448 585
R3424 VSS.n1450 VSS.n1449 585
R3425 VSS.n1455 VSS.n1418 585
R3426 VSS.n1418 VSS.n1417 585
R3427 VSS.n1463 VSS.n1414 585
R3428 VSS.n1414 VSS.n1413 585
R3429 VSS.n1478 VSS.n1477 585
R3430 VSS.n1477 VSS.t73 585
R3431 VSS.n1490 VSS.n1489 585
R3432 VSS.n1491 VSS.n1490 585
R3433 VSS.n1462 VSS.n1461 585
R3434 VSS.n1461 VSS.n1460 585
R3435 VSS.n1457 VSS.n1456 585
R3436 VSS.n1458 VSS.n1457 585
R3437 VSS.n1447 VSS.n1421 585
R3438 VSS.n1451 VSS.n1421 585
R3439 VSS.n1412 VSS.n1411 585
R3440 VSS.n1476 VSS.n1412 585
R3441 VSS.n1403 VSS.n1402 585
R3442 VSS.n1492 VSS.n1403 585
R3443 VSS.n1363 VSS.n1362 585
R3444 VSS.n1362 VSS.n1361 585
R3445 VSS.n1500 VSS.n1497 585
R3446 VSS.n1718 VSS.n1497 585
R3447 VSS.n1527 VSS.n1526 585
R3448 VSS.n1702 VSS.n1527 585
R3449 VSS.n1689 VSS.n1688 585
R3450 VSS.n1688 VSS.n1687 585
R3451 VSS.n1610 VSS.n1609 585
R3452 VSS.n1611 VSS.n1610 585
R3453 VSS.n1618 VSS.n1617 585
R3454 VSS.t13 VSS.n1618 585
R3455 VSS.n1599 VSS.n1597 585
R3456 VSS.n1651 VSS.n1599 585
R3457 VSS.n1649 VSS.n1648 585
R3458 VSS.n1650 VSS.n1649 585
R3459 VSS.n1616 VSS.n1598 585
R3460 VSS.n1619 VSS.n1598 585
R3461 VSS.n1613 VSS.n1580 585
R3462 VSS.n1613 VSS.n1612 585
R3463 VSS.n1705 VSS.n1704 585
R3464 VSS.n1704 VSS.n1703 585
R3465 VSS.n1690 VSS.n1529 585
R3466 VSS.n1529 VSS.n1528 585
R3467 VSS.n1627 VSS.n1626 585
R3468 VSS.n1494 VSS.n1493 585
R3469 VSS.n1716 VSS.n1715 585
R3470 VSS.n1717 VSS.n1716 585
R3471 VSS.n1719 VSS.n1718 403.461
R3472 VSS.n1701 VSS.n1528 403.461
R3473 VSS.n1612 VSS.n1600 403.461
R3474 VSS.n1652 VSS.n1619 403.461
R3475 VSS.n1650 VSS.n1620 403.461
R3476 VSS.n1452 VSS.n1451 396.599
R3477 VSS.n1459 VSS.n1458 396.599
R3478 VSS.n1460 VSS.n1459 396.599
R3479 VSS.n1476 VSS.n1475 396.599
R3480 VSS.n1491 VSS.n1404 396.599
R3481 VSS.n1686 VSS.n1685 395.849
R3482 VSS.n1685 VSS.n1546 395.849
R3483 VSS.n735 VSS.n734 338.954
R3484 VSS.n574 VSS.n564 338.954
R3485 VSS.n653 VSS.n587 338.954
R3486 VSS.n654 VSS.n642 338.954
R3487 VSS.n663 VSS.n661 338.954
R3488 VSS.n1308 VSS.n1307 338.954
R3489 VSS.n1166 VSS.n1156 338.954
R3490 VSS.n1220 VSS.n1179 338.954
R3491 VSS.n1233 VSS.n1231 338.954
R3492 VSS.n2190 VSS.n9 338.954
R3493 VSS.n2041 VSS.n2040 338.954
R3494 VSS.n2099 VSS.n74 338.954
R3495 VSS.n2141 VSS.n2137 338.954
R3496 VSS.n2140 VSS.n18 338.954
R3497 VSS.n2182 VSS.n2181 338.954
R3498 VSS.n699 VSS.n586 332.558
R3499 VSS.n699 VSS.n698 332.558
R3500 VSS.n1272 VSS.n1178 332.558
R3501 VSS.n1272 VSS.n1271 332.558
R3502 VSS.n2102 VSS.n2101 332.558
R3503 VSS.n2101 VSS.n46 332.558
R3504 VSS.n467 VSS.n466 329.38
R3505 VSS.n474 VSS.n473 329.38
R3506 VSS.n475 VSS.n474 329.38
R3507 VSS.n491 VSS.n490 329.38
R3508 VSS.n506 VSS.n419 329.38
R3509 VSS.n1059 VSS.n1058 329.38
R3510 VSS.n1066 VSS.n1065 329.38
R3511 VSS.n1067 VSS.n1066 329.38
R3512 VSS.n1083 VSS.n1082 329.38
R3513 VSS.n1098 VSS.n1011 329.38
R3514 VSS.n1956 VSS.n140 329.38
R3515 VSS.n1979 VSS.n1977 329.38
R3516 VSS.n1979 VSS.n1978 329.38
R3517 VSS.n2008 VSS.n2007 329.38
R3518 VSS.n2029 VSS.n104 329.38
R3519 VSS.n1851 VSS.n217 329.38
R3520 VSS.n1874 VSS.n1872 329.38
R3521 VSS.n1874 VSS.n1873 329.38
R3522 VSS.n1903 VSS.n1902 329.38
R3523 VSS.n1925 VSS.n179 329.38
R3524 VSS.n333 VSS.n332 329.38
R3525 VSS.n340 VSS.n339 329.38
R3526 VSS.n341 VSS.n340 329.38
R3527 VSS.n357 VSS.n356 329.38
R3528 VSS.n373 VSS.n286 329.38
R3529 VSS.t24 VSS.n1498 304.498
R3530 VSS.n701 VSS.n700 292.5
R3531 VSS.n700 VSS.n699 292.5
R3532 VSS.n1274 VSS.n1273 292.5
R3533 VSS.n1273 VSS.n1272 292.5
R3534 VSS.n73 VSS.n57 292.5
R3535 VSS.n2101 VSS.n73 292.5
R3536 VSS.n1684 VSS.n1683 292.5
R3537 VSS.n1685 VSS.n1684 292.5
R3538 VSS.n738 VSS.n737 290.906
R3539 VSS.n665 VSS.n639 290.906
R3540 VSS.n1311 VSS.n1310 290.906
R3541 VSS.n2192 VSS.n6 290.906
R3542 VSS.n2044 VSS.n2043 290.906
R3543 VSS.n2185 VSS.n2184 290.906
R3544 VSS.n1722 VSS.n1721 290.906
R3545 VSS.n1629 VSS.n1628 290.906
R3546 VSS.n1724 VSS.t22 269.807
R3547 VSS.t31 VSS.n513 255.815
R3548 VSS.t27 VSS.n1105 255.815
R3549 VSS.t53 VSS.n2075 255.815
R3550 VSS.t46 VSS.n1422 239.457
R3551 VSS.n2187 VSS.t34 223.941
R3552 VSS.t50 VSS.n437 198.87
R3553 VSS.t58 VSS.n1029 198.87
R3554 VSS.n1954 VSS.t37 198.87
R3555 VSS.n1849 VSS.t1 192.655
R3556 VSS.t10 VSS.n305 192.655
R3557 VSS.n740 VSS.t33 188.758
R3558 VSS.n1313 VSS.t29 188.758
R3559 VSS.n2046 VSS.t55 188.758
R3560 VSS.n1424 VSS.t46 157.143
R3561 VSS.t34 VSS.t8 137.948
R3562 VSS.n1824 VSS.t1 136.724
R3563 VSS.n307 VSS.t10 136.724
R3564 VSS.t3 VSS.t35 130.782
R3565 VSS.n439 VSS.t50 130.508
R3566 VSS.n1031 VSS.t58 130.508
R3567 VSS.n168 VSS.t37 130.508
R3568 VSS.t8 VSS.t3 128.99
R3569 VSS.n901 VSS.n897 128.415
R3570 VSS.n899 VSS.n830 128.415
R3571 VSS.n930 VSS.n830 128.415
R3572 VSS.n934 VSS.n933 128.415
R3573 VSS.n963 VSS.n962 128.415
R3574 VSS.n1687 VSS.n1686 121.799
R3575 VSS.n1611 VSS.n1546 121.799
R3576 VSS.n1458 VSS.n1417 112.246
R3577 VSS.n1460 VSS.n1413 112.246
R3578 VSS.n1702 VSS.n1701 106.575
R3579 VSS.t13 VSS.n1600 106.575
R3580 VSS.n586 VSS.n585 102.326
R3581 VSS.n698 VSS.n697 102.326
R3582 VSS.n1178 VSS.n1177 102.326
R3583 VSS.n1271 VSS.n1270 102.326
R3584 VSS.n2102 VSS.n2100 102.326
R3585 VSS.n2136 VSS.n46 102.326
R3586 VSS.n1703 VSS.t24 98.9624
R3587 VSS.n1451 VSS.n1450 97.2794
R3588 VSS.t73 VSS.n1476 97.2794
R3589 VSS.n473 VSS.n432 93.2208
R3590 VSS.n475 VSS.n428 93.2208
R3591 VSS.n1065 VSS.n1024 93.2208
R3592 VSS.n1067 VSS.n1020 93.2208
R3593 VSS.n1977 VSS.n1976 93.2208
R3594 VSS.n1978 VSS.n119 93.2208
R3595 VSS.n1872 VSS.n1871 93.2208
R3596 VSS.n1873 VSS.n194 93.2208
R3597 VSS.n339 VSS.n300 93.2208
R3598 VSS.n341 VSS.n295 93.2208
R3599 VSS.n1717 VSS.n1498 91.35
R3600 VSS.n1652 VSS.n1651 91.35
R3601 VSS.n574 VSS.n573 89.5354
R3602 VSS.t6 VSS.n653 89.5354
R3603 VSS.n1166 VSS.n1165 89.5354
R3604 VSS.t67 VSS.n1220 89.5354
R3605 VSS.n2077 VSS.n74 89.5354
R3606 VSS.n2141 VSS.t42 89.5354
R3607 VSS.n572 VSS.t31 83.14
R3608 VSS.n1164 VSS.t27 83.14
R3609 VSS.n2076 VSS.t53 83.14
R3610 VSS.n1424 VSS.n1361 82.3134
R3611 VSS.n1492 VSS.n1491 82.3134
R3612 VSS.n736 VSS.n512 81.5708
R3613 VSS.n571 VSS.n514 81.5708
R3614 VSS.n576 VSS.n575 81.5708
R3615 VSS.n652 VSS.n588 81.5708
R3616 VSS.n656 VSS.n655 81.5708
R3617 VSS.n664 VSS.n640 81.5708
R3618 VSS.n1309 VSS.n1104 81.5708
R3619 VSS.n1163 VSS.n1106 81.5708
R3620 VSS.n1168 VSS.n1167 81.5708
R3621 VSS.n1221 VSS.n1180 81.5708
R3622 VSS.n1234 VSS.n1218 81.5708
R3623 VSS.n2191 VSS.n7 81.5708
R3624 VSS.n2042 VSS.n2039 81.5708
R3625 VSS.n2074 VSS.n85 81.5708
R3626 VSS.n2098 VSS.n75 81.5708
R3627 VSS.n2142 VSS.n44 81.5708
R3628 VSS.n2139 VSS.n19 81.5708
R3629 VSS.n2183 VSS.n17 81.5708
R3630 VSS.n1720 VSS.n1497 81.5708
R3631 VSS.n1704 VSS.n1499 81.5708
R3632 VSS.n1700 VSS.n1529 81.5708
R3633 VSS.n1614 VSS.n1613 81.5708
R3634 VSS.n1653 VSS.n1598 81.5708
R3635 VSS.n1649 VSS.n1621 81.5708
R3636 VSS.n466 VSS.n465 80.7915
R3637 VSS.t20 VSS.n491 80.7915
R3638 VSS.n1058 VSS.n1057 80.7915
R3639 VSS.t76 VSS.n1083 80.7915
R3640 VSS.n1956 VSS.n1955 80.7915
R3641 VSS.t39 VSS.n2008 80.7915
R3642 VSS.n1851 VSS.n1850 80.7915
R3643 VSS.n1904 VSS.n1903 80.7915
R3644 VSS.n332 VSS.n331 80.7915
R3645 VSS.n358 VSS.n357 80.7915
R3646 VSS.n700 VSS.n562 80.0317
R3647 VSS.n700 VSS.n563 80.0317
R3648 VSS.n1273 VSS.n1154 80.0317
R3649 VSS.n1273 VSS.n1155 80.0317
R3650 VSS.n2103 VSS.n73 80.0317
R3651 VSS.n73 VSS.n47 80.0317
R3652 VSS.n1684 VSS.n1545 80.0317
R3653 VSS.n1684 VSS.n1547 80.0317
R3654 VSS.n733 VSS.n513 76.7447
R3655 VSS.n660 VSS.n642 76.7447
R3656 VSS.n1306 VSS.n1105 76.7447
R3657 VSS.n1233 VSS.n1232 76.7447
R3658 VSS.n2075 VSS.n86 76.7447
R3659 VSS.n2180 VSS.n18 76.7447
R3660 VSS.n1719 VSS.n1493 76.1251
R3661 VSS.n1626 VSS.n1620 76.1251
R3662 VSS.t62 VSS.n853 75.1106
R3663 VSS.n1425 VSS.n1423 74.5791
R3664 VSS.n1453 VSS.n1421 74.5791
R3665 VSS.n1457 VSS.n1416 74.5791
R3666 VSS.n1461 VSS.n1416 74.5791
R3667 VSS.n1474 VSS.n1412 74.5791
R3668 VSS.n1490 VSS.n1405 74.5791
R3669 VSS.n867 VSS.n854 74.5791
R3670 VSS.n902 VSS.n851 74.5791
R3671 VSS.n898 VSS.n831 74.5791
R3672 VSS.n929 VSS.n831 74.5791
R3673 VSS.n935 VSS.n829 74.5791
R3674 VSS.n961 VSS.n798 74.5791
R3675 VSS.n308 VSS.n306 74.5791
R3676 VSS.n334 VSS.n304 74.5791
R3677 VSS.n338 VSS.n299 74.5791
R3678 VSS.n342 VSS.n299 74.5791
R3679 VSS.n355 VSS.n294 74.5791
R3680 VSS.n372 VSS.n287 74.5791
R3681 VSS.n1848 VSS.n230 74.5791
R3682 VSS.n1852 VSS.n218 74.5791
R3683 VSS.n1875 VSS.n215 74.5791
R3684 VSS.n1875 VSS.n216 74.5791
R3685 VSS.n1901 VSS.n193 74.5791
R3686 VSS.n1924 VSS.n180 74.5791
R3687 VSS.n440 VSS.n438 74.5791
R3688 VSS.n468 VSS.n436 74.5791
R3689 VSS.n472 VSS.n431 74.5791
R3690 VSS.n476 VSS.n431 74.5791
R3691 VSS.n489 VSS.n427 74.5791
R3692 VSS.n505 VSS.n420 74.5791
R3693 VSS.n1032 VSS.n1030 74.5791
R3694 VSS.n1060 VSS.n1028 74.5791
R3695 VSS.n1064 VSS.n1023 74.5791
R3696 VSS.n1068 VSS.n1023 74.5791
R3697 VSS.n1081 VSS.n1019 74.5791
R3698 VSS.n1097 VSS.n1012 74.5791
R3699 VSS.n1953 VSS.n155 74.5791
R3700 VSS.n1957 VSS.n141 74.5791
R3701 VSS.n1980 VSS.n138 74.5791
R3702 VSS.n1980 VSS.n139 74.5791
R3703 VSS.n2006 VSS.n118 74.5791
R3704 VSS.n2028 VSS.n105 74.5791
R3705 VSS.n439 VSS.n375 68.3621
R3706 VSS.n507 VSS.n506 68.3621
R3707 VSS.n1031 VSS.n789 68.3621
R3708 VSS.n1099 VSS.n1098 68.3621
R3709 VSS.n169 VSS.n168 68.3621
R3710 VSS.n2030 VSS.n2029 68.3621
R3711 VSS.n1825 VSS.n1824 68.3621
R3712 VSS.n1926 VSS.n1925 68.3621
R3713 VSS.n307 VSS.n242 68.3621
R3714 VSS.n374 VSS.n373 68.3621
R3715 VSS.n735 VSS.n508 63.954
R3716 VSS.n663 VSS.n662 63.954
R3717 VSS.n1308 VSS.n1100 63.954
R3718 VSS.n2190 VSS.n2189 63.954
R3719 VSS.n2041 VSS.n2031 63.954
R3720 VSS.n2182 VSS.n13 63.954
R3721 VSS.n869 VSS.t62 53.3045
R3722 VSS.n1723 VSS.n1493 53.2877
R3723 VSS.n1626 VSS.n10 53.2877
R3724 VSS.n176 VSS.t71 46.866
R3725 VSS.n282 VSS.t45 46.866
R3726 VSS.n796 VSS.t17 46.866
R3727 VSS.n1400 VSS.t74 46.863
R3728 VSS.n415 VSS.t21 46.863
R3729 VSS.n1007 VSS.t77 46.863
R3730 VSS.n101 VSS.t40 46.863
R3731 VSS.n1371 VSS.t47 46.8459
R3732 VSS.n386 VSS.t51 46.8459
R3733 VSS.n978 VSS.t59 46.8459
R3734 VSS.n151 VSS.t38 46.8459
R3735 VSS.n227 VSS.t2 46.8455
R3736 VSS.n252 VSS.t11 46.8455
R3737 VSS.n858 VSS.t63 46.8455
R3738 VSS.n629 VSS.t7 46.8085
R3739 VSS.n1240 VSS.t68 46.8085
R3740 VSS.n2164 VSS.t43 46.8085
R3741 VSS.n1636 VSS.t14 46.8085
R3742 VSS.n710 VSS.t32 46.808
R3743 VSS.n1283 VSS.t28 46.808
R3744 VSS.n63 VSS.t54 46.808
R3745 VSS.n1543 VSS.t25 46.808
R3746 VSS.n1771 VSS.n1361 44.8985
R3747 VSS.n1726 VSS.n1492 44.8985
R3748 VSS.n739 VSS.n508 44.7679
R3749 VSS.n662 VSS.n11 44.7679
R3750 VSS.n1312 VSS.n1100 44.7679
R3751 VSS.n2189 VSS.n2188 44.7679
R3752 VSS.n2045 VSS.n2031 44.7679
R3753 VSS.n2186 VSS.n13 44.7679
R3754 VSS.n1718 VSS.n1717 38.0628
R3755 VSS.n1651 VSS.n1650 38.0628
R3756 VSS.n787 VSS.n375 37.2886
R3757 VSS.n742 VSS.n507 37.2886
R3758 VSS.n1360 VSS.n789 37.2886
R3759 VSS.n1315 VSS.n1099 37.2886
R3760 VSS.n169 VSS.n167 37.2886
R3761 VSS.n2048 VSS.n2030 37.2886
R3762 VSS.n1825 VSS.n1823 37.2886
R3763 VSS.n1927 VSS.n1926 37.2886
R3764 VSS.n1820 VSS.n242 37.2886
R3765 VSS.n1775 VSS.n374 37.2886
R3766 VSS.n900 VSS.n899 36.3441
R3767 VSS.n931 VSS.n930 36.3441
R3768 VSS.n1725 VSS.n1724 33.5883
R3769 VSS.n734 VSS.n733 31.9772
R3770 VSS.n661 VSS.n660 31.9772
R3771 VSS.n1307 VSS.n1306 31.9772
R3772 VSS.n1232 VSS.n9 31.9772
R3773 VSS.n2040 VSS.n86 31.9772
R3774 VSS.n2181 VSS.n2180 31.9772
R3775 VSS.n897 VSS.n896 31.4983
R3776 VSS.n933 VSS.n932 31.4983
R3777 VSS.n1450 VSS.n1422 29.9325
R3778 VSS.t73 VSS.n1404 29.9325
R3779 VSS.n870 VSS.n869 26.6525
R3780 VSS.n964 VSS.n963 26.6525
R3781 VSS.n465 VSS.n437 24.8593
R3782 VSS.t20 VSS.n419 24.8593
R3783 VSS.n1057 VSS.n1029 24.8593
R3784 VSS.t76 VSS.n1011 24.8593
R3785 VSS.n1955 VSS.n1954 24.8593
R3786 VSS.t39 VSS.n104 24.8593
R3787 VSS.n1850 VSS.n1849 24.8593
R3788 VSS.n331 VSS.n305 24.8593
R3789 VSS.n584 VSS.n562 24.6255
R3790 VSS.n696 VSS.n563 24.6255
R3791 VSS.n1176 VSS.n1154 24.6255
R3792 VSS.n1269 VSS.n1155 24.6255
R3793 VSS.n2103 VSS.n72 24.6255
R3794 VSS.n2135 VSS.n47 24.6255
R3795 VSS.n1688 VSS.n1545 24.6255
R3796 VSS.n1610 VSS.n1547 24.6255
R3797 VSS.n1703 VSS.n1702 22.8379
R3798 VSS.n1619 VSS.t13 22.8379
R3799 VSS.n575 VSS.n565 21.5474
R3800 VSS.n652 VSS.n643 21.5474
R3801 VSS.n1167 VSS.n1157 21.5474
R3802 VSS.n1230 VSS.n1221 21.5474
R3803 VSS.n2078 VSS.n75 21.5474
R3804 VSS.n2142 VSS.n45 21.5474
R3805 VSS.n1700 VSS.n1527 21.5474
R3806 VSS.n1618 VSS.n1614 21.5474
R3807 VSS.n1457 VSS.n1418 21.1076
R3808 VSS.n1461 VSS.n1414 21.1076
R3809 VSS.n898 VSS.n852 21.1076
R3810 VSS.n929 VSS.n822 21.1076
R3811 VSS.n338 VSS.n301 21.1076
R3812 VSS.n342 VSS.n296 21.1076
R3813 VSS.n1870 VSS.n215 21.1076
R3814 VSS.n216 VSS.n195 21.1076
R3815 VSS.n472 VSS.n433 21.1076
R3816 VSS.n476 VSS.n429 21.1076
R3817 VSS.n1064 VSS.n1025 21.1076
R3818 VSS.n1068 VSS.n1021 21.1076
R3819 VSS.n1975 VSS.n138 21.1076
R3820 VSS.n139 VSS.n120 21.1076
R3821 VSS.n573 VSS.n572 19.1865
R3822 VSS.n654 VSS.t6 19.1865
R3823 VSS.n1165 VSS.n1164 19.1865
R3824 VSS.n1231 VSS.t67 19.1865
R3825 VSS.n2077 VSS.n2076 19.1865
R3826 VSS.t42 VSS.n2140 19.1865
R3827 VSS.t70 VSS.n179 18.6446
R3828 VSS.t44 VSS.n286 18.6446
R3829 VSS.n732 VSS.n514 18.4693
R3830 VSS.n659 VSS.n656 18.4693
R3831 VSS.n1305 VSS.n1106 18.4693
R3832 VSS.n1234 VSS.n1219 18.4693
R3833 VSS.n2074 VSS.n87 18.4693
R3834 VSS.n2179 VSS.n19 18.4693
R3835 VSS.n1716 VSS.n1499 18.4693
R3836 VSS.n1653 VSS.n1599 18.4693
R3837 VSS.n1449 VSS.n1421 18.2934
R3838 VSS.n1477 VSS.n1412 18.2934
R3839 VSS.n895 VSS.n851 18.2934
R3840 VSS.n829 VSS.n799 18.2934
R3841 VSS.n330 VSS.n304 18.2934
R3842 VSS.n359 VSS.n294 18.2934
R3843 VSS.n1852 VSS.n229 18.2934
R3844 VSS.n1905 VSS.n193 18.2934
R3845 VSS.n464 VSS.n436 18.2934
R3846 VSS.n492 VSS.n427 18.2934
R3847 VSS.n1056 VSS.n1028 18.2934
R3848 VSS.n1084 VSS.n1019 18.2934
R3849 VSS.n1957 VSS.n154 18.2934
R3850 VSS.n2009 VSS.n118 18.2934
R3851 VSS.n1425 VSS.n1362 15.4791
R3852 VSS.n1490 VSS.n1403 15.4791
R3853 VSS.n871 VSS.n867 15.4791
R3854 VSS.n965 VSS.n798 15.4791
R3855 VSS.n308 VSS.n243 15.4791
R3856 VSS.n372 VSS.n285 15.4791
R3857 VSS.n1826 VSS.n230 15.4791
R3858 VSS.n1924 VSS.n178 15.4791
R3859 VSS.n440 VSS.n376 15.4791
R3860 VSS.n505 VSS.n418 15.4791
R3861 VSS.n1032 VSS.n790 15.4791
R3862 VSS.n1097 VSS.n1010 15.4791
R3863 VSS.n170 VSS.n155 15.4791
R3864 VSS.n2028 VSS.n103 15.4791
R3865 VSS.n736 VSS.n509 15.3911
R3866 VSS.n664 VSS.n641 15.3911
R3867 VSS.n1309 VSS.n1101 15.3911
R3868 VSS.n2191 VSS.n8 15.3911
R3869 VSS.n2042 VSS.n2032 15.3911
R3870 VSS.n2183 VSS.n14 15.3911
R3871 VSS.n1720 VSS.n1494 15.3911
R3872 VSS.n1627 VSS.n1621 15.3911
R3873 VSS.n1452 VSS.n1417 14.9665
R3874 VSS.n1475 VSS.n1413 14.9665
R3875 VSS.n870 VSS.n868 14.5379
R3876 VSS.n964 VSS.n788 14.5379
R3877 VSS.n467 VSS.n432 12.4299
R3878 VSS.n490 VSS.n428 12.4299
R3879 VSS.n1059 VSS.n1024 12.4299
R3880 VSS.n1082 VSS.n1020 12.4299
R3881 VSS.n1976 VSS.n140 12.4299
R3882 VSS.n2007 VSS.n119 12.4299
R3883 VSS.n1871 VSS.n217 12.4299
R3884 VSS.n1902 VSS.n194 12.4299
R3885 VSS.n333 VSS.n300 12.4299
R3886 VSS.n356 VSS.n295 12.4299
R3887 VSS.n896 VSS.n853 9.69213
R3888 VSS.n1770 VSS.n1769 9.38145
R3889 VSS.n1819 VSS.n1818 9.38145
R3890 VSS.n786 VSS.n785 9.38145
R3891 VSS.n873 VSS.n865 9.38145
R3892 VSS.n1359 VSS.n1358 9.38145
R3893 VSS.n172 VSS.n165 9.38145
R3894 VSS.n1828 VSS.n240 9.38145
R3895 VSS.n665 VSS.n635 9.30555
R3896 VSS.n737 VSS.n511 9.30555
R3897 VSS.n2192 VSS.n3 9.30555
R3898 VSS.n1310 VSS.n1103 9.30555
R3899 VSS.n2184 VSS.n16 9.30555
R3900 VSS.n2043 VSS.n2036 9.30555
R3901 VSS.n1630 VSS.n1629 9.30555
R3902 VSS.n1721 VSS.n1496 9.30555
R3903 VSS.n1446 VSS.n1445 9.3005
R3904 VSS.n1467 VSS.n1466 9.3005
R3905 VSS.n1407 VSS.n1406 9.3005
R3906 VSS.n1488 VSS.n1487 9.3005
R3907 VSS.n327 VSS.n326 9.3005
R3908 VSS.n348 VSS.n347 9.3005
R3909 VSS.n289 VSS.n288 9.3005
R3910 VSS.n370 VSS.n369 9.3005
R3911 VSS.n712 VSS.n711 9.3005
R3912 VSS.n638 VSS.n637 9.3005
R3913 VSS.n693 VSS.n692 9.3005
R3914 VSS.n605 VSS.n599 9.3005
R3915 VSS.n560 VSS.n558 9.3005
R3916 VSS.n685 VSS.n684 9.3005
R3917 VSS.n683 VSS.n622 9.3005
R3918 VSS.n691 VSS.n590 9.3005
R3919 VSS.n713 VSS.n545 9.3005
R3920 VSS.n579 VSS.n578 9.3005
R3921 VSS.n607 VSS.n606 9.3005
R3922 VSS.n526 VSS.n525 9.3005
R3923 VSS.n567 VSS.n566 9.3005
R3924 VSS.n568 VSS.n542 9.3005
R3925 VSS.n461 VSS.n460 9.3005
R3926 VSS.n482 VSS.n481 9.3005
R3927 VSS.n422 VSS.n421 9.3005
R3928 VSS.n503 VSS.n502 9.3005
R3929 VSS.n488 VSS.n487 9.3005
R3930 VSS.n489 VSS.n488 9.3005
R3931 VSS.n490 VSS.n489 9.3005
R3932 VSS.n469 VSS.n435 9.3005
R3933 VSS.n469 VSS.n468 9.3005
R3934 VSS.n468 VSS.n467 9.3005
R3935 VSS.n454 VSS.n438 9.3005
R3936 VSS.n438 VSS.n437 9.3005
R3937 VSS.n494 VSS.n425 9.3005
R3938 VSS.n494 VSS.n420 9.3005
R3939 VSS.n420 VSS.n419 9.3005
R3940 VSS.n744 VSS.n743 9.3005
R3941 VSS.n743 VSS.n742 9.3005
R3942 VSS.n787 VSS.n786 9.3005
R3943 VSS.n626 VSS.n624 9.3005
R3944 VSS.n656 VSS.n624 9.3005
R3945 VSS.n656 VSS.n642 9.3005
R3946 VSS.n651 VSS.n650 9.3005
R3947 VSS.n652 VSS.n651 9.3005
R3948 VSS.n653 VSS.n652 9.3005
R3949 VSS.n610 VSS.n589 9.3005
R3950 VSS.n589 VSS.n563 9.3005
R3951 VSS.n698 VSS.n563 9.3005
R3952 VSS.n546 VSS.n543 9.3005
R3953 VSS.n575 VSS.n546 9.3005
R3954 VSS.n575 VSS.n574 9.3005
R3955 VSS.n582 VSS.n581 9.3005
R3956 VSS.n582 VSS.n562 9.3005
R3957 VSS.n586 VSS.n562 9.3005
R3958 VSS.n665 VSS.n664 9.3005
R3959 VSS.n664 VSS.n663 9.3005
R3960 VSS.n737 VSS.n736 9.3005
R3961 VSS.n736 VSS.n735 9.3005
R3962 VSS.n730 VSS.n729 9.3005
R3963 VSS.n730 VSS.n514 9.3005
R3964 VSS.n514 VSS.n513 9.3005
R3965 VSS.n849 VSS.n845 9.3005
R3966 VSS.n827 VSS.n826 9.3005
R3967 VSS.n807 VSS.n806 9.3005
R3968 VSS.n810 VSS.n809 9.3005
R3969 VSS.n1285 VSS.n1284 9.3005
R3970 VSS.n5 VSS.n4 9.3005
R3971 VSS.n1266 VSS.n1265 9.3005
R3972 VSS.n1197 VSS.n1191 9.3005
R3973 VSS.n1152 VSS.n1150 9.3005
R3974 VSS.n1258 VSS.n1257 9.3005
R3975 VSS.n1256 VSS.n1214 9.3005
R3976 VSS.n1264 VSS.n1182 9.3005
R3977 VSS.n1286 VSS.n1137 9.3005
R3978 VSS.n1171 VSS.n1170 9.3005
R3979 VSS.n1199 VSS.n1198 9.3005
R3980 VSS.n1118 VSS.n1117 9.3005
R3981 VSS.n1159 VSS.n1158 9.3005
R3982 VSS.n1160 VSS.n1134 9.3005
R3983 VSS.n1053 VSS.n1052 9.3005
R3984 VSS.n1074 VSS.n1073 9.3005
R3985 VSS.n1014 VSS.n1013 9.3005
R3986 VSS.n1095 VSS.n1094 9.3005
R3987 VSS.n1080 VSS.n1079 9.3005
R3988 VSS.n1081 VSS.n1080 9.3005
R3989 VSS.n1082 VSS.n1081 9.3005
R3990 VSS.n1061 VSS.n1027 9.3005
R3991 VSS.n1061 VSS.n1060 9.3005
R3992 VSS.n1060 VSS.n1059 9.3005
R3993 VSS.n1046 VSS.n1030 9.3005
R3994 VSS.n1030 VSS.n1029 9.3005
R3995 VSS.n1086 VSS.n1017 9.3005
R3996 VSS.n1086 VSS.n1012 9.3005
R3997 VSS.n1012 VSS.n1011 9.3005
R3998 VSS.n1317 VSS.n1316 9.3005
R3999 VSS.n1316 VSS.n1315 9.3005
R4000 VSS.n1360 VSS.n1359 9.3005
R4001 VSS.n1237 VSS.n1235 9.3005
R4002 VSS.n1235 VSS.n1234 9.3005
R4003 VSS.n1234 VSS.n1233 9.3005
R4004 VSS.n1228 VSS.n1227 9.3005
R4005 VSS.n1228 VSS.n1221 9.3005
R4006 VSS.n1221 VSS.n1220 9.3005
R4007 VSS.n1202 VSS.n1181 9.3005
R4008 VSS.n1181 VSS.n1155 9.3005
R4009 VSS.n1271 VSS.n1155 9.3005
R4010 VSS.n1138 VSS.n1135 9.3005
R4011 VSS.n1167 VSS.n1138 9.3005
R4012 VSS.n1167 VSS.n1166 9.3005
R4013 VSS.n1174 VSS.n1173 9.3005
R4014 VSS.n1174 VSS.n1154 9.3005
R4015 VSS.n1178 VSS.n1154 9.3005
R4016 VSS.n2192 VSS.n2191 9.3005
R4017 VSS.n2191 VSS.n2190 9.3005
R4018 VSS.n1310 VSS.n1309 9.3005
R4019 VSS.n1309 VSS.n1308 9.3005
R4020 VSS.n1303 VSS.n1302 9.3005
R4021 VSS.n1303 VSS.n1106 9.3005
R4022 VSS.n1106 VSS.n1105 9.3005
R4023 VSS.n1960 VSS.n1959 9.3005
R4024 VSS.n1998 VSS.n1997 9.3005
R4025 VSS.n107 VSS.n106 9.3005
R4026 VSS.n2026 VSS.n2025 9.3005
R4027 VSS.n2005 VSS.n2004 9.3005
R4028 VSS.n2006 VSS.n2005 9.3005
R4029 VSS.n2007 VSS.n2006 9.3005
R4030 VSS.n1973 VSS.n1972 9.3005
R4031 VSS.n1973 VSS.n141 9.3005
R4032 VSS.n141 VSS.n140 9.3005
R4033 VSS.n1953 VSS.n1952 9.3005
R4034 VSS.n1954 VSS.n1953 9.3005
R4035 VSS.n2013 VSS.n2012 9.3005
R4036 VSS.n2012 VSS.n105 9.3005
R4037 VSS.n105 VSS.n104 9.3005
R4038 VSS.n2050 VSS.n2049 9.3005
R4039 VSS.n2049 VSS.n2048 9.3005
R4040 VSS.n167 VSS.n165 9.3005
R4041 VSS.n2176 VSS.n2175 9.3005
R4042 VSS.n2156 VSS.n2155 9.3005
R4043 VSS.n2132 VSS.n36 9.3005
R4044 VSS.n2146 VSS.n37 9.3005
R4045 VSS.n2119 VSS.n2118 9.3005
R4046 VSS.n68 VSS.n67 9.3005
R4047 VSS.n2067 VSS.n2066 9.3005
R4048 VSS.n2043 VSS.n2042 9.3005
R4049 VSS.n2042 VSS.n2041 9.3005
R4050 VSS.n2037 VSS.n96 9.3005
R4051 VSS.n2065 VSS.n83 9.3005
R4052 VSS.n2073 VSS.n2072 9.3005
R4053 VSS.n2074 VSS.n2073 9.3005
R4054 VSS.n2075 VSS.n2074 9.3005
R4055 VSS.n2082 VSS.n2081 9.3005
R4056 VSS.n2081 VSS.n75 9.3005
R4057 VSS.n75 VSS.n74 9.3005
R4058 VSS.n2094 VSS.n76 9.3005
R4059 VSS.n2096 VSS.n2095 9.3005
R4060 VSS.n2105 VSS.n2104 9.3005
R4061 VSS.n2104 VSS.n2103 9.3005
R4062 VSS.n2103 VSS.n2102 9.3005
R4063 VSS.n70 VSS.n69 9.3005
R4064 VSS.n2117 VSS.n56 9.3005
R4065 VSS.n2131 VSS.n2130 9.3005
R4066 VSS.n2131 VSS.n47 9.3005
R4067 VSS.n47 VSS.n46 9.3005
R4068 VSS.n2143 VSS.n43 9.3005
R4069 VSS.n2143 VSS.n2142 9.3005
R4070 VSS.n2142 VSS.n2141 9.3005
R4071 VSS.n2154 VSS.n29 9.3005
R4072 VSS.n26 VSS.n20 9.3005
R4073 VSS.n20 VSS.n19 9.3005
R4074 VSS.n19 VSS.n18 9.3005
R4075 VSS.n2184 VSS.n2183 9.3005
R4076 VSS.n2183 VSS.n2182 9.3005
R4077 VSS.n1855 VSS.n1854 9.3005
R4078 VSS.n1893 VSS.n1892 9.3005
R4079 VSS.n182 VSS.n181 9.3005
R4080 VSS.n1922 VSS.n1921 9.3005
R4081 VSS.n1900 VSS.n1899 9.3005
R4082 VSS.n1901 VSS.n1900 9.3005
R4083 VSS.n1902 VSS.n1901 9.3005
R4084 VSS.n1868 VSS.n1867 9.3005
R4085 VSS.n1868 VSS.n218 9.3005
R4086 VSS.n218 VSS.n217 9.3005
R4087 VSS.n1848 VSS.n1847 9.3005
R4088 VSS.n1849 VSS.n1848 9.3005
R4089 VSS.n1909 VSS.n1908 9.3005
R4090 VSS.n1908 VSS.n180 9.3005
R4091 VSS.n180 VSS.n179 9.3005
R4092 VSS.n1929 VSS.n1928 9.3005
R4093 VSS.n1928 VSS.n1927 9.3005
R4094 VSS.n1823 VSS.n240 9.3005
R4095 VSS.n354 VSS.n353 9.3005
R4096 VSS.n355 VSS.n354 9.3005
R4097 VSS.n356 VSS.n355 9.3005
R4098 VSS.n335 VSS.n303 9.3005
R4099 VSS.n335 VSS.n334 9.3005
R4100 VSS.n334 VSS.n333 9.3005
R4101 VSS.n322 VSS.n306 9.3005
R4102 VSS.n306 VSS.n305 9.3005
R4103 VSS.n361 VSS.n292 9.3005
R4104 VSS.n361 VSS.n287 9.3005
R4105 VSS.n287 VSS.n286 9.3005
R4106 VSS.n1777 VSS.n1776 9.3005
R4107 VSS.n1776 VSS.n1775 9.3005
R4108 VSS.n1820 VSS.n1819 9.3005
R4109 VSS.n937 VSS.n936 9.3005
R4110 VSS.n936 VSS.n935 9.3005
R4111 VSS.n935 VSS.n934 9.3005
R4112 VSS.n903 VSS.n848 9.3005
R4113 VSS.n903 VSS.n902 9.3005
R4114 VSS.n902 VSS.n901 9.3005
R4115 VSS.n892 VSS.n854 9.3005
R4116 VSS.n854 VSS.n853 9.3005
R4117 VSS.n960 VSS.n959 9.3005
R4118 VSS.n961 VSS.n960 9.3005
R4119 VSS.n962 VSS.n961 9.3005
R4120 VSS.n967 VSS.n966 9.3005
R4121 VSS.n966 VSS.n788 9.3005
R4122 VSS.n868 VSS.n865 9.3005
R4123 VSS.n1473 VSS.n1472 9.3005
R4124 VSS.n1474 VSS.n1473 9.3005
R4125 VSS.n1475 VSS.n1474 9.3005
R4126 VSS.n1454 VSS.n1420 9.3005
R4127 VSS.n1454 VSS.n1453 9.3005
R4128 VSS.n1453 VSS.n1452 9.3005
R4129 VSS.n1439 VSS.n1423 9.3005
R4130 VSS.n1423 VSS.n1422 9.3005
R4131 VSS.n1479 VSS.n1410 9.3005
R4132 VSS.n1479 VSS.n1405 9.3005
R4133 VSS.n1405 VSS.n1404 9.3005
R4134 VSS.n1728 VSS.n1727 9.3005
R4135 VSS.n1727 VSS.n1726 9.3005
R4136 VSS.n1771 VSS.n1770 9.3005
R4137 VSS.n1692 VSS.n1691 9.3005
R4138 VSS.n1647 VSS.n1646 9.3005
R4139 VSS.n1673 VSS.n1672 9.3005
R4140 VSS.n1551 VSS.n1549 9.3005
R4141 VSS.n1569 VSS.n1568 9.3005
R4142 VSS.n1654 VSS.n1595 9.3005
R4143 VSS.n1654 VSS.n1653 9.3005
R4144 VSS.n1653 VSS.n1652 9.3005
R4145 VSS.n1615 VSS.n1586 9.3005
R4146 VSS.n1596 VSS.n1594 9.3005
R4147 VSS.n1585 VSS.n1581 9.3005
R4148 VSS.n1614 VSS.n1581 9.3005
R4149 VSS.n1614 VSS.n1600 9.3005
R4150 VSS.n1671 VSS.n1579 9.3005
R4151 VSS.n1608 VSS.n1607 9.3005
R4152 VSS.n1608 VSS.n1547 9.3005
R4153 VSS.n1547 VSS.n1546 9.3005
R4154 VSS.n1699 VSS.n1698 9.3005
R4155 VSS.n1700 VSS.n1699 9.3005
R4156 VSS.n1701 VSS.n1700 9.3005
R4157 VSS.n1693 VSS.n1542 9.3005
R4158 VSS.n1564 VSS.n1544 9.3005
R4159 VSS.n1545 VSS.n1544 9.3005
R4160 VSS.n1686 VSS.n1545 9.3005
R4161 VSS.n1567 VSS.n1556 9.3005
R4162 VSS.n1603 VSS.n1602 9.3005
R4163 VSS.n1629 VSS.n1621 9.3005
R4164 VSS.n1621 VSS.n1620 9.3005
R4165 VSS.n1510 VSS.n1509 9.3005
R4166 VSS.n1721 VSS.n1720 9.3005
R4167 VSS.n1720 VSS.n1719 9.3005
R4168 VSS.n1714 VSS.n1713 9.3005
R4169 VSS.n1714 VSS.n1499 9.3005
R4170 VSS.n1499 VSS.n1498 9.3005
R4171 VSS.n1708 VSS.n1707 9.3005
R4172 VSS.n1706 VSS.n1525 9.3005
R4173 VSS.n431 VSS.n430 9.15497
R4174 VSS.n474 VSS.n431 9.15497
R4175 VSS.n1023 VSS.n1022 9.15497
R4176 VSS.n1066 VSS.n1023 9.15497
R4177 VSS.n1981 VSS.n1980 9.15497
R4178 VSS.n1980 VSS.n1979 9.15497
R4179 VSS.n1876 VSS.n1875 9.15497
R4180 VSS.n1875 VSS.n1874 9.15497
R4181 VSS.n299 VSS.n298 9.15497
R4182 VSS.n340 VSS.n299 9.15497
R4183 VSS.n927 VSS.n831 9.15497
R4184 VSS.n831 VSS.n830 9.15497
R4185 VSS.n1416 VSS.n1415 9.15497
R4186 VSS.n1459 VSS.n1416 9.15497
R4187 VSS.n1770 VSS.n1362 8.44336
R4188 VSS.n1727 VSS.n1403 8.44336
R4189 VSS.n871 VSS.n865 8.44336
R4190 VSS.n966 VSS.n965 8.44336
R4191 VSS.n1819 VSS.n243 8.44336
R4192 VSS.n1776 VSS.n285 8.44336
R4193 VSS.n1826 VSS.n240 8.44336
R4194 VSS.n1928 VSS.n178 8.44336
R4195 VSS.n786 VSS.n376 8.44336
R4196 VSS.n743 VSS.n418 8.44336
R4197 VSS.n1359 VSS.n790 8.44336
R4198 VSS.n1316 VSS.n1010 8.44336
R4199 VSS.n170 VSS.n165 8.44336
R4200 VSS.n2049 VSS.n103 8.44336
R4201 VSS.n732 VSS.n512 7.69581
R4202 VSS.n659 VSS.n640 7.69581
R4203 VSS.n1305 VSS.n1104 7.69581
R4204 VSS.n1219 VSS.n7 7.69581
R4205 VSS.n2039 VSS.n87 7.69581
R4206 VSS.n2179 VSS.n17 7.69581
R4207 VSS.n1716 VSS.n1497 7.69581
R4208 VSS.n1649 VSS.n1599 7.69581
R4209 VSS.n1687 VSS.n1528 7.61296
R4210 VSS.n1612 VSS.n1611 7.61296
R4211 VSS.n962 VSS.t16 7.26922
R4212 VSS.n585 VSS.n564 6.39585
R4213 VSS.n697 VSS.n587 6.39585
R4214 VSS.n1177 VSS.n1156 6.39585
R4215 VSS.n1270 VSS.n1179 6.39585
R4216 VSS.n2100 VSS.n2099 6.39585
R4217 VSS.n2137 VSS.n2136 6.39585
R4218 VSS.n1904 VSS.t70 6.21519
R4219 VSS.n358 VSS.t44 6.21519
R4220 VSS.n1449 VSS.n1423 5.62907
R4221 VSS.n1477 VSS.n1405 5.62907
R4222 VSS.n895 VSS.n854 5.62907
R4223 VSS.n961 VSS.n799 5.62907
R4224 VSS.n330 VSS.n306 5.62907
R4225 VSS.n359 VSS.n287 5.62907
R4226 VSS.n1848 VSS.n229 5.62907
R4227 VSS.n1905 VSS.n180 5.62907
R4228 VSS.n464 VSS.n438 5.62907
R4229 VSS.n492 VSS.n420 5.62907
R4230 VSS.n1056 VSS.n1030 5.62907
R4231 VSS.n1084 VSS.n1012 5.62907
R4232 VSS.n1953 VSS.n154 5.62907
R4233 VSS.n2009 VSS.n105 5.62907
R4234 VSS.n641 VSS.n639 5.33568
R4235 VSS.n738 VSS.n509 5.33568
R4236 VSS.n8 VSS.n6 5.33568
R4237 VSS.n1311 VSS.n1101 5.33568
R4238 VSS.n2044 VSS.n2032 5.33568
R4239 VSS.n2185 VSS.n14 5.33568
R4240 VSS.n1628 VSS.n1627 5.33568
R4241 VSS.n1722 VSS.n1494 5.33568
R4242 VSS.n901 VSS.n900 4.84631
R4243 VSS.n934 VSS.n931 4.84631
R4244 VSS.n1456 VSS.n1415 4.84621
R4245 VSS.n1462 VSS.n1415 4.84621
R4246 VSS.n337 VSS.n298 4.84621
R4247 VSS.n343 VSS.n298 4.84621
R4248 VSS.n471 VSS.n430 4.84621
R4249 VSS.n477 VSS.n430 4.84621
R4250 VSS.n927 VSS.n832 4.84621
R4251 VSS.n928 VSS.n927 4.84621
R4252 VSS.n1063 VSS.n1022 4.84621
R4253 VSS.n1069 VSS.n1022 4.84621
R4254 VSS.n1981 VSS.n136 4.84621
R4255 VSS.n1981 VSS.n137 4.84621
R4256 VSS.n1876 VSS.n213 4.84621
R4257 VSS.n1876 VSS.n214 4.84621
R4258 VSS.n1433 VSS.n1427 4.6505
R4259 VSS.n316 VSS.n310 4.6505
R4260 VSS.n448 VSS.n442 4.6505
R4261 VSS.n877 VSS.n855 4.6505
R4262 VSS.n1040 VSS.n1034 4.6505
R4263 VSS.n1937 VSS.n156 4.6505
R4264 VSS.n1832 VSS.n231 4.6505
R4265 VSS.n571 VSS.n565 4.61769
R4266 VSS.n655 VSS.n643 4.61769
R4267 VSS.n1163 VSS.n1157 4.61769
R4268 VSS.n1230 VSS.n1218 4.61769
R4269 VSS.n2078 VSS.n85 4.61769
R4270 VSS.n2139 VSS.n45 4.61769
R4271 VSS.n1704 VSS.n1527 4.61769
R4272 VSS.n1618 VSS.n1598 4.61769
R4273 VSS.n1483 VSS.n1482 4.5005
R4274 VSS.n1486 VSS.n1485 4.5005
R4275 VSS.n1469 VSS.n1468 4.5005
R4276 VSS.n1444 VSS.n1443 4.5005
R4277 VSS.n1435 VSS.n1434 4.5005
R4278 VSS.n1436 VSS.n1428 4.5005
R4279 VSS.n1432 VSS.n1429 4.5005
R4280 VSS.n1393 VSS.n1391 4.5005
R4281 VSS.n1738 VSS.n1737 4.5005
R4282 VSS.n1745 VSS.n1383 4.5005
R4283 VSS.n1752 VSS.n1751 4.5005
R4284 VSS.n1753 VSS.n1375 4.5005
R4285 VSS.n1440 VSS.n1372 4.5005
R4286 VSS.n1760 VSS.n1759 4.5005
R4287 VSS.n1744 VSS.n1743 4.5005
R4288 VSS.n1484 VSS.n1408 4.5005
R4289 VSS.n1768 VSS.n1767 4.5005
R4290 VSS.n1481 VSS.n1409 4.5005
R4291 VSS.n1481 VSS.n1480 4.5005
R4292 VSS.n1442 VSS.n1441 4.5005
R4293 VSS.n1441 VSS.n1419 4.5005
R4294 VSS.n1438 VSS.n1437 4.5005
R4295 VSS.n1471 VSS.n1470 4.5005
R4296 VSS.n1471 VSS.n1464 4.5005
R4297 VSS.n1730 VSS.n1401 4.5005
R4298 VSS.n1730 VSS.n1729 4.5005
R4299 VSS.n365 VSS.n364 4.5005
R4300 VSS.n368 VSS.n367 4.5005
R4301 VSS.n350 VSS.n349 4.5005
R4302 VSS.n325 VSS.n253 4.5005
R4303 VSS.n318 VSS.n317 4.5005
R4304 VSS.n319 VSS.n311 4.5005
R4305 VSS.n1817 VSS.n1816 4.5005
R4306 VSS.n315 VSS.n312 4.5005
R4307 VSS.n363 VSS.n291 4.5005
R4308 VSS.n363 VSS.n362 4.5005
R4309 VSS.n275 VSS.n273 4.5005
R4310 VSS.n1787 VSS.n1786 4.5005
R4311 VSS.n1794 VSS.n265 4.5005
R4312 VSS.n1801 VSS.n1800 4.5005
R4313 VSS.n297 VSS.n261 4.5005
R4314 VSS.n1802 VSS.n256 4.5005
R4315 VSS.n324 VSS.n323 4.5005
R4316 VSS.n324 VSS.n302 4.5005
R4317 VSS.n1809 VSS.n1808 4.5005
R4318 VSS.n321 VSS.n320 4.5005
R4319 VSS.n1793 VSS.n1792 4.5005
R4320 VSS.n352 VSS.n351 4.5005
R4321 VSS.n352 VSS.n345 4.5005
R4322 VSS.n366 VSS.n290 4.5005
R4323 VSS.n1779 VSS.n283 4.5005
R4324 VSS.n1779 VSS.n1778 4.5005
R4325 VSS.n678 VSS.n677 4.5005
R4326 VSS.n600 VSS.n597 4.5005
R4327 VSS.n717 VSS.n716 4.5005
R4328 VSS.n527 VSS.n510 4.5005
R4329 VSS.n535 VSS.n534 4.5005
R4330 VSS.n728 VSS.n727 4.5005
R4331 VSS.n728 VSS.n516 4.5005
R4332 VSS.n580 VSS.n577 4.5005
R4333 VSS.n720 VSS.n541 4.5005
R4334 VSS.n715 VSS.n544 4.5005
R4335 VSS.n715 VSS.n714 4.5005
R4336 VSS.n636 VSS.n634 4.5005
R4337 VSS.n594 VSS.n592 4.5005
R4338 VSS.n644 VSS.n592 4.5005
R4339 VSS.n621 VSS.n619 4.5005
R4340 VSS.n609 VSS.n598 4.5005
R4341 VSS.n609 VSS.n608 4.5005
R4342 VSS.n614 VSS.n591 4.5005
R4343 VSS.n704 VSS.n703 4.5005
R4344 VSS.n703 VSS.n702 4.5005
R4345 VSS.n676 VSS.n628 4.5005
R4346 VSS.n681 VSS.n680 4.5005
R4347 VSS.n682 VSS.n681 4.5005
R4348 VSS.n604 VSS.n603 4.5005
R4349 VSS.n604 VSS.n561 4.5005
R4350 VSS.n647 VSS.n646 4.5005
R4351 VSS.n667 VSS.n666 4.5005
R4352 VSS.n523 VSS.n517 4.5005
R4353 VSS.n536 VSS.n524 4.5005
R4354 VSS.n498 VSS.n497 4.5005
R4355 VSS.n501 VSS.n500 4.5005
R4356 VSS.n484 VSS.n483 4.5005
R4357 VSS.n459 VSS.n458 4.5005
R4358 VSS.n450 VSS.n449 4.5005
R4359 VSS.n451 VSS.n443 4.5005
R4360 VSS.n447 VSS.n444 4.5005
R4361 VSS.n408 VSS.n406 4.5005
R4362 VSS.n754 VSS.n753 4.5005
R4363 VSS.n761 VSS.n398 4.5005
R4364 VSS.n768 VSS.n767 4.5005
R4365 VSS.n769 VSS.n390 4.5005
R4366 VSS.n455 VSS.n387 4.5005
R4367 VSS.n776 VSS.n775 4.5005
R4368 VSS.n760 VSS.n759 4.5005
R4369 VSS.n499 VSS.n423 4.5005
R4370 VSS.n784 VSS.n783 4.5005
R4371 VSS.n496 VSS.n424 4.5005
R4372 VSS.n496 VSS.n495 4.5005
R4373 VSS.n457 VSS.n456 4.5005
R4374 VSS.n456 VSS.n434 4.5005
R4375 VSS.n453 VSS.n452 4.5005
R4376 VSS.n486 VSS.n485 4.5005
R4377 VSS.n486 VSS.n479 4.5005
R4378 VSS.n746 VSS.n416 4.5005
R4379 VSS.n746 VSS.n745 4.5005
R4380 VSS.n956 VSS.n803 4.5005
R4381 VSS.n955 VSS.n954 4.5005
R4382 VSS.n825 VSS.n824 4.5005
R4383 VSS.n907 VSS.n906 4.5005
R4384 VSS.n880 VSS.n878 4.5005
R4385 VSS.n879 VSS.n856 4.5005
R4386 VSS.n876 VSS.n875 4.5005
R4387 VSS.n882 VSS.n881 4.5005
R4388 VSS.n958 VSS.n957 4.5005
R4389 VSS.n958 VSS.n801 4.5005
R4390 VSS.n814 VSS.n813 4.5005
R4391 VSS.n945 VSS.n944 4.5005
R4392 VSS.n837 VSS.n836 4.5005
R4393 VSS.n916 VSS.n915 4.5005
R4394 VSS.n926 VSS.n834 4.5005
R4395 VSS.n914 VSS.n913 4.5005
R4396 VSS.n905 VSS.n844 4.5005
R4397 VSS.n905 VSS.n904 4.5005
R4398 VSS.n859 VSS.n843 4.5005
R4399 VSS.n891 VSS.n857 4.5005
R4400 VSS.n818 VSS.n816 4.5005
R4401 VSS.n823 VSS.n819 4.5005
R4402 VSS.n821 VSS.n819 4.5005
R4403 VSS.n953 VSS.n805 4.5005
R4404 VSS.n970 VSS.n969 4.5005
R4405 VSS.n969 VSS.n968 4.5005
R4406 VSS.n1251 VSS.n1250 4.5005
R4407 VSS.n1192 VSS.n1189 4.5005
R4408 VSS.n1290 VSS.n1289 4.5005
R4409 VSS.n1119 VSS.n1102 4.5005
R4410 VSS.n1127 VSS.n1126 4.5005
R4411 VSS.n1301 VSS.n1300 4.5005
R4412 VSS.n1301 VSS.n1108 4.5005
R4413 VSS.n1172 VSS.n1169 4.5005
R4414 VSS.n1293 VSS.n1133 4.5005
R4415 VSS.n1288 VSS.n1136 4.5005
R4416 VSS.n1288 VSS.n1287 4.5005
R4417 VSS.n1242 VSS.n1241 4.5005
R4418 VSS.n1186 VSS.n1184 4.5005
R4419 VSS.n1222 VSS.n1184 4.5005
R4420 VSS.n1213 VSS.n1211 4.5005
R4421 VSS.n1201 VSS.n1190 4.5005
R4422 VSS.n1201 VSS.n1200 4.5005
R4423 VSS.n1206 VSS.n1183 4.5005
R4424 VSS.n1277 VSS.n1276 4.5005
R4425 VSS.n1276 VSS.n1275 4.5005
R4426 VSS.n1249 VSS.n1239 4.5005
R4427 VSS.n1254 VSS.n1253 4.5005
R4428 VSS.n1255 VSS.n1254 4.5005
R4429 VSS.n1196 VSS.n1195 4.5005
R4430 VSS.n1196 VSS.n1153 4.5005
R4431 VSS.n1224 VSS.n1223 4.5005
R4432 VSS.n2194 VSS.n2193 4.5005
R4433 VSS.n1115 VSS.n1109 4.5005
R4434 VSS.n1128 VSS.n1116 4.5005
R4435 VSS.n1090 VSS.n1089 4.5005
R4436 VSS.n1093 VSS.n1092 4.5005
R4437 VSS.n1076 VSS.n1075 4.5005
R4438 VSS.n1051 VSS.n1050 4.5005
R4439 VSS.n1042 VSS.n1041 4.5005
R4440 VSS.n1043 VSS.n1035 4.5005
R4441 VSS.n1039 VSS.n1036 4.5005
R4442 VSS.n1000 VSS.n998 4.5005
R4443 VSS.n1327 VSS.n1326 4.5005
R4444 VSS.n1334 VSS.n990 4.5005
R4445 VSS.n1341 VSS.n1340 4.5005
R4446 VSS.n1342 VSS.n982 4.5005
R4447 VSS.n1047 VSS.n979 4.5005
R4448 VSS.n1349 VSS.n1348 4.5005
R4449 VSS.n1333 VSS.n1332 4.5005
R4450 VSS.n1091 VSS.n1015 4.5005
R4451 VSS.n1357 VSS.n1356 4.5005
R4452 VSS.n1088 VSS.n1016 4.5005
R4453 VSS.n1088 VSS.n1087 4.5005
R4454 VSS.n1049 VSS.n1048 4.5005
R4455 VSS.n1048 VSS.n1026 4.5005
R4456 VSS.n1045 VSS.n1044 4.5005
R4457 VSS.n1078 VSS.n1077 4.5005
R4458 VSS.n1078 VSS.n1071 4.5005
R4459 VSS.n1319 VSS.n1008 4.5005
R4460 VSS.n1319 VSS.n1318 4.5005
R4461 VSS.n114 VSS.n109 4.5005
R4462 VSS.n2024 VSS.n2023 4.5005
R4463 VSS.n2001 VSS.n124 4.5005
R4464 VSS.n152 VSS.n150 4.5005
R4465 VSS.n1940 VSS.n1938 4.5005
R4466 VSS.n1939 VSS.n157 4.5005
R4467 VSS.n1942 VSS.n1941 4.5005
R4468 VSS.n2000 VSS.n1999 4.5005
R4469 VSS.n126 VSS.n113 4.5005
R4470 VSS.n1990 VSS.n1989 4.5005
R4471 VSS.n135 VSS.n133 4.5005
R4472 VSS.n147 VSS.n146 4.5005
R4473 VSS.n1962 VSS.n1961 4.5005
R4474 VSS.n159 VSS.n149 4.5005
R4475 VSS.n1991 VSS.n128 4.5005
R4476 VSS.n2022 VSS.n108 4.5005
R4477 VSS.n1936 VSS.n1935 4.5005
R4478 VSS.n116 VSS.n115 4.5005
R4479 VSS.n2011 VSS.n116 4.5005
R4480 VSS.n145 VSS.n143 4.5005
R4481 VSS.n143 VSS.n142 4.5005
R4482 VSS.n1951 VSS.n158 4.5005
R4483 VSS.n2003 VSS.n2002 4.5005
R4484 VSS.n2003 VSS.n122 4.5005
R4485 VSS.n2053 VSS.n2052 4.5005
R4486 VSS.n2052 VSS.n2051 4.5005
R4487 VSS.n2167 VSS.n21 4.5005
R4488 VSS.n2163 VSS.n25 4.5005
R4489 VSS.n53 VSS.n52 4.5005
R4490 VSS.n78 VSS.n77 4.5005
R4491 VSS.n2080 VSS.n77 4.5005
R4492 VSS.n2059 VSS.n2058 4.5005
R4493 VSS.n2035 VSS.n2033 4.5005
R4494 VSS.n2087 VSS.n82 4.5005
R4495 VSS.n2060 VSS.n95 4.5005
R4496 VSS.n2070 VSS.n91 4.5005
R4497 VSS.n91 VSS.n89 4.5005
R4498 VSS.n71 VSS.n64 4.5005
R4499 VSS.n2112 VSS.n58 4.5005
R4500 VSS.n66 VSS.n58 4.5005
R4501 VSS.n2115 VSS.n55 4.5005
R4502 VSS.n2116 VSS.n2115 4.5005
R4503 VSS.n51 VSS.n49 4.5005
R4504 VSS.n49 VSS.n48 4.5005
R4505 VSS.n2145 VSS.n35 4.5005
R4506 VSS.n2145 VSS.n2144 4.5005
R4507 VSS.n31 VSS.n30 4.5005
R4508 VSS.n2159 VSS.n2158 4.5005
R4509 VSS.n2158 VSS.n2157 4.5005
R4510 VSS.n22 VSS.n15 4.5005
R4511 VSS.n40 VSS.n38 4.5005
R4512 VSS.n92 VSS.n90 4.5005
R4513 VSS.n2162 VSS.n2161 4.5005
R4514 VSS.n2121 VSS.n2120 4.5005
R4515 VSS.n2084 VSS.n2083 4.5005
R4516 VSS.n189 VSS.n184 4.5005
R4517 VSS.n1920 VSS.n1919 4.5005
R4518 VSS.n1896 VSS.n199 4.5005
R4519 VSS.n1857 VSS.n1856 4.5005
R4520 VSS.n1835 VSS.n1833 4.5005
R4521 VSS.n1834 VSS.n232 4.5005
R4522 VSS.n1837 VSS.n1836 4.5005
R4523 VSS.n1895 VSS.n1894 4.5005
R4524 VSS.n201 VSS.n188 4.5005
R4525 VSS.n1885 VSS.n1884 4.5005
R4526 VSS.n210 VSS.n208 4.5005
R4527 VSS.n224 VSS.n223 4.5005
R4528 VSS.n234 VSS.n226 4.5005
R4529 VSS.n1886 VSS.n203 4.5005
R4530 VSS.n1918 VSS.n183 4.5005
R4531 VSS.n1831 VSS.n1830 4.5005
R4532 VSS.n191 VSS.n190 4.5005
R4533 VSS.n1907 VSS.n191 4.5005
R4534 VSS.n1877 VSS.n209 4.5005
R4535 VSS.n222 VSS.n220 4.5005
R4536 VSS.n220 VSS.n219 4.5005
R4537 VSS.n1846 VSS.n233 4.5005
R4538 VSS.n1898 VSS.n1897 4.5005
R4539 VSS.n1898 VSS.n197 4.5005
R4540 VSS.n1932 VSS.n1931 4.5005
R4541 VSS.n1931 VSS.n1930 4.5005
R4542 VSS.n1634 VSS.n1633 4.5005
R4543 VSS.n1604 VSS.n1553 4.5005
R4544 VSS.n1697 VSS.n1696 4.5005
R4545 VSS.n1511 VSS.n1495 4.5005
R4546 VSS.n1519 VSS.n1518 4.5005
R4547 VSS.n1711 VSS.n1503 4.5005
R4548 VSS.n1503 VSS.n1501 4.5005
R4549 VSS.n1566 VSS.n1565 4.5005
R4550 VSS.n1537 VSS.n1536 4.5005
R4551 VSS.n1695 VSS.n1532 4.5005
R4552 VSS.n1532 VSS.n1530 4.5005
R4553 VSS.n1639 VSS.n1623 4.5005
R4554 VSS.n1669 VSS.n1668 4.5005
R4555 VSS.n1670 VSS.n1669 4.5005
R4556 VSS.n1664 VSS.n1584 4.5005
R4557 VSS.n1606 VSS.n1605 4.5005
R4558 VSS.n1606 VSS.n1601 4.5005
R4559 VSS.n1674 VSS.n1577 4.5005
R4560 VSS.n1571 VSS.n1570 4.5005
R4561 VSS.n1570 VSS.n1548 4.5005
R4562 VSS.n1635 VSS.n1631 4.5005
R4563 VSS.n1656 VSS.n1593 4.5005
R4564 VSS.n1656 VSS.n1655 4.5005
R4565 VSS.n1681 VSS.n1680 4.5005
R4566 VSS.n1682 VSS.n1681 4.5005
R4567 VSS.n1667 VSS.n1582 4.5005
R4568 VSS.n1624 VSS.n1622 4.5005
R4569 VSS.n1504 VSS.n1502 4.5005
R4570 VSS.n1520 VSS.n1508 4.5005
R4571 VSS.n744 VSS.n415 3.69976
R4572 VSS.n1317 VSS.n1007 3.69976
R4573 VSS.n2050 VSS.n101 3.69976
R4574 VSS.n1728 VSS.n1400 3.69976
R4575 VSS.n1929 VSS.n176 3.69922
R4576 VSS.n1777 VSS.n282 3.69922
R4577 VSS.n967 VSS.n796 3.69922
R4578 VSS.n1767 VSS.n1365 3.42389
R4579 VSS.n379 VSS.n283 3.42389
R4580 VSS.n783 VSS.n380 3.42389
R4581 VSS.n971 VSS.n970 3.42389
R4582 VSS.n1356 VSS.n972 3.42389
R4583 VSS.n1935 VSS.n1934 3.42389
R4584 VSS.n1933 VSS.n1932 3.42389
R4585 VSS.n1514 VSS.n1401 3.423
R4586 VSS.n1816 VSS.n246 3.423
R4587 VSS.n530 VSS.n416 3.423
R4588 VSS.n875 VSS.n874 3.423
R4589 VSS.n1122 VSS.n1008 3.423
R4590 VSS.n2054 VSS.n2053 3.423
R4591 VSS.n1830 VSS.n1829 3.423
R4592 VSS.n674 VSS.n673 3.4105
R4593 VSS.n675 VSS.n674 3.4105
R4594 VSS.n672 VSS.n630 3.4105
R4595 VSS.n669 VSS.n633 3.4105
R4596 VSS.n669 VSS.n668 3.4105
R4597 VSS.n688 VSS.n687 3.4105
R4598 VSS.n687 VSS.n686 3.4105
R4599 VSS.n631 VSS.n627 3.4105
R4600 VSS.n627 VSS.n625 3.4105
R4601 VSS.n613 VSS.n595 3.4105
R4602 VSS.n613 VSS.n612 3.4105
R4603 VSS.n617 VSS.n593 3.4105
R4604 VSS.n690 VSS.n689 3.4105
R4605 VSS.n691 VSS.n690 3.4105
R4606 VSS.n706 VSS.n705 3.4105
R4607 VSS.n602 VSS.n601 3.4105
R4608 VSS.n551 VSS.n540 3.4105
R4609 VSS.n551 VSS.n545 3.4105
R4610 VSS.n553 VSS.n552 3.4105
R4611 VSS.n708 VSS.n707 3.4105
R4612 VSS.n726 VSS.n725 3.4105
R4613 VSS.n726 VSS.n519 3.4105
R4614 VSS.n723 VSS.n722 3.4105
R4615 VSS.n722 VSS.n721 3.4105
R4616 VSS.n1782 VSS.n1781 3.4105
R4617 VSS.n1781 VSS.n1780 3.4105
R4618 VSS.n1789 VSS.n1788 3.4105
R4619 VSS.n1784 VSS.n1783 3.4105
R4620 VSS.n1785 VSS.n1784 3.4105
R4621 VSS.n1797 VSS.n1796 3.4105
R4622 VSS.n1796 VSS.n1795 3.4105
R4623 VSS.n268 VSS.n263 3.4105
R4624 VSS.n1791 VSS.n1790 3.4105
R4625 VSS.n1791 VSS.n267 3.4105
R4626 VSS.n1805 VSS.n1804 3.4105
R4627 VSS.n1804 VSS.n1803 3.4105
R4628 VSS.n262 VSS.n260 3.4105
R4629 VSS.n1799 VSS.n1798 3.4105
R4630 VSS.n1799 VSS.n258 3.4105
R4631 VSS.n1812 VSS.n1811 3.4105
R4632 VSS.n1811 VSS.n1810 3.4105
R4633 VSS.n1807 VSS.n1806 3.4105
R4634 VSS.n1813 VSS.n247 3.4105
R4635 VSS.n247 VSS.n245 3.4105
R4636 VSS.n531 VSS.n529 3.4105
R4637 VSS.n529 VSS.n528 3.4105
R4638 VSS.n522 VSS.n521 3.4105
R4639 VSS.n539 VSS.n538 3.4105
R4640 VSS.n538 VSS.n537 3.4105
R4641 VSS.n749 VSS.n748 3.4105
R4642 VSS.n748 VSS.n747 3.4105
R4643 VSS.n756 VSS.n755 3.4105
R4644 VSS.n751 VSS.n750 3.4105
R4645 VSS.n752 VSS.n751 3.4105
R4646 VSS.n764 VSS.n763 3.4105
R4647 VSS.n763 VSS.n762 3.4105
R4648 VSS.n401 VSS.n397 3.4105
R4649 VSS.n758 VSS.n757 3.4105
R4650 VSS.n758 VSS.n400 3.4105
R4651 VSS.n772 VSS.n771 3.4105
R4652 VSS.n771 VSS.n770 3.4105
R4653 VSS.n396 VSS.n394 3.4105
R4654 VSS.n766 VSS.n765 3.4105
R4655 VSS.n766 VSS.n392 3.4105
R4656 VSS.n779 VSS.n778 3.4105
R4657 VSS.n778 VSS.n777 3.4105
R4658 VSS.n774 VSS.n773 3.4105
R4659 VSS.n780 VSS.n381 3.4105
R4660 VSS.n381 VSS.n378 3.4105
R4661 VSS.n1247 VSS.n1246 3.4105
R4662 VSS.n1248 VSS.n1247 3.4105
R4663 VSS.n1245 VSS.n1243 3.4105
R4664 VSS.n2197 VSS.n2196 3.4105
R4665 VSS.n2196 VSS.n2195 3.4105
R4666 VSS.n1261 VSS.n1260 3.4105
R4667 VSS.n1260 VSS.n1259 3.4105
R4668 VSS.n1244 VSS.n1238 3.4105
R4669 VSS.n1238 VSS.n1236 3.4105
R4670 VSS.n1205 VSS.n1187 3.4105
R4671 VSS.n1205 VSS.n1204 3.4105
R4672 VSS.n1209 VSS.n1185 3.4105
R4673 VSS.n1263 VSS.n1262 3.4105
R4674 VSS.n1264 VSS.n1263 3.4105
R4675 VSS.n1279 VSS.n1278 3.4105
R4676 VSS.n1194 VSS.n1193 3.4105
R4677 VSS.n1143 VSS.n1132 3.4105
R4678 VSS.n1143 VSS.n1137 3.4105
R4679 VSS.n1145 VSS.n1144 3.4105
R4680 VSS.n1281 VSS.n1280 3.4105
R4681 VSS.n1299 VSS.n1298 3.4105
R4682 VSS.n1299 VSS.n1111 3.4105
R4683 VSS.n1296 VSS.n1295 3.4105
R4684 VSS.n1295 VSS.n1294 3.4105
R4685 VSS.n950 VSS.n949 3.4105
R4686 VSS.n950 VSS.n795 3.4105
R4687 VSS.n943 VSS.n942 3.4105
R4688 VSS.n948 VSS.n947 3.4105
R4689 VSS.n947 VSS.n946 3.4105
R4690 VSS.n923 VSS.n922 3.4105
R4691 VSS.n923 VSS.n835 3.4105
R4692 VSS.n921 VSS.n920 3.4105
R4693 VSS.n941 VSS.n940 3.4105
R4694 VSS.n940 VSS.n939 3.4105
R4695 VSS.n910 VSS.n841 3.4105
R4696 VSS.n841 VSS.n840 3.4105
R4697 VSS.n839 VSS.n838 3.4105
R4698 VSS.n918 VSS.n917 3.4105
R4699 VSS.n917 VSS.n833 3.4105
R4700 VSS.n888 VSS.n887 3.4105
R4701 VSS.n888 VSS.n860 3.4105
R4702 VSS.n909 VSS.n908 3.4105
R4703 VSS.n886 VSS.n885 3.4105
R4704 VSS.n885 VSS.n884 3.4105
R4705 VSS.n1123 VSS.n1121 3.4105
R4706 VSS.n1121 VSS.n1120 3.4105
R4707 VSS.n1114 VSS.n1113 3.4105
R4708 VSS.n1131 VSS.n1130 3.4105
R4709 VSS.n1130 VSS.n1129 3.4105
R4710 VSS.n1322 VSS.n1321 3.4105
R4711 VSS.n1321 VSS.n1320 3.4105
R4712 VSS.n1329 VSS.n1328 3.4105
R4713 VSS.n1324 VSS.n1323 3.4105
R4714 VSS.n1325 VSS.n1324 3.4105
R4715 VSS.n1337 VSS.n1336 3.4105
R4716 VSS.n1336 VSS.n1335 3.4105
R4717 VSS.n993 VSS.n989 3.4105
R4718 VSS.n1331 VSS.n1330 3.4105
R4719 VSS.n1331 VSS.n992 3.4105
R4720 VSS.n1345 VSS.n1344 3.4105
R4721 VSS.n1344 VSS.n1343 3.4105
R4722 VSS.n988 VSS.n986 3.4105
R4723 VSS.n1339 VSS.n1338 3.4105
R4724 VSS.n1339 VSS.n984 3.4105
R4725 VSS.n1352 VSS.n1351 3.4105
R4726 VSS.n1351 VSS.n1350 3.4105
R4727 VSS.n1347 VSS.n1346 3.4105
R4728 VSS.n1353 VSS.n973 3.4105
R4729 VSS.n973 VSS.n792 3.4105
R4730 VSS.n2169 VSS.n2168 3.4105
R4731 VSS.n2152 VSS.n2151 3.4105
R4732 VSS.n2153 VSS.n2152 3.4105
R4733 VSS.n2149 VSS.n27 3.4105
R4734 VSS.n28 VSS.n27 3.4105
R4735 VSS.n2127 VSS.n2126 3.4105
R4736 VSS.n2127 VSS.n50 3.4105
R4737 VSS.n34 VSS.n33 3.4105
R4738 VSS.n2148 VSS.n2147 3.4105
R4739 VSS.n2147 VSS.n2146 3.4105
R4740 VSS.n2111 VSS.n2110 3.4105
R4741 VSS.n2123 VSS.n2122 3.4105
R4742 VSS.n2093 VSS.n2092 3.4105
R4743 VSS.n2094 VSS.n2093 3.4105
R4744 VSS.n2091 VSS.n79 3.4105
R4745 VSS.n2109 VSS.n2108 3.4105
R4746 VSS.n2069 VSS.n2064 3.4105
R4747 VSS.n2069 VSS.n2068 3.4105
R4748 VSS.n2090 VSS.n2089 3.4105
R4749 VSS.n2089 VSS.n2088 3.4105
R4750 VSS.n2055 VSS.n97 3.4105
R4751 VSS.n2034 VSS.n97 3.4105
R4752 VSS.n94 VSS.n93 3.4105
R4753 VSS.n2063 VSS.n2062 3.4105
R4754 VSS.n2062 VSS.n2061 3.4105
R4755 VSS.n2166 VSS.n24 3.4105
R4756 VSS.n2166 VSS.n2165 3.4105
R4757 VSS.n2019 VSS.n2018 3.4105
R4758 VSS.n2019 VSS.n100 3.4105
R4759 VSS.n1996 VSS.n1995 3.4105
R4760 VSS.n2017 VSS.n2016 3.4105
R4761 VSS.n2016 VSS.n2015 3.4105
R4762 VSS.n1986 VSS.n130 3.4105
R4763 VSS.n130 VSS.n129 3.4105
R4764 VSS.n1988 VSS.n1987 3.4105
R4765 VSS.n1994 VSS.n1993 3.4105
R4766 VSS.n1993 VSS.n1992 3.4105
R4767 VSS.n1969 VSS.n1968 3.4105
R4768 VSS.n1969 VSS.n144 3.4105
R4769 VSS.n1965 VSS.n132 3.4105
R4770 VSS.n1985 VSS.n1984 3.4105
R4771 VSS.n1984 VSS.n1983 3.4105
R4772 VSS.n1948 VSS.n1947 3.4105
R4773 VSS.n1948 VSS.n160 3.4105
R4774 VSS.n1964 VSS.n1963 3.4105
R4775 VSS.n1946 VSS.n1945 3.4105
R4776 VSS.n1945 VSS.n1944 3.4105
R4777 VSS.n2173 VSS.n2172 3.4105
R4778 VSS.n2174 VSS.n2173 3.4105
R4779 VSS.n1915 VSS.n1914 3.4105
R4780 VSS.n1915 VSS.n175 3.4105
R4781 VSS.n1891 VSS.n1890 3.4105
R4782 VSS.n1913 VSS.n1912 3.4105
R4783 VSS.n1912 VSS.n1911 3.4105
R4784 VSS.n1881 VSS.n205 3.4105
R4785 VSS.n205 VSS.n204 3.4105
R4786 VSS.n1883 VSS.n1882 3.4105
R4787 VSS.n1889 VSS.n1888 3.4105
R4788 VSS.n1888 VSS.n1887 3.4105
R4789 VSS.n1864 VSS.n1863 3.4105
R4790 VSS.n1864 VSS.n221 3.4105
R4791 VSS.n1860 VSS.n207 3.4105
R4792 VSS.n1880 VSS.n1879 3.4105
R4793 VSS.n1879 VSS.n1878 3.4105
R4794 VSS.n1843 VSS.n1842 3.4105
R4795 VSS.n1843 VSS.n235 3.4105
R4796 VSS.n1859 VSS.n1858 3.4105
R4797 VSS.n1841 VSS.n1840 3.4105
R4798 VSS.n1840 VSS.n1839 3.4105
R4799 VSS.n1638 VSS.n1592 3.4105
R4800 VSS.n1638 VSS.n1637 3.4105
R4801 VSS.n1641 VSS.n1640 3.4105
R4802 VSS.n1644 VSS.n1643 3.4105
R4803 VSS.n1645 VSS.n1644 3.4105
R4804 VSS.n1662 VSS.n1661 3.4105
R4805 VSS.n1663 VSS.n1662 3.4105
R4806 VSS.n1659 VSS.n1658 3.4105
R4807 VSS.n1658 VSS.n1657 3.4105
R4808 VSS.n1677 VSS.n1676 3.4105
R4809 VSS.n1676 VSS.n1675 3.4105
R4810 VSS.n1590 VSS.n1589 3.4105
R4811 VSS.n1591 VSS.n1583 3.4105
R4812 VSS.n1583 VSS.n1579 3.4105
R4813 VSS.n1573 VSS.n1572 3.4105
R4814 VSS.n1679 VSS.n1678 3.4105
R4815 VSS.n1694 VSS.n1541 3.4105
R4816 VSS.n1694 VSS.n1693 3.4105
R4817 VSS.n1558 VSS.n1534 3.4105
R4818 VSS.n1561 VSS.n1554 3.4105
R4819 VSS.n1710 VSS.n1524 3.4105
R4820 VSS.n1710 VSS.n1709 3.4105
R4821 VSS.n1540 VSS.n1539 3.4105
R4822 VSS.n1539 VSS.n1538 3.4105
R4823 VSS.n1733 VSS.n1732 3.4105
R4824 VSS.n1732 VSS.n1731 3.4105
R4825 VSS.n1740 VSS.n1739 3.4105
R4826 VSS.n1735 VSS.n1734 3.4105
R4827 VSS.n1736 VSS.n1735 3.4105
R4828 VSS.n1748 VSS.n1747 3.4105
R4829 VSS.n1747 VSS.n1746 3.4105
R4830 VSS.n1386 VSS.n1382 3.4105
R4831 VSS.n1742 VSS.n1741 3.4105
R4832 VSS.n1742 VSS.n1385 3.4105
R4833 VSS.n1756 VSS.n1755 3.4105
R4834 VSS.n1755 VSS.n1754 3.4105
R4835 VSS.n1381 VSS.n1379 3.4105
R4836 VSS.n1750 VSS.n1749 3.4105
R4837 VSS.n1750 VSS.n1377 3.4105
R4838 VSS.n1763 VSS.n1762 3.4105
R4839 VSS.n1762 VSS.n1761 3.4105
R4840 VSS.n1758 VSS.n1757 3.4105
R4841 VSS.n1764 VSS.n1366 3.4105
R4842 VSS.n1366 VSS.n1364 3.4105
R4843 VSS.n1515 VSS.n1513 3.4105
R4844 VSS.n1513 VSS.n1512 3.4105
R4845 VSS.n1507 VSS.n1506 3.4105
R4846 VSS.n1523 VSS.n1522 3.4105
R4847 VSS.n1522 VSS.n1521 3.4105
R4848 VSS.n1427 VSS.n1426 3.29193
R4849 VSS.n1447 VSS.n1446 3.29193
R4850 VSS.n1466 VSS.n1411 3.29193
R4851 VSS.n310 VSS.n309 3.29193
R4852 VSS.n328 VSS.n327 3.29193
R4853 VSS.n347 VSS.n293 3.29193
R4854 VSS.n525 VSS.n515 3.29193
R4855 VSS.n657 VSS.n638 3.29193
R4856 VSS.n442 VSS.n441 3.29193
R4857 VSS.n462 VSS.n461 3.29193
R4858 VSS.n481 VSS.n426 3.29193
R4859 VSS.n866 VSS.n855 3.29193
R4860 VSS.n893 VSS.n849 3.29193
R4861 VSS.n828 VSS.n827 3.29193
R4862 VSS.n1117 VSS.n1107 3.29193
R4863 VSS.n1216 VSS.n5 3.29193
R4864 VSS.n1034 VSS.n1033 3.29193
R4865 VSS.n1054 VSS.n1053 3.29193
R4866 VSS.n1073 VSS.n1018 3.29193
R4867 VSS.n166 VSS.n156 3.29193
R4868 VSS.n1959 VSS.n1958 3.29193
R4869 VSS.n1997 VSS.n117 3.29193
R4870 VSS.n2038 VSS.n2037 3.29193
R4871 VSS.n2177 VSS.n2176 3.29193
R4872 VSS.n241 VSS.n231 3.29193
R4873 VSS.n1854 VSS.n1853 3.29193
R4874 VSS.n1892 VSS.n192 3.29193
R4875 VSS.n1509 VSS.n1500 3.29193
R4876 VSS.n1648 VSS.n1647 3.29193
R4877 VSS.n1489 VSS.n1488 3.2005
R4878 VSS.n371 VSS.n370 3.2005
R4879 VSS.n504 VSS.n503 3.2005
R4880 VSS.n809 VSS.n808 3.2005
R4881 VSS.n1096 VSS.n1095 3.2005
R4882 VSS.n2027 VSS.n2026 3.2005
R4883 VSS.n1923 VSS.n1922 3.2005
R4884 VSS.n430 VSS.n399 3.03311
R4885 VSS.n454 VSS.n453 3.03311
R4886 VSS.n1022 VSS.n991 3.03311
R4887 VSS.n1046 VSS.n1045 3.03311
R4888 VSS.n1982 VSS.n1981 3.03311
R4889 VSS.n1952 VSS.n1951 3.03311
R4890 VSS.n1877 VSS.n1876 3.03311
R4891 VSS.n1847 VSS.n1846 3.03311
R4892 VSS.n298 VSS.n297 3.03311
R4893 VSS.n322 VSS.n321 3.03311
R4894 VSS.n927 VSS.n926 3.03311
R4895 VSS.n892 VSS.n891 3.03311
R4896 VSS.n1415 VSS.n1384 3.03311
R4897 VSS.n1439 VSS.n1438 3.03311
R4898 VSS.n1453 VSS.n1418 2.81479
R4899 VSS.n1474 VSS.n1414 2.81479
R4900 VSS.n902 VSS.n852 2.81479
R4901 VSS.n935 VSS.n822 2.81479
R4902 VSS.n334 VSS.n301 2.81479
R4903 VSS.n355 VSS.n296 2.81479
R4904 VSS.n1870 VSS.n218 2.81479
R4905 VSS.n1901 VSS.n195 2.81479
R4906 VSS.n468 VSS.n433 2.81479
R4907 VSS.n489 VSS.n429 2.81479
R4908 VSS.n1060 VSS.n1025 2.81479
R4909 VSS.n1081 VSS.n1021 2.81479
R4910 VSS.n1975 VSS.n141 2.81479
R4911 VSS.n2006 VSS.n120 2.81479
R4912 VSS.n694 VSS.n693 2.5605
R4913 VSS.n1267 VSS.n1266 2.5605
R4914 VSS.n2133 VSS.n2132 2.5605
R4915 VSS.n1672 VSS.n1580 2.5605
R4916 VSS.n712 VSS.n547 2.46907
R4917 VSS.n1285 VSS.n1139 2.46907
R4918 VSS.n2097 VSS.n2096 2.46907
R4919 VSS.n1691 VSS.n1690 2.46907
R4920 VSS.n932 VSS.t16 2.42341
R4921 VSS.n684 VSS.n623 2.37764
R4922 VSS.n1257 VSS.n1215 2.37764
R4923 VSS.n2138 VSS.n29 2.37764
R4924 VSS.n1616 VSS.n1615 2.37764
R4925 VSS.n570 VSS.n568 2.28621
R4926 VSS.n1162 VSS.n1160 2.28621
R4927 VSS.n2065 VSS.n84 2.28621
R4928 VSS.n1706 VSS.n1705 2.28621
R4929 VSS.n2200 VSS.n2199 2.27261
R4930 VSS.n1399 VSS.n1397 2.2505
R4931 VSS.n1465 VSS.n1388 2.2505
R4932 VSS.n1395 VSS.n1394 2.2505
R4933 VSS.n1370 VSS.n1368 2.2505
R4934 VSS.n1376 VSS.n1374 2.2505
R4935 VSS.n1431 VSS.n1430 2.2505
R4936 VSS.n281 VSS.n279 2.2505
R4937 VSS.n346 VSS.n270 2.2505
R4938 VSS.n277 VSS.n276 2.2505
R4939 VSS.n251 VSS.n249 2.2505
R4940 VSS.n257 VSS.n255 2.2505
R4941 VSS.n314 VSS.n313 2.2505
R4942 VSS.n679 VSS.n626 2.2505
R4943 VSS.n611 VSS.n596 2.2505
R4944 VSS.n649 VSS.n648 2.2505
R4945 VSS.n719 VSS.n718 2.2505
R4946 VSS.n550 VSS.n548 2.2505
R4947 VSS.n580 VSS.n556 2.2505
R4948 VSS.n729 VSS.n518 2.2505
R4949 VSS.n414 VSS.n412 2.2505
R4950 VSS.n480 VSS.n403 2.2505
R4951 VSS.n410 VSS.n409 2.2505
R4952 VSS.n385 VSS.n383 2.2505
R4953 VSS.n391 VSS.n389 2.2505
R4954 VSS.n446 VSS.n445 2.2505
R4955 VSS.n952 VSS.n951 2.2505
R4956 VSS.n938 VSS.n817 2.2505
R4957 VSS.n804 VSS.n802 2.2505
R4958 VSS.n890 VSS.n889 2.2505
R4959 VSS.n847 VSS.n846 2.2505
R4960 VSS.n883 VSS.n864 2.2505
R4961 VSS.n1252 VSS.n1237 2.2505
R4962 VSS.n1203 VSS.n1188 2.2505
R4963 VSS.n1226 VSS.n1225 2.2505
R4964 VSS.n1292 VSS.n1291 2.2505
R4965 VSS.n1142 VSS.n1140 2.2505
R4966 VSS.n1172 VSS.n1148 2.2505
R4967 VSS.n1302 VSS.n1110 2.2505
R4968 VSS.n1006 VSS.n1004 2.2505
R4969 VSS.n1072 VSS.n995 2.2505
R4970 VSS.n1002 VSS.n1001 2.2505
R4971 VSS.n977 VSS.n975 2.2505
R4972 VSS.n983 VSS.n981 2.2505
R4973 VSS.n1038 VSS.n1037 2.2505
R4974 VSS.n2021 VSS.n2020 2.2505
R4975 VSS.n125 VSS.n123 2.2505
R4976 VSS.n2014 VSS.n112 2.2505
R4977 VSS.n1950 VSS.n1949 2.2505
R4978 VSS.n1971 VSS.n1970 2.2505
R4979 VSS.n1943 VSS.n164 2.2505
R4980 VSS.n2072 VSS.n2071 2.2505
R4981 VSS.n2086 VSS.n2085 2.2505
R4982 VSS.n2106 VSS.n62 2.2505
R4983 VSS.n2129 VSS.n2128 2.2505
R4984 VSS.n42 VSS.n41 2.2505
R4985 VSS.n2160 VSS.n26 2.2505
R4986 VSS.n64 VSS.n59 2.2505
R4987 VSS.n1917 VSS.n1916 2.2505
R4988 VSS.n200 VSS.n198 2.2505
R4989 VSS.n1910 VSS.n187 2.2505
R4990 VSS.n1845 VSS.n1844 2.2505
R4991 VSS.n1866 VSS.n1865 2.2505
R4992 VSS.n1838 VSS.n239 2.2505
R4993 VSS.n1632 VSS.n1595 2.2505
R4994 VSS.n1578 VSS.n1576 2.2505
R4995 VSS.n1666 VSS.n1665 2.2505
R4996 VSS.n1533 VSS.n1531 2.2505
R4997 VSS.n1563 VSS.n1562 2.2505
R4998 VSS.n1565 VSS.n1555 2.2505
R4999 VSS.n1713 VSS.n1712 2.2505
R5000 VSS.n2199 VSS.n0 2.24315
R5001 VSS.n701 VSS.n561 2.10336
R5002 VSS.n1274 VSS.n1153 2.10336
R5003 VSS.n2116 VSS.n57 2.10336
R5004 VSS.n1683 VSS.n1682 2.10336
R5005 VSS.n702 VSS.n701 2.01193
R5006 VSS.n1275 VSS.n1274 2.01193
R5007 VSS.n66 VSS.n57 2.01193
R5008 VSS.n1683 VSS.n1548 2.01193
R5009 VSS.n1769 VSS.n1768 1.98071
R5010 VSS.n1831 VSS.n1828 1.98071
R5011 VSS.n785 VSS.n784 1.98071
R5012 VSS.n1818 VSS.n1817 1.98071
R5013 VSS.n1358 VSS.n1357 1.98071
R5014 VSS.n876 VSS.n873 1.98071
R5015 VSS.n1936 VSS.n172 1.98071
R5016 VSS.n709 VSS.n708 1.94045
R5017 VSS.n1282 VSS.n1281 1.94045
R5018 VSS.n2108 VSS.n2107 1.94045
R5019 VSS.n1561 VSS.n1557 1.94045
R5020 VSS VSS.n0 1.85712
R5021 VSS.n1439 VSS.n1427 1.55479
R5022 VSS.n322 VSS.n310 1.55479
R5023 VSS.n454 VSS.n442 1.55479
R5024 VSS.n892 VSS.n855 1.55479
R5025 VSS.n1046 VSS.n1034 1.55479
R5026 VSS.n1952 VSS.n156 1.55479
R5027 VSS.n1847 VSS.n231 1.55479
R5028 VSS.n584 VSS.n576 1.53956
R5029 VSS.n696 VSS.n588 1.53956
R5030 VSS.n1176 VSS.n1168 1.53956
R5031 VSS.n1269 VSS.n1180 1.53956
R5032 VSS.n2098 VSS.n72 1.53956
R5033 VSS.n2135 VSS.n44 1.53956
R5034 VSS.n1688 VSS.n1529 1.53956
R5035 VSS.n1613 VSS.n1610 1.53956
R5036 VSS.n266 VSS.n264 1.5005
R5037 VSS.n925 VSS.n924 1.5005
R5038 VSS.n212 VSS.n211 1.5005
R5039 VSS.n1480 VSS.n1406 1.46336
R5040 VSS.n362 VSS.n288 1.46336
R5041 VSS.n583 VSS.n582 1.46336
R5042 VSS.n695 VSS.n589 1.46336
R5043 VSS.n495 VSS.n421 1.46336
R5044 VSS.n807 VSS.n801 1.46336
R5045 VSS.n1175 VSS.n1174 1.46336
R5046 VSS.n1268 VSS.n1181 1.46336
R5047 VSS.n1087 VSS.n1013 1.46336
R5048 VSS.n2011 VSS.n106 1.46336
R5049 VSS.n2104 VSS.n65 1.46336
R5050 VSS.n2134 VSS.n2131 1.46336
R5051 VSS.n1907 VSS.n181 1.46336
R5052 VSS.n1689 VSS.n1544 1.46336
R5053 VSS.n1609 VSS.n1608 1.46336
R5054 VSS.n1446 VSS.n1419 1.37193
R5055 VSS.n1456 VSS.n1455 1.37193
R5056 VSS.n1463 VSS.n1462 1.37193
R5057 VSS.n1466 VSS.n1464 1.37193
R5058 VSS.n327 VSS.n302 1.37193
R5059 VSS.n337 VSS.n336 1.37193
R5060 VSS.n344 VSS.n343 1.37193
R5061 VSS.n347 VSS.n345 1.37193
R5062 VSS.n461 VSS.n434 1.37193
R5063 VSS.n471 VSS.n470 1.37193
R5064 VSS.n478 VSS.n477 1.37193
R5065 VSS.n481 VSS.n479 1.37193
R5066 VSS.n904 VSS.n849 1.37193
R5067 VSS.n850 VSS.n832 1.37193
R5068 VSS.n928 VSS.n820 1.37193
R5069 VSS.n827 VSS.n821 1.37193
R5070 VSS.n1053 VSS.n1026 1.37193
R5071 VSS.n1063 VSS.n1062 1.37193
R5072 VSS.n1070 VSS.n1069 1.37193
R5073 VSS.n1073 VSS.n1071 1.37193
R5074 VSS.n1959 VSS.n142 1.37193
R5075 VSS.n1974 VSS.n136 1.37193
R5076 VSS.n137 VSS.n121 1.37193
R5077 VSS.n1997 VSS.n122 1.37193
R5078 VSS.n1854 VSS.n219 1.37193
R5079 VSS.n1869 VSS.n213 1.37193
R5080 VSS.n214 VSS.n196 1.37193
R5081 VSS.n1892 VSS.n197 1.37193
R5082 VSS.n569 VSS.n546 1.2805
R5083 VSS.n651 VSS.n645 1.2805
R5084 VSS.n1161 VSS.n1138 1.2805
R5085 VSS.n1229 VSS.n1228 1.2805
R5086 VSS.n2081 VSS.n2079 1.2805
R5087 VSS.n2143 VSS.n39 1.2805
R5088 VSS.n1699 VSS.n1526 1.2805
R5089 VSS.n1617 VSS.n1581 1.2805
R5090 VSS.n1448 VSS.n1447 1.18907
R5091 VSS.n1478 VSS.n1411 1.18907
R5092 VSS.n329 VSS.n328 1.18907
R5093 VSS.n360 VSS.n293 1.18907
R5094 VSS.n463 VSS.n462 1.18907
R5095 VSS.n493 VSS.n426 1.18907
R5096 VSS.n894 VSS.n893 1.18907
R5097 VSS.n828 VSS.n800 1.18907
R5098 VSS.n1055 VSS.n1054 1.18907
R5099 VSS.n1085 VSS.n1018 1.18907
R5100 VSS.n1958 VSS.n153 1.18907
R5101 VSS.n2010 VSS.n117 1.18907
R5102 VSS.n1853 VSS.n228 1.18907
R5103 VSS.n1906 VSS.n192 1.18907
R5104 VSS.n1815 VSS.n1814 1.13717
R5105 VSS.n250 VSS.n248 1.13717
R5106 VSS.n259 VSS.n254 1.13717
R5107 VSS.n271 VSS.n269 1.13717
R5108 VSS.n274 VSS.n272 1.13717
R5109 VSS.n280 VSS.n278 1.13717
R5110 VSS.n533 VSS.n532 1.13717
R5111 VSS.n554 VSS.n549 1.13717
R5112 VSS.n616 VSS.n615 1.13717
R5113 VSS.n671 VSS.n670 1.13717
R5114 VSS.n782 VSS.n781 1.13717
R5115 VSS.n384 VSS.n382 1.13717
R5116 VSS.n393 VSS.n388 1.13717
R5117 VSS.n404 VSS.n402 1.13717
R5118 VSS.n407 VSS.n405 1.13717
R5119 VSS.n413 VSS.n411 1.13717
R5120 VSS.n863 VSS.n862 1.13717
R5121 VSS.n861 VSS.n842 1.13717
R5122 VSS.n912 VSS.n911 1.13717
R5123 VSS.n919 VSS.n815 1.13717
R5124 VSS.n812 VSS.n811 1.13717
R5125 VSS.n794 VSS.n793 1.13717
R5126 VSS.n1125 VSS.n1124 1.13717
R5127 VSS.n1146 VSS.n1141 1.13717
R5128 VSS.n1208 VSS.n1207 1.13717
R5129 VSS.n2 VSS.n1 1.13717
R5130 VSS.n1355 VSS.n1354 1.13717
R5131 VSS.n976 VSS.n974 1.13717
R5132 VSS.n985 VSS.n980 1.13717
R5133 VSS.n996 VSS.n994 1.13717
R5134 VSS.n999 VSS.n997 1.13717
R5135 VSS.n1005 VSS.n1003 1.13717
R5136 VSS.n2170 VSS.n23 1.13717
R5137 VSS.n163 VSS.n162 1.13717
R5138 VSS.n161 VSS.n148 1.13717
R5139 VSS.n1967 VSS.n1966 1.13717
R5140 VSS.n131 VSS.n127 1.13717
R5141 VSS.n111 VSS.n110 1.13717
R5142 VSS.n99 VSS.n98 1.13717
R5143 VSS.n2057 VSS.n2056 1.13717
R5144 VSS.n61 VSS.n60 1.13717
R5145 VSS.n2125 VSS.n2124 1.13717
R5146 VSS.n238 VSS.n237 1.13717
R5147 VSS.n236 VSS.n225 1.13717
R5148 VSS.n1862 VSS.n1861 1.13717
R5149 VSS.n206 VSS.n202 1.13717
R5150 VSS.n186 VSS.n185 1.13717
R5151 VSS.n174 VSS.n173 1.13717
R5152 VSS.n1766 VSS.n1765 1.13717
R5153 VSS.n1369 VSS.n1367 1.13717
R5154 VSS.n1378 VSS.n1373 1.13717
R5155 VSS.n1389 VSS.n1387 1.13717
R5156 VSS.n1392 VSS.n1390 1.13717
R5157 VSS.n1398 VSS.n1396 1.13717
R5158 VSS.n1517 VSS.n1516 1.13717
R5159 VSS.n1560 VSS.n1559 1.13717
R5160 VSS.n1588 VSS.n1575 1.13717
R5161 VSS.n1642 VSS.n1625 1.13717
R5162 VSS.n1384 VSS.n1380 1.1255
R5163 VSS.n399 VSS.n395 1.1255
R5164 VSS.n991 VSS.n987 1.1255
R5165 VSS.n1982 VSS.n134 1.1255
R5166 VSS.n731 VSS.n730 1.09764
R5167 VSS.n658 VSS.n624 1.09764
R5168 VSS.n1304 VSS.n1303 1.09764
R5169 VSS.n1235 VSS.n1217 1.09764
R5170 VSS.n2073 VSS.n88 1.09764
R5171 VSS.n2178 VSS.n20 1.09764
R5172 VSS.n1715 VSS.n1714 1.09764
R5173 VSS.n1654 VSS.n1597 1.09764
R5174 VSS.n559 VSS.n557 1.04225
R5175 VSS.n1151 VSS.n1149 1.04225
R5176 VSS.n2114 VSS.n2113 1.04225
R5177 VSS.n1552 VSS.n1550 1.04225
R5178 VSS.n1426 VSS.n1363 1.00621
R5179 VSS.n1489 VSS.n1402 1.00621
R5180 VSS.n309 VSS.n244 1.00621
R5181 VSS.n371 VSS.n284 1.00621
R5182 VSS.n730 VSS.n516 1.00621
R5183 VSS.n568 VSS.n567 1.00621
R5184 VSS.n608 VSS.n607 1.00621
R5185 VSS.n441 VSS.n377 1.00621
R5186 VSS.n504 VSS.n417 1.00621
R5187 VSS.n872 VSS.n866 1.00621
R5188 VSS.n808 VSS.n797 1.00621
R5189 VSS.n1303 VSS.n1108 1.00621
R5190 VSS.n1160 VSS.n1159 1.00621
R5191 VSS.n1200 VSS.n1199 1.00621
R5192 VSS.n1033 VSS.n791 1.00621
R5193 VSS.n1096 VSS.n1009 1.00621
R5194 VSS.n171 VSS.n166 1.00621
R5195 VSS.n2027 VSS.n102 1.00621
R5196 VSS.n2073 VSS.n89 1.00621
R5197 VSS.n2066 VSS.n2065 1.00621
R5198 VSS.n2118 VSS.n48 1.00621
R5199 VSS.n1827 VSS.n241 1.00621
R5200 VSS.n1923 VSS.n177 1.00621
R5201 VSS.n1714 VSS.n1501 1.00621
R5202 VSS.n1707 VSS.n1706 1.00621
R5203 VSS.n1602 VSS.n1601 1.00621
R5204 VSS.n737 VSS.n510 0.914786
R5205 VSS.n578 VSS.n577 0.914786
R5206 VSS.n702 VSS.n560 0.914786
R5207 VSS.n684 VSS.n683 0.914786
R5208 VSS.n682 VSS.n624 0.914786
R5209 VSS.n666 VSS.n665 0.914786
R5210 VSS.n1310 VSS.n1102 0.914786
R5211 VSS.n1170 VSS.n1169 0.914786
R5212 VSS.n1275 VSS.n1152 0.914786
R5213 VSS.n1257 VSS.n1256 0.914786
R5214 VSS.n1255 VSS.n1235 0.914786
R5215 VSS.n2193 VSS.n2192 0.914786
R5216 VSS.n2043 VSS.n2033 0.914786
R5217 VSS.n71 VSS.n70 0.914786
R5218 VSS.n67 VSS.n66 0.914786
R5219 VSS.n2156 VSS.n29 0.914786
R5220 VSS.n2157 VSS.n20 0.914786
R5221 VSS.n2184 VSS.n15 0.914786
R5222 VSS.n1721 VSS.n1495 0.914786
R5223 VSS.n1567 VSS.n1566 0.914786
R5224 VSS.n1568 VSS.n1548 0.914786
R5225 VSS.n1615 VSS.n1596 0.914786
R5226 VSS.n1655 VSS.n1654 0.914786
R5227 VSS.n1629 VSS.n1622 0.914786
R5228 VSS.n669 VSS.n635 0.908949
R5229 VSS.n2196 VSS.n3 0.908949
R5230 VSS.n2173 VSS.n16 0.908949
R5231 VSS.n1644 VSS.n1630 0.908949
R5232 VSS.n529 VSS.n511 0.908879
R5233 VSS.n1121 VSS.n1103 0.908879
R5234 VSS.n2036 VSS.n97 0.908879
R5235 VSS.n1513 VSS.n1496 0.908879
R5236 VSS.n724 VSS.n520 0.853
R5237 VSS.n557 VSS.n555 0.853
R5238 VSS.n620 VSS.n618 0.853
R5239 VSS.n1297 VSS.n1112 0.853
R5240 VSS.n1149 VSS.n1147 0.853
R5241 VSS.n1212 VSS.n1210 0.853
R5242 VSS.n81 VSS.n80 0.853
R5243 VSS.n2113 VSS.n54 0.853
R5244 VSS.n2150 VSS.n32 0.853
R5245 VSS.n1535 VSS.n1505 0.853
R5246 VSS.n1574 VSS.n1552 0.853
R5247 VSS.n1660 VSS.n1587 0.853
R5248 VSS.n714 VSS.n546 0.823357
R5249 VSS.n713 VSS.n712 0.823357
R5250 VSS.n599 VSS.n561 0.823357
R5251 VSS.n644 VSS.n590 0.823357
R5252 VSS.n1287 VSS.n1138 0.823357
R5253 VSS.n1286 VSS.n1285 0.823357
R5254 VSS.n1191 VSS.n1153 0.823357
R5255 VSS.n1222 VSS.n1182 0.823357
R5256 VSS.n2081 VSS.n2080 0.823357
R5257 VSS.n2096 VSS.n76 0.823357
R5258 VSS.n2117 VSS.n2116 0.823357
R5259 VSS.n2144 VSS.n37 0.823357
R5260 VSS.n1699 VSS.n1530 0.823357
R5261 VSS.n1691 VSS.n1542 0.823357
R5262 VSS.n1682 VSS.n1549 0.823357
R5263 VSS.n1671 VSS.n1670 0.823357
R5264 VSS.n714 VSS.n713 0.731929
R5265 VSS.n693 VSS.n590 0.731929
R5266 VSS.n651 VSS.n644 0.731929
R5267 VSS.n1287 VSS.n1286 0.731929
R5268 VSS.n1266 VSS.n1182 0.731929
R5269 VSS.n1228 VSS.n1222 0.731929
R5270 VSS.n2080 VSS.n76 0.731929
R5271 VSS.n2132 VSS.n37 0.731929
R5272 VSS.n2144 VSS.n2143 0.731929
R5273 VSS.n1542 VSS.n1530 0.731929
R5274 VSS.n1672 VSS.n1671 0.731929
R5275 VSS.n1670 VSS.n1581 0.731929
R5276 VSS.n525 VSS.n510 0.6405
R5277 VSS.n582 VSS.n577 0.6405
R5278 VSS.n683 VSS.n682 0.6405
R5279 VSS.n666 VSS.n638 0.6405
R5280 VSS.n1117 VSS.n1102 0.6405
R5281 VSS.n1174 VSS.n1169 0.6405
R5282 VSS.n1256 VSS.n1255 0.6405
R5283 VSS.n2193 VSS.n5 0.6405
R5284 VSS.n2037 VSS.n2033 0.6405
R5285 VSS.n2104 VSS.n71 0.6405
R5286 VSS.n2157 VSS.n2156 0.6405
R5287 VSS.n2176 VSS.n15 0.6405
R5288 VSS.n1509 VSS.n1495 0.6405
R5289 VSS.n1566 VSS.n1544 0.6405
R5290 VSS.n1655 VSS.n1596 0.6405
R5291 VSS.n1647 VSS.n1622 0.6405
R5292 VSS.n567 VSS.n516 0.549071
R5293 VSS.n608 VSS.n589 0.549071
R5294 VSS.n1159 VSS.n1108 0.549071
R5295 VSS.n1200 VSS.n1181 0.549071
R5296 VSS.n2066 VSS.n89 0.549071
R5297 VSS.n2131 VSS.n48 0.549071
R5298 VSS.n1707 VSS.n1501 0.549071
R5299 VSS.n1608 VSS.n1601 0.549071
R5300 VSS.n531 VSS 0.517836
R5301 VSS.n1123 VSS 0.517836
R5302 VSS.n2055 VSS 0.517836
R5303 VSS.n1515 VSS 0.517836
R5304 VSS.n1769 VSS.n1363 0.465127
R5305 VSS.n1818 VSS.n244 0.465127
R5306 VSS.n785 VSS.n377 0.465127
R5307 VSS.n873 VSS.n872 0.465127
R5308 VSS.n1358 VSS.n791 0.465127
R5309 VSS.n172 VSS.n171 0.465127
R5310 VSS.n1828 VSS.n1827 0.465127
R5311 VSS.n1729 VSS.n1402 0.457643
R5312 VSS.n1778 VSS.n284 0.457643
R5313 VSS.n731 VSS.n515 0.457643
R5314 VSS.n658 VSS.n657 0.457643
R5315 VSS.n745 VSS.n417 0.457643
R5316 VSS.n968 VSS.n797 0.457643
R5317 VSS.n1304 VSS.n1107 0.457643
R5318 VSS.n1217 VSS.n1216 0.457643
R5319 VSS.n1318 VSS.n1009 0.457643
R5320 VSS.n2051 VSS.n102 0.457643
R5321 VSS.n2038 VSS.n88 0.457643
R5322 VSS.n2178 VSS.n2177 0.457643
R5323 VSS.n1930 VSS.n177 0.457643
R5324 VSS.n1715 VSS.n1500 0.457643
R5325 VSS.n1648 VSS.n1597 0.457643
R5326 VSS.n2171 VSS 0.415989
R5327 VSS.n1448 VSS.n1439 0.366214
R5328 VSS.n1479 VSS.n1478 0.366214
R5329 VSS.n329 VSS.n322 0.366214
R5330 VSS.n361 VSS.n360 0.366214
R5331 VSS.n463 VSS.n454 0.366214
R5332 VSS.n494 VSS.n493 0.366214
R5333 VSS.n894 VSS.n892 0.366214
R5334 VSS.n960 VSS.n800 0.366214
R5335 VSS.n1055 VSS.n1046 0.366214
R5336 VSS.n1086 VSS.n1085 0.366214
R5337 VSS.n1952 VSS.n153 0.366214
R5338 VSS.n2012 VSS.n2010 0.366214
R5339 VSS.n1847 VSS.n228 0.366214
R5340 VSS.n1908 VSS.n1906 0.366214
R5341 VSS.n246 VSS 0.301636
R5342 VSS.n874 VSS 0.301636
R5343 VSS.n1829 VSS 0.301636
R5344 VSS.n1365 VSS 0.301636
R5345 VSS.n633 VSS 0.300964
R5346 VSS VSS.n2197 0.300964
R5347 VSS.n2172 VSS 0.300964
R5348 VSS.n1643 VSS 0.300964
R5349 VSS.n380 VSS 0.29425
R5350 VSS.n972 VSS 0.29425
R5351 VSS.n1934 VSS 0.29425
R5352 VSS.n570 VSS.n569 0.274786
R5353 VSS.n578 VSS.n560 0.274786
R5354 VSS.n607 VSS.n599 0.274786
R5355 VSS.n645 VSS.n623 0.274786
R5356 VSS.n1162 VSS.n1161 0.274786
R5357 VSS.n1170 VSS.n1152 0.274786
R5358 VSS.n1199 VSS.n1191 0.274786
R5359 VSS.n1229 VSS.n1215 0.274786
R5360 VSS.n2079 VSS.n84 0.274786
R5361 VSS.n70 VSS.n67 0.274786
R5362 VSS.n2118 VSS.n2117 0.274786
R5363 VSS.n2138 VSS.n39 0.274786
R5364 VSS.n1705 VSS.n1526 0.274786
R5365 VSS.n1568 VSS.n1567 0.274786
R5366 VSS.n1602 VSS.n1549 0.274786
R5367 VSS.n1617 VSS.n1616 0.274786
R5368 VSS VSS.n379 0.206964
R5369 VSS VSS.n971 0.206964
R5370 VSS VSS.n1933 0.206964
R5371 VSS.n1454 VSS.n1419 0.183357
R5372 VSS.n1455 VSS.n1454 0.183357
R5373 VSS.n1473 VSS.n1463 0.183357
R5374 VSS.n1473 VSS.n1464 0.183357
R5375 VSS.n335 VSS.n302 0.183357
R5376 VSS.n336 VSS.n335 0.183357
R5377 VSS.n354 VSS.n344 0.183357
R5378 VSS.n354 VSS.n345 0.183357
R5379 VSS.n469 VSS.n434 0.183357
R5380 VSS.n470 VSS.n469 0.183357
R5381 VSS.n488 VSS.n478 0.183357
R5382 VSS.n488 VSS.n479 0.183357
R5383 VSS.n904 VSS.n903 0.183357
R5384 VSS.n903 VSS.n850 0.183357
R5385 VSS.n936 VSS.n820 0.183357
R5386 VSS.n936 VSS.n821 0.183357
R5387 VSS.n1061 VSS.n1026 0.183357
R5388 VSS.n1062 VSS.n1061 0.183357
R5389 VSS.n1080 VSS.n1070 0.183357
R5390 VSS.n1080 VSS.n1071 0.183357
R5391 VSS.n1973 VSS.n142 0.183357
R5392 VSS.n1974 VSS.n1973 0.183357
R5393 VSS.n2005 VSS.n121 0.183357
R5394 VSS.n2005 VSS.n122 0.183357
R5395 VSS.n1868 VSS.n219 0.183357
R5396 VSS.n1869 VSS.n1868 0.183357
R5397 VSS.n1900 VSS.n196 0.183357
R5398 VSS.n1900 VSS.n197 0.183357
R5399 VSS VSS.n632 0.107929
R5400 VSS.n2198 VSS 0.107929
R5401 VSS VSS.n2171 0.107929
R5402 VSS.n2200 VSS 0.107929
R5403 VSS VSS.n530 0.107593
R5404 VSS VSS.n1122 0.107593
R5405 VSS VSS.n2054 0.107593
R5406 VSS VSS.n1514 0.107593
R5407 VSS.n1480 VSS.n1479 0.0919286
R5408 VSS.n1488 VSS.n1406 0.0919286
R5409 VSS.n1729 VSS.n1728 0.0919286
R5410 VSS.n362 VSS.n361 0.0919286
R5411 VSS.n370 VSS.n288 0.0919286
R5412 VSS.n1778 VSS.n1777 0.0919286
R5413 VSS.n583 VSS.n547 0.0919286
R5414 VSS.n695 VSS.n694 0.0919286
R5415 VSS.n495 VSS.n494 0.0919286
R5416 VSS.n503 VSS.n421 0.0919286
R5417 VSS.n745 VSS.n744 0.0919286
R5418 VSS.n960 VSS.n801 0.0919286
R5419 VSS.n809 VSS.n807 0.0919286
R5420 VSS.n968 VSS.n967 0.0919286
R5421 VSS.n1175 VSS.n1139 0.0919286
R5422 VSS.n1268 VSS.n1267 0.0919286
R5423 VSS.n1087 VSS.n1086 0.0919286
R5424 VSS.n1095 VSS.n1013 0.0919286
R5425 VSS.n1318 VSS.n1317 0.0919286
R5426 VSS.n2012 VSS.n2011 0.0919286
R5427 VSS.n2026 VSS.n106 0.0919286
R5428 VSS.n2051 VSS.n2050 0.0919286
R5429 VSS.n2097 VSS.n65 0.0919286
R5430 VSS.n2134 VSS.n2133 0.0919286
R5431 VSS.n1908 VSS.n1907 0.0919286
R5432 VSS.n1922 VSS.n181 0.0919286
R5433 VSS.n1930 VSS.n1929 0.0919286
R5434 VSS.n1690 VSS.n1689 0.0919286
R5435 VSS.n1609 VSS.n1580 0.0919286
R5436 VSS.n1813 VSS.n1812 0.024
R5437 VSS.n1783 VSS.n1782 0.024
R5438 VSS.n780 VSS.n779 0.024
R5439 VSS.n750 VSS.n749 0.024
R5440 VSS.n887 VSS.n886 0.024
R5441 VSS.n949 VSS.n948 0.024
R5442 VSS.n1353 VSS.n1352 0.024
R5443 VSS.n1323 VSS.n1322 0.024
R5444 VSS.n1842 VSS.n1841 0.024
R5445 VSS.n1914 VSS.n1913 0.024
R5446 VSS.n1947 VSS.n1946 0.024
R5447 VSS.n2018 VSS.n2017 0.024
R5448 VSS.n1764 VSS.n1763 0.024
R5449 VSS.n1734 VSS.n1733 0.024
R5450 VSS.n1753 VSS.n1752 0.0228214
R5451 VSS.n1745 VSS.n1744 0.0228214
R5452 VSS.n1737 VSS.n1393 0.0228214
R5453 VSS.n223 VSS.n210 0.0228214
R5454 VSS.n1886 VSS.n1885 0.0228214
R5455 VSS.n1894 VSS.n188 0.0228214
R5456 VSS.n769 VSS.n768 0.0228214
R5457 VSS.n761 VSS.n760 0.0228214
R5458 VSS.n753 VSS.n408 0.0228214
R5459 VSS.n1802 VSS.n1801 0.0228214
R5460 VSS.n1794 VSS.n1793 0.0228214
R5461 VSS.n1786 VSS.n275 0.0228214
R5462 VSS.n692 VSS.n591 0.0228214
R5463 VSS.n1342 VSS.n1341 0.0228214
R5464 VSS.n1334 VSS.n1333 0.0228214
R5465 VSS.n1326 VSS.n1000 0.0228214
R5466 VSS.n915 VSS.n914 0.0228214
R5467 VSS.n836 VSS.n818 0.0228214
R5468 VSS.n945 VSS.n813 0.0228214
R5469 VSS.n1265 VSS.n1183 0.0228214
R5470 VSS.n146 VSS.n135 0.0228214
R5471 VSS.n1991 VSS.n1990 0.0228214
R5472 VSS.n1999 VSS.n113 0.0228214
R5473 VSS.n52 VSS.n36 0.0228214
R5474 VSS.n1674 VSS.n1673 0.0228214
R5475 VSS.n1760 VSS.n1371 0.0210357
R5476 VSS.n234 VSS.n227 0.0210357
R5477 VSS.n776 VSS.n386 0.0210357
R5478 VSS.n1809 VSS.n252 0.0210357
R5479 VSS.n711 VSS.n710 0.0210357
R5480 VSS.n604 VSS.n559 0.0210357
R5481 VSS.n603 VSS.n557 0.0210357
R5482 VSS.n1349 VSS.n978 0.0210357
R5483 VSS.n859 VSS.n858 0.0210357
R5484 VSS.n1284 VSS.n1283 0.0210357
R5485 VSS.n1196 VSS.n1151 0.0210357
R5486 VSS.n1195 VSS.n1149 0.0210357
R5487 VSS.n159 VSS.n151 0.0210357
R5488 VSS.n2095 VSS.n63 0.0210357
R5489 VSS.n2115 VSS.n2114 0.0210357
R5490 VSS.n2113 VSS.n55 0.0210357
R5491 VSS.n1692 VSS.n1543 0.0210357
R5492 VSS.n1681 VSS.n1550 0.0210357
R5493 VSS.n1680 VSS.n1552 0.0210357
R5494 VSS.n703 VSS.n559 0.0201429
R5495 VSS.n686 VSS.n685 0.0201429
R5496 VSS.n704 VSS.n557 0.0201429
R5497 VSS.n1276 VSS.n1151 0.0201429
R5498 VSS.n1259 VSS.n1258 0.0201429
R5499 VSS.n1277 VSS.n1149 0.0201429
R5500 VSS.n2114 VSS.n58 0.0201429
R5501 VSS.n2154 VSS.n2153 0.0201429
R5502 VSS.n2113 VSS.n2112 0.0201429
R5503 VSS.n1570 VSS.n1550 0.0201429
R5504 VSS.n1663 VSS.n1586 0.0201429
R5505 VSS.n1571 VSS.n1552 0.0201429
R5506 VSS.n721 VSS.n542 0.01925
R5507 VSS.n1294 VSS.n1134 0.01925
R5508 VSS.n2088 VSS.n83 0.01925
R5509 VSS.n1538 VSS.n1525 0.01925
R5510 VSS.n1384 VSS.n1377 0.0174643
R5511 VSS.n1746 VSS.n1384 0.0174643
R5512 VSS.n1750 VSS.n1380 0.0174643
R5513 VSS.n1747 VSS.n1380 0.0174643
R5514 VSS.n212 VSS.n204 0.0174643
R5515 VSS.n399 VSS.n392 0.0174643
R5516 VSS.n762 VSS.n399 0.0174643
R5517 VSS.n1795 VSS.n266 0.0174643
R5518 VSS.n1796 VSS.n264 0.0174643
R5519 VSS.n556 VSS.n550 0.0174643
R5520 VSS.n766 VSS.n395 0.0174643
R5521 VSS.n763 VSS.n395 0.0174643
R5522 VSS.n991 VSS.n984 0.0174643
R5523 VSS.n1335 VSS.n991 0.0174643
R5524 VSS.n925 VSS.n835 0.0174643
R5525 VSS.n924 VSS.n923 0.0174643
R5526 VSS.n1148 VSS.n1142 0.0174643
R5527 VSS.n1339 VSS.n987 0.0174643
R5528 VSS.n1336 VSS.n987 0.0174643
R5529 VSS.n1983 VSS.n1982 0.0174643
R5530 VSS.n1982 VSS.n129 0.0174643
R5531 VSS.n1984 VSS.n134 0.0174643
R5532 VSS.n134 VSS.n130 0.0174643
R5533 VSS.n62 VSS.n59 0.0174643
R5534 VSS.n211 VSS.n205 0.0174643
R5535 VSS.n1562 VSS.n1555 0.0174643
R5536 VSS.n1436 VSS.n1435 0.0165714
R5537 VSS.n1739 VSS.n1738 0.0165714
R5538 VSS.n1485 VSS.n1483 0.0165714
R5539 VSS.n1878 VSS.n1877 0.0165714
R5540 VSS.n297 VSS.n258 0.0165714
R5541 VSS.n319 VSS.n318 0.0165714
R5542 VSS.n1808 VSS.n1807 0.0165714
R5543 VSS.n1807 VSS.n253 0.0165714
R5544 VSS.n1799 VSS.n261 0.0165714
R5545 VSS.n367 VSS.n365 0.0165714
R5546 VSS.n705 VSS.n556 0.0165714
R5547 VSS.n602 VSS.n600 0.0165714
R5548 VSS.n598 VSS.n596 0.0165714
R5549 VSS.n451 VSS.n450 0.0165714
R5550 VSS.n755 VSS.n754 0.0165714
R5551 VSS.n500 VSS.n498 0.0165714
R5552 VSS.n926 VSS.n833 0.0165714
R5553 VSS.n880 VSS.n879 0.0165714
R5554 VSS.n908 VSS.n843 0.0165714
R5555 VSS.n908 VSS.n907 0.0165714
R5556 VSS.n917 VSS.n834 0.0165714
R5557 VSS.n956 VSS.n955 0.0165714
R5558 VSS.n1278 VSS.n1148 0.0165714
R5559 VSS.n1194 VSS.n1192 0.0165714
R5560 VSS.n1190 VSS.n1188 0.0165714
R5561 VSS.n1043 VSS.n1042 0.0165714
R5562 VSS.n1328 VSS.n1327 0.0165714
R5563 VSS.n1092 VSS.n1090 0.0165714
R5564 VSS.n1940 VSS.n1939 0.0165714
R5565 VSS.n1996 VSS.n126 0.0165714
R5566 VSS.n2023 VSS.n109 0.0165714
R5567 VSS.n2111 VSS.n59 0.0165714
R5568 VSS.n2122 VSS.n2121 0.0165714
R5569 VSS.n2128 VSS.n51 0.0165714
R5570 VSS.n1835 VSS.n1834 0.0165714
R5571 VSS.n1858 VSS.n226 0.0165714
R5572 VSS.n1858 VSS.n1857 0.0165714
R5573 VSS.n1879 VSS.n209 0.0165714
R5574 VSS.n1919 VSS.n184 0.0165714
R5575 VSS.n1572 VSS.n1555 0.0165714
R5576 VSS.n1679 VSS.n1553 0.0165714
R5577 VSS.n1605 VSS.n1576 0.0165714
R5578 VSS.n1759 VSS.n1758 0.0156786
R5579 VSS.n1788 VSS.n1787 0.0156786
R5580 VSS.n537 VSS.n535 0.0156786
R5581 VSS.n726 VSS.n520 0.0156786
R5582 VSS.n722 VSS.n520 0.0156786
R5583 VSS.n687 VSS.n620 0.0156786
R5584 VSS.n627 VSS.n620 0.0156786
R5585 VSS.n775 VSS.n774 0.0156786
R5586 VSS.n944 VSS.n943 0.0156786
R5587 VSS.n1129 VSS.n1127 0.0156786
R5588 VSS.n1299 VSS.n1112 0.0156786
R5589 VSS.n1295 VSS.n1112 0.0156786
R5590 VSS.n1260 VSS.n1212 0.0156786
R5591 VSS.n1238 VSS.n1212 0.0156786
R5592 VSS.n1348 VSS.n1347 0.0156786
R5593 VSS.n1963 VSS.n149 0.0156786
R5594 VSS.n2061 VSS.n2059 0.0156786
R5595 VSS.n2069 VSS.n81 0.0156786
R5596 VSS.n2089 VSS.n81 0.0156786
R5597 VSS.n2152 VSS.n32 0.0156786
R5598 VSS.n32 VSS.n27 0.0156786
R5599 VSS.n1891 VSS.n201 0.0156786
R5600 VSS.n1521 VSS.n1519 0.0156786
R5601 VSS.n1710 VSS.n1505 0.0156786
R5602 VSS.n1539 VSS.n1505 0.0156786
R5603 VSS.n1662 VSS.n1587 0.0156786
R5604 VSS.n1658 VSS.n1587 0.0156786
R5605 VSS.n1806 VSS.n1805 0.0152714
R5606 VSS.n1790 VSS.n1789 0.0152714
R5607 VSS.n773 VSS.n772 0.0152714
R5608 VSS.n757 VSS.n756 0.0152714
R5609 VSS.n707 VSS.n706 0.0152714
R5610 VSS.n601 VSS.n595 0.0152714
R5611 VSS.n910 VSS.n909 0.0152714
R5612 VSS.n942 VSS.n941 0.0152714
R5613 VSS.n1346 VSS.n1345 0.0152714
R5614 VSS.n1330 VSS.n1329 0.0152714
R5615 VSS.n1280 VSS.n1279 0.0152714
R5616 VSS.n1193 VSS.n1187 0.0152714
R5617 VSS.n1863 VSS.n1859 0.0152714
R5618 VSS.n1890 VSS.n1889 0.0152714
R5619 VSS.n1968 VSS.n1964 0.0152714
R5620 VSS.n1995 VSS.n1994 0.0152714
R5621 VSS.n2110 VSS.n2109 0.0152714
R5622 VSS.n2126 VSS.n2123 0.0152714
R5623 VSS.n1757 VSS.n1756 0.0152714
R5624 VSS.n1741 VSS.n1740 0.0152714
R5625 VSS.n1573 VSS.n1554 0.0152714
R5626 VSS.n1678 VSS.n1677 0.0152714
R5627 VSS.n552 VSS.n549 0.0147857
R5628 VSS.n615 VSS.n593 0.0147857
R5629 VSS.n1144 VSS.n1141 0.0147857
R5630 VSS.n1207 VSS.n1185 0.0147857
R5631 VSS.n79 VSS.n61 0.0147857
R5632 VSS.n2124 VSS.n34 0.0147857
R5633 VSS.n1560 VSS.n1534 0.0147857
R5634 VSS.n1589 VSS.n1588 0.0147857
R5635 VSS.n636 VSS.n629 0.0138929
R5636 VSS.n1241 VSS.n1240 0.0138929
R5637 VSS.n2164 VSS.n21 0.0138929
R5638 VSS.n1636 VSS.n1623 0.0138929
R5639 VSS.n1798 VSS.n1797 0.0132571
R5640 VSS.n765 VSS.n764 0.0132571
R5641 VSS.n725 VSS.n539 0.0132571
R5642 VSS.n723 VSS.n540 0.0132571
R5643 VSS.n689 VSS.n688 0.0132571
R5644 VSS.n673 VSS.n631 0.0132571
R5645 VSS.n922 VSS.n918 0.0132571
R5646 VSS.n1338 VSS.n1337 0.0132571
R5647 VSS.n1298 VSS.n1131 0.0132571
R5648 VSS.n1296 VSS.n1132 0.0132571
R5649 VSS.n1262 VSS.n1261 0.0132571
R5650 VSS.n1246 VSS.n1244 0.0132571
R5651 VSS.n1881 VSS.n1880 0.0132571
R5652 VSS.n1986 VSS.n1985 0.0132571
R5653 VSS.n2064 VSS.n2063 0.0132571
R5654 VSS.n2092 VSS.n2090 0.0132571
R5655 VSS.n2151 VSS.n2148 0.0132571
R5656 VSS.n2149 VSS.n24 0.0132571
R5657 VSS.n1749 VSS.n1748 0.0132571
R5658 VSS.n1524 VSS.n1523 0.0132571
R5659 VSS.n1541 VSS.n1540 0.0132571
R5660 VSS.n1661 VSS.n1591 0.0132571
R5661 VSS.n1659 VSS.n1592 0.0132571
R5662 VSS.n1486 VSS.n1408 0.013
R5663 VSS.n1731 VSS.n1730 0.013
R5664 VSS.n1485 VSS.n1484 0.013
R5665 VSS.n1839 VSS.n1831 0.013
R5666 VSS.n1837 VSS.n1833 0.013
R5667 VSS.n501 VSS.n423 0.013
R5668 VSS.n747 VSS.n746 0.013
R5669 VSS.n1817 VSS.n245 0.013
R5670 VSS.n317 VSS.n315 0.013
R5671 VSS.n318 VSS.n312 0.013
R5672 VSS.n500 VSS.n499 0.013
R5673 VSS.n1093 VSS.n1015 0.013
R5674 VSS.n1320 VSS.n1319 0.013
R5675 VSS.n884 VSS.n876 0.013
R5676 VSS.n882 VSS.n878 0.013
R5677 VSS.n881 VSS.n880 0.013
R5678 VSS.n1092 VSS.n1091 0.013
R5679 VSS.n2024 VSS.n108 0.013
R5680 VSS.n2052 VSS.n100 0.013
R5681 VSS.n2023 VSS.n2022 0.013
R5682 VSS.n1836 VSS.n1835 0.013
R5683 VSS.n1768 VSS.n1364 0.0121071
R5684 VSS.n1434 VSS.n1432 0.0121071
R5685 VSS.n1435 VSS.n1429 0.0121071
R5686 VSS.n1409 VSS.n1395 0.0121071
R5687 VSS.n1846 VSS.n1845 0.0121071
R5688 VSS.n1920 VSS.n183 0.0121071
R5689 VSS.n1931 VSS.n175 0.0121071
R5690 VSS.n784 VSS.n378 0.0121071
R5691 VSS.n449 VSS.n447 0.0121071
R5692 VSS.n321 VSS.n251 0.0121071
R5693 VSS.n368 VSS.n290 0.0121071
R5694 VSS.n1780 VSS.n1779 0.0121071
R5695 VSS.n320 VSS.n249 0.0121071
R5696 VSS.n367 VSS.n366 0.0121071
R5697 VSS.n535 VSS.n526 0.0121071
R5698 VSS.n450 VSS.n444 0.0121071
R5699 VSS.n424 VSS.n410 0.0121071
R5700 VSS.n1357 VSS.n792 0.0121071
R5701 VSS.n1041 VSS.n1039 0.0121071
R5702 VSS.n891 VSS.n890 0.0121071
R5703 VSS.n954 VSS.n953 0.0121071
R5704 VSS.n969 VSS.n795 0.0121071
R5705 VSS.n889 VSS.n857 0.0121071
R5706 VSS.n955 VSS.n805 0.0121071
R5707 VSS.n1127 VSS.n1118 0.0121071
R5708 VSS.n1042 VSS.n1036 0.0121071
R5709 VSS.n1016 VSS.n1002 0.0121071
R5710 VSS.n1944 VSS.n1936 0.0121071
R5711 VSS.n1942 VSS.n1938 0.0121071
R5712 VSS.n1941 VSS.n1940 0.0121071
R5713 VSS.n115 VSS.n112 0.0121071
R5714 VSS.n2059 VSS.n96 0.0121071
R5715 VSS.n1844 VSS.n233 0.0121071
R5716 VSS.n1919 VSS.n1918 0.0121071
R5717 VSS.n1519 VSS.n1510 0.0121071
R5718 VSS.n1434 VSS.n1433 0.0112143
R5719 VSS.n1438 VSS.n1370 0.0112143
R5720 VSS.n1410 VSS.n1394 0.0112143
R5721 VSS.n1437 VSS.n1368 0.0112143
R5722 VSS.n1921 VSS.n1920 0.0112143
R5723 VSS.n449 VSS.n448 0.0112143
R5724 VSS.n453 VSS.n385 0.0112143
R5725 VSS.n425 VSS.n409 0.0112143
R5726 VSS.n369 VSS.n368 0.0112143
R5727 VSS.n291 VSS.n277 0.0112143
R5728 VSS.n581 VSS.n548 0.0112143
R5729 VSS.n611 VSS.n610 0.0112143
R5730 VSS.n649 VSS.n621 0.0112143
R5731 VSS.n637 VSS.n636 0.0112143
R5732 VSS.n648 VSS.n619 0.0112143
R5733 VSS.n452 VSS.n383 0.0112143
R5734 VSS.n1041 VSS.n1040 0.0112143
R5735 VSS.n1045 VSS.n977 0.0112143
R5736 VSS.n1017 VSS.n1001 0.0112143
R5737 VSS.n954 VSS.n810 0.0112143
R5738 VSS.n957 VSS.n804 0.0112143
R5739 VSS.n1173 VSS.n1140 0.0112143
R5740 VSS.n1203 VSS.n1202 0.0112143
R5741 VSS.n1226 VSS.n1213 0.0112143
R5742 VSS.n1241 VSS.n4 0.0112143
R5743 VSS.n1225 VSS.n1211 0.0112143
R5744 VSS.n1044 VSS.n975 0.0112143
R5745 VSS.n1938 VSS.n1937 0.0112143
R5746 VSS.n1951 VSS.n1950 0.0112143
R5747 VSS.n2014 VSS.n2013 0.0112143
R5748 VSS.n1949 VSS.n158 0.0112143
R5749 VSS.n2106 VSS.n2105 0.0112143
R5750 VSS.n2130 VSS.n2129 0.0112143
R5751 VSS.n42 VSS.n30 0.0112143
R5752 VSS.n2175 VSS.n21 0.0112143
R5753 VSS.n41 VSS.n31 0.0112143
R5754 VSS.n190 VSS.n187 0.0112143
R5755 VSS.n1564 VSS.n1563 0.0112143
R5756 VSS.n1607 VSS.n1578 0.0112143
R5757 VSS.n1665 VSS.n1664 0.0112143
R5758 VSS.n1646 VSS.n1623 0.0112143
R5759 VSS.n1666 VSS.n1584 0.0112143
R5760 VSS.n1438 VSS.n1428 0.0103214
R5761 VSS.n1761 VSS.n1760 0.0103214
R5762 VSS.n1754 VSS.n1376 0.0103214
R5763 VSS.n1465 VSS.n1385 0.0103214
R5764 VSS.n1487 VSS.n1486 0.0103214
R5765 VSS.n1437 VSS.n1436 0.0103214
R5766 VSS.n1755 VSS.n1374 0.0103214
R5767 VSS.n1751 VSS.n1379 0.0103214
R5768 VSS.n1742 VSS.n1388 0.0103214
R5769 VSS.n1469 VSS.n1391 0.0103214
R5770 VSS.n1833 VSS.n1832 0.0103214
R5771 VSS.n1866 VSS.n221 0.0103214
R5772 VSS.n1887 VSS.n198 0.0103214
R5773 VSS.n1911 VSS.n188 0.0103214
R5774 VSS.n1910 VSS.n1909 0.0103214
R5775 VSS.n191 VSS.n189 0.0103214
R5776 VSS.n453 VSS.n443 0.0103214
R5777 VSS.n777 VSS.n776 0.0103214
R5778 VSS.n770 VSS.n391 0.0103214
R5779 VSS.n480 VSS.n400 0.0103214
R5780 VSS.n502 VSS.n501 0.0103214
R5781 VSS.n317 VSS.n316 0.0103214
R5782 VSS.n1803 VSS.n257 0.0103214
R5783 VSS.n346 VSS.n267 0.0103214
R5784 VSS.n1786 VSS.n1785 0.0103214
R5785 VSS.n292 VSS.n276 0.0103214
R5786 VSS.n364 VSS.n363 0.0103214
R5787 VSS.n1804 VSS.n255 0.0103214
R5788 VSS.n268 VSS.n265 0.0103214
R5789 VSS.n1791 VSS.n270 0.0103214
R5790 VSS.n365 VSS.n291 0.0103214
R5791 VSS.n729 VSS.n728 0.0103214
R5792 VSS.n566 VSS.n542 0.0103214
R5793 VSS.n720 VSS.n719 0.0103214
R5794 VSS.n727 VSS.n518 0.0103214
R5795 VSS.n718 VSS.n541 0.0103214
R5796 VSS.n452 VSS.n451 0.0103214
R5797 VSS.n771 VSS.n389 0.0103214
R5798 VSS.n767 VSS.n394 0.0103214
R5799 VSS.n758 VSS.n403 0.0103214
R5800 VSS.n484 VSS.n406 0.0103214
R5801 VSS.n1045 VSS.n1035 0.0103214
R5802 VSS.n1350 VSS.n1349 0.0103214
R5803 VSS.n1343 VSS.n983 0.0103214
R5804 VSS.n1072 VSS.n992 0.0103214
R5805 VSS.n1094 VSS.n1093 0.0103214
R5806 VSS.n878 VSS.n877 0.0103214
R5807 VSS.n847 VSS.n840 0.0103214
R5808 VSS.n939 VSS.n938 0.0103214
R5809 VSS.n946 VSS.n945 0.0103214
R5810 VSS.n959 VSS.n802 0.0103214
R5811 VSS.n958 VSS.n803 0.0103214
R5812 VSS.n846 VSS.n841 0.0103214
R5813 VSS.n920 VSS.n837 0.0103214
R5814 VSS.n940 VSS.n817 0.0103214
R5815 VSS.n957 VSS.n956 0.0103214
R5816 VSS.n1302 VSS.n1301 0.0103214
R5817 VSS.n1158 VSS.n1134 0.0103214
R5818 VSS.n1293 VSS.n1292 0.0103214
R5819 VSS.n1300 VSS.n1110 0.0103214
R5820 VSS.n1291 VSS.n1133 0.0103214
R5821 VSS.n1044 VSS.n1043 0.0103214
R5822 VSS.n1344 VSS.n981 0.0103214
R5823 VSS.n1340 VSS.n986 0.0103214
R5824 VSS.n1331 VSS.n995 0.0103214
R5825 VSS.n1076 VSS.n998 0.0103214
R5826 VSS.n1951 VSS.n157 0.0103214
R5827 VSS.n160 VSS.n159 0.0103214
R5828 VSS.n1971 VSS.n144 0.0103214
R5829 VSS.n1992 VSS.n123 0.0103214
R5830 VSS.n2025 VSS.n2024 0.0103214
R5831 VSS.n1939 VSS.n158 0.0103214
R5832 VSS.n1970 VSS.n1969 0.0103214
R5833 VSS.n1965 VSS.n133 0.0103214
R5834 VSS.n1993 VSS.n125 0.0103214
R5835 VSS.n2001 VSS.n2000 0.0103214
R5836 VSS.n2072 VSS.n91 0.0103214
R5837 VSS.n2067 VSS.n83 0.0103214
R5838 VSS.n2087 VSS.n2086 0.0103214
R5839 VSS.n2071 VSS.n2070 0.0103214
R5840 VSS.n2085 VSS.n82 0.0103214
R5841 VSS.n1865 VSS.n1864 0.0103214
R5842 VSS.n1884 VSS.n1883 0.0103214
R5843 VSS.n1888 VSS.n200 0.0103214
R5844 VSS.n190 VSS.n184 0.0103214
R5845 VSS.n1713 VSS.n1503 0.0103214
R5846 VSS.n1708 VSS.n1525 0.0103214
R5847 VSS.n1537 VSS.n1531 0.0103214
R5848 VSS.n1712 VSS.n1711 0.0103214
R5849 VSS.n1536 VSS.n1533 0.0103214
R5850 VSS.n706 VSS.n555 0.00956429
R5851 VSS.n601 VSS.n555 0.00956429
R5852 VSS.n1279 VSS.n1147 0.00956429
R5853 VSS.n1193 VSS.n1147 0.00956429
R5854 VSS.n2110 VSS.n54 0.00956429
R5855 VSS.n2123 VSS.n54 0.00956429
R5856 VSS.n1574 VSS.n1573 0.00956429
R5857 VSS.n1678 VSS.n1574 0.00956429
R5858 VSS.n1432 VSS.n1431 0.00942857
R5859 VSS.n1737 VSS.n1736 0.00942857
R5860 VSS.n1482 VSS.n1481 0.00942857
R5861 VSS.n1430 VSS.n1429 0.00942857
R5862 VSS.n1443 VSS.n1372 0.00942857
R5863 VSS.n1386 VSS.n1383 0.00942857
R5864 VSS.n1483 VSS.n1409 0.00942857
R5865 VSS.n1846 VSS.n232 0.00942857
R5866 VSS.n235 VSS.n234 0.00942857
R5867 VSS.n1916 VSS.n183 0.00942857
R5868 VSS.n447 VSS.n446 0.00942857
R5869 VSS.n753 VSS.n752 0.00942857
R5870 VSS.n497 VSS.n496 0.00942857
R5871 VSS.n321 VSS.n311 0.00942857
R5872 VSS.n1810 VSS.n1809 0.00942857
R5873 VSS.n290 VSS.n281 0.00942857
R5874 VSS.n320 VSS.n319 0.00942857
R5875 VSS.n1800 VSS.n260 0.00942857
R5876 VSS.n350 VSS.n273 0.00942857
R5877 VSS.n366 VSS.n279 0.00942857
R5878 VSS.n580 VSS.n579 0.00942857
R5879 VSS.n703 VSS.n558 0.00942857
R5880 VSS.n606 VSS.n597 0.00942857
R5881 VSS.n685 VSS.n622 0.00942857
R5882 VSS.n681 VSS.n626 0.00942857
R5883 VSS.n680 VSS.n679 0.00942857
R5884 VSS.n445 VSS.n444 0.00942857
R5885 VSS.n458 VSS.n387 0.00942857
R5886 VSS.n401 VSS.n398 0.00942857
R5887 VSS.n498 VSS.n424 0.00942857
R5888 VSS.n1039 VSS.n1038 0.00942857
R5889 VSS.n1326 VSS.n1325 0.00942857
R5890 VSS.n1089 VSS.n1088 0.00942857
R5891 VSS.n891 VSS.n856 0.00942857
R5892 VSS.n860 VSS.n859 0.00942857
R5893 VSS.n953 VSS.n952 0.00942857
R5894 VSS.n879 VSS.n857 0.00942857
R5895 VSS.n916 VSS.n839 0.00942857
R5896 VSS.n824 VSS.n814 0.00942857
R5897 VSS.n951 VSS.n805 0.00942857
R5898 VSS.n1172 VSS.n1171 0.00942857
R5899 VSS.n1276 VSS.n1150 0.00942857
R5900 VSS.n1198 VSS.n1189 0.00942857
R5901 VSS.n1258 VSS.n1214 0.00942857
R5902 VSS.n1254 VSS.n1237 0.00942857
R5903 VSS.n1253 VSS.n1252 0.00942857
R5904 VSS.n1037 VSS.n1036 0.00942857
R5905 VSS.n1050 VSS.n979 0.00942857
R5906 VSS.n993 VSS.n990 0.00942857
R5907 VSS.n1090 VSS.n1016 0.00942857
R5908 VSS.n1943 VSS.n1942 0.00942857
R5909 VSS.n2015 VSS.n113 0.00942857
R5910 VSS.n116 VSS.n114 0.00942857
R5911 VSS.n1941 VSS.n164 0.00942857
R5912 VSS.n1962 VSS.n150 0.00942857
R5913 VSS.n1989 VSS.n1988 0.00942857
R5914 VSS.n115 VSS.n109 0.00942857
R5915 VSS.n69 VSS.n64 0.00942857
R5916 VSS.n68 VSS.n58 0.00942857
R5917 VSS.n2120 VSS.n2119 0.00942857
R5918 VSS.n2155 VSS.n2154 0.00942857
R5919 VSS.n2158 VSS.n26 0.00942857
R5920 VSS.n2160 VSS.n2159 0.00942857
R5921 VSS.n1834 VSS.n233 0.00942857
R5922 VSS.n1860 VSS.n208 0.00942857
R5923 VSS.n1896 VSS.n1895 0.00942857
R5924 VSS.n1918 VSS.n1917 0.00942857
R5925 VSS.n1565 VSS.n1556 0.00942857
R5926 VSS.n1570 VSS.n1569 0.00942857
R5927 VSS.n1604 VSS.n1603 0.00942857
R5928 VSS.n1594 VSS.n1586 0.00942857
R5929 VSS.n1656 VSS.n1595 0.00942857
R5930 VSS.n1632 VSS.n1593 0.00942857
R5931 VSS.n1408 VSS.n1399 0.00853571
R5932 VSS.n1484 VSS.n1397 0.00853571
R5933 VSS.n1401 VSS.n1398 0.00853571
R5934 VSS.n1838 VSS.n1837 0.00853571
R5935 VSS.n1856 VSS.n1855 0.00853571
R5936 VSS.n423 VSS.n414 0.00853571
R5937 VSS.n315 VSS.n314 0.00853571
R5938 VSS.n326 VSS.n325 0.00853571
R5939 VSS.n1816 VSS.n1815 0.00853571
R5940 VSS.n313 VSS.n312 0.00853571
R5941 VSS.n323 VSS.n255 0.00853571
R5942 VSS.n711 VSS.n545 0.00853571
R5943 VSS.n605 VSS.n604 0.00853571
R5944 VSS.n691 VSS.n592 0.00853571
R5945 VSS.n533 VSS.n529 0.00853571
R5946 VSS.n538 VSS.n522 0.00853571
R5947 VSS.n552 VSS.n551 0.00853571
R5948 VSS.n708 VSS.n549 0.00853571
R5949 VSS.n690 VSS.n593 0.00853571
R5950 VSS.n690 VSS.n594 0.00853571
R5951 VSS.n674 VSS.n630 0.00853571
R5952 VSS.n634 VSS.n630 0.00853571
R5953 VSS.n670 VSS.n669 0.00853571
R5954 VSS.n499 VSS.n412 0.00853571
R5955 VSS.n416 VSS.n413 0.00853571
R5956 VSS.n1015 VSS.n1006 0.00853571
R5957 VSS.n883 VSS.n882 0.00853571
R5958 VSS.n906 VSS.n845 0.00853571
R5959 VSS.n875 VSS.n863 0.00853571
R5960 VSS.n881 VSS.n864 0.00853571
R5961 VSS.n846 VSS.n844 0.00853571
R5962 VSS.n1284 VSS.n1137 0.00853571
R5963 VSS.n1197 VSS.n1196 0.00853571
R5964 VSS.n1264 VSS.n1184 0.00853571
R5965 VSS.n1125 VSS.n1121 0.00853571
R5966 VSS.n1130 VSS.n1114 0.00853571
R5967 VSS.n1144 VSS.n1143 0.00853571
R5968 VSS.n1281 VSS.n1141 0.00853571
R5969 VSS.n1263 VSS.n1185 0.00853571
R5970 VSS.n1263 VSS.n1186 0.00853571
R5971 VSS.n1247 VSS.n1243 0.00853571
R5972 VSS.n1243 VSS.n1242 0.00853571
R5973 VSS.n2196 VSS.n2 0.00853571
R5974 VSS.n1091 VSS.n1004 0.00853571
R5975 VSS.n1008 VSS.n1005 0.00853571
R5976 VSS.n2020 VSS.n108 0.00853571
R5977 VSS.n2022 VSS.n2021 0.00853571
R5978 VSS.n2053 VSS.n99 0.00853571
R5979 VSS.n2095 VSS.n2094 0.00853571
R5980 VSS.n2115 VSS.n56 0.00853571
R5981 VSS.n2146 VSS.n2145 0.00853571
R5982 VSS.n2057 VSS.n97 0.00853571
R5983 VSS.n2062 VSS.n94 0.00853571
R5984 VSS.n2093 VSS.n79 0.00853571
R5985 VSS.n2108 VSS.n61 0.00853571
R5986 VSS.n2147 VSS.n34 0.00853571
R5987 VSS.n2147 VSS.n35 0.00853571
R5988 VSS.n2168 VSS.n2166 0.00853571
R5989 VSS.n2168 VSS.n2167 0.00853571
R5990 VSS.n2173 VSS.n23 0.00853571
R5991 VSS.n1830 VSS.n238 0.00853571
R5992 VSS.n1836 VSS.n239 0.00853571
R5993 VSS.n1865 VSS.n222 0.00853571
R5994 VSS.n1693 VSS.n1692 0.00853571
R5995 VSS.n1681 VSS.n1551 0.00853571
R5996 VSS.n1669 VSS.n1579 0.00853571
R5997 VSS.n1517 VSS.n1513 0.00853571
R5998 VSS.n1522 VSS.n1507 0.00853571
R5999 VSS.n1694 VSS.n1534 0.00853571
R6000 VSS.n1561 VSS.n1560 0.00853571
R6001 VSS.n1589 VSS.n1583 0.00853571
R6002 VSS.n1668 VSS.n1583 0.00853571
R6003 VSS.n1640 VSS.n1638 0.00853571
R6004 VSS.n1640 VSS.n1639 0.00853571
R6005 VSS.n1644 VSS.n1625 0.00853571
R6006 VSS.n1814 VSS.n246 0.00822143
R6007 VSS.n1806 VSS.n248 0.00822143
R6008 VSS.n1789 VSS.n272 0.00822143
R6009 VSS.n379 VSS.n278 0.00822143
R6010 VSS.n781 VSS.n380 0.00822143
R6011 VSS.n773 VSS.n382 0.00822143
R6012 VSS.n756 VSS.n405 0.00822143
R6013 VSS.n530 VSS.n411 0.00822143
R6014 VSS.n874 VSS.n862 0.00822143
R6015 VSS.n909 VSS.n842 0.00822143
R6016 VSS.n942 VSS.n811 0.00822143
R6017 VSS.n971 VSS.n793 0.00822143
R6018 VSS.n1354 VSS.n972 0.00822143
R6019 VSS.n1346 VSS.n974 0.00822143
R6020 VSS.n1329 VSS.n997 0.00822143
R6021 VSS.n1122 VSS.n1003 0.00822143
R6022 VSS.n1829 VSS.n237 0.00822143
R6023 VSS.n1859 VSS.n225 0.00822143
R6024 VSS.n1890 VSS.n185 0.00822143
R6025 VSS.n1933 VSS.n173 0.00822143
R6026 VSS.n1934 VSS.n162 0.00822143
R6027 VSS.n1964 VSS.n148 0.00822143
R6028 VSS.n1995 VSS.n110 0.00822143
R6029 VSS.n2054 VSS.n98 0.00822143
R6030 VSS.n1765 VSS.n1365 0.00822143
R6031 VSS.n1757 VSS.n1367 0.00822143
R6032 VSS.n1740 VSS.n1390 0.00822143
R6033 VSS.n1514 VSS.n1396 0.00822143
R6034 VSS.n1445 VSS.n1444 0.00764286
R6035 VSS.n1468 VSS.n1467 0.00764286
R6036 VSS.n1767 VSS.n1766 0.00764286
R6037 VSS.n1758 VSS.n1372 0.00764286
R6038 VSS.n1442 VSS.n1374 0.00764286
R6039 VSS.n1379 VSS.n1378 0.00764286
R6040 VSS.n1387 VSS.n1386 0.00764286
R6041 VSS.n1470 VSS.n1388 0.00764286
R6042 VSS.n1898 VSS.n199 0.00764286
R6043 VSS.n460 VSS.n459 0.00764286
R6044 VSS.n483 VSS.n482 0.00764286
R6045 VSS.n352 VSS.n349 0.00764286
R6046 VSS.n260 VSS.n259 0.00764286
R6047 VSS.n269 VSS.n268 0.00764286
R6048 VSS.n351 VSS.n350 0.00764286
R6049 VSS.n1788 VSS.n273 0.00764286
R6050 VSS.n283 VSS.n280 0.00764286
R6051 VSS.n537 VSS.n536 0.00764286
R6052 VSS.n729 VSS.n517 0.00764286
R6053 VSS.n715 VSS.n545 0.00764286
R6054 VSS.n692 VSS.n691 0.00764286
R6055 VSS.n677 VSS.n626 0.00764286
R6056 VSS.n677 VSS.n676 0.00764286
R6057 VSS.n534 VSS.n533 0.00764286
R6058 VSS.n534 VSS.n522 0.00764286
R6059 VSS.n538 VSS.n524 0.00764286
R6060 VSS.n523 VSS.n518 0.00764286
R6061 VSS.n718 VSS.n717 0.00764286
R6062 VSS.n551 VSS.n544 0.00764286
R6063 VSS.n615 VSS.n614 0.00764286
R6064 VSS.n648 VSS.n647 0.00764286
R6065 VSS.n679 VSS.n678 0.00764286
R6066 VSS.n678 VSS.n628 0.00764286
R6067 VSS.n783 VSS.n782 0.00764286
R6068 VSS.n774 VSS.n387 0.00764286
R6069 VSS.n457 VSS.n389 0.00764286
R6070 VSS.n394 VSS.n393 0.00764286
R6071 VSS.n402 VSS.n401 0.00764286
R6072 VSS.n485 VSS.n403 0.00764286
R6073 VSS.n1052 VSS.n1051 0.00764286
R6074 VSS.n1075 VSS.n1074 0.00764286
R6075 VSS.n825 VSS.n819 0.00764286
R6076 VSS.n912 VSS.n839 0.00764286
R6077 VSS.n920 VSS.n919 0.00764286
R6078 VSS.n824 VSS.n823 0.00764286
R6079 VSS.n943 VSS.n814 0.00764286
R6080 VSS.n970 VSS.n794 0.00764286
R6081 VSS.n1129 VSS.n1128 0.00764286
R6082 VSS.n1302 VSS.n1109 0.00764286
R6083 VSS.n1288 VSS.n1137 0.00764286
R6084 VSS.n1265 VSS.n1264 0.00764286
R6085 VSS.n1250 VSS.n1237 0.00764286
R6086 VSS.n1250 VSS.n1249 0.00764286
R6087 VSS.n1126 VSS.n1125 0.00764286
R6088 VSS.n1126 VSS.n1114 0.00764286
R6089 VSS.n1130 VSS.n1116 0.00764286
R6090 VSS.n1115 VSS.n1110 0.00764286
R6091 VSS.n1291 VSS.n1290 0.00764286
R6092 VSS.n1143 VSS.n1136 0.00764286
R6093 VSS.n1207 VSS.n1206 0.00764286
R6094 VSS.n1225 VSS.n1224 0.00764286
R6095 VSS.n1252 VSS.n1251 0.00764286
R6096 VSS.n1251 VSS.n1239 0.00764286
R6097 VSS.n1356 VSS.n1355 0.00764286
R6098 VSS.n1347 VSS.n979 0.00764286
R6099 VSS.n1049 VSS.n981 0.00764286
R6100 VSS.n986 VSS.n985 0.00764286
R6101 VSS.n994 VSS.n993 0.00764286
R6102 VSS.n1077 VSS.n995 0.00764286
R6103 VSS.n1960 VSS.n152 0.00764286
R6104 VSS.n1998 VSS.n124 0.00764286
R6105 VSS.n1935 VSS.n163 0.00764286
R6106 VSS.n1963 VSS.n1962 0.00764286
R6107 VSS.n1970 VSS.n145 0.00764286
R6108 VSS.n1966 VSS.n1965 0.00764286
R6109 VSS.n1988 VSS.n131 0.00764286
R6110 VSS.n2002 VSS.n125 0.00764286
R6111 VSS.n2061 VSS.n2060 0.00764286
R6112 VSS.n2072 VSS.n90 0.00764286
R6113 VSS.n2094 VSS.n77 0.00764286
R6114 VSS.n2146 VSS.n36 0.00764286
R6115 VSS.n2162 VSS.n26 0.00764286
R6116 VSS.n2163 VSS.n2162 0.00764286
R6117 VSS.n2058 VSS.n2057 0.00764286
R6118 VSS.n2058 VSS.n94 0.00764286
R6119 VSS.n2062 VSS.n95 0.00764286
R6120 VSS.n2071 VSS.n92 0.00764286
R6121 VSS.n2085 VSS.n2084 0.00764286
R6122 VSS.n2093 VSS.n78 0.00764286
R6123 VSS.n2124 VSS.n53 0.00764286
R6124 VSS.n41 VSS.n40 0.00764286
R6125 VSS.n2161 VSS.n2160 0.00764286
R6126 VSS.n2161 VSS.n25 0.00764286
R6127 VSS.n1861 VSS.n1860 0.00764286
R6128 VSS.n1883 VSS.n206 0.00764286
R6129 VSS.n1897 VSS.n1896 0.00764286
R6130 VSS.n1895 VSS.n1891 0.00764286
R6131 VSS.n1932 VSS.n174 0.00764286
R6132 VSS.n1521 VSS.n1520 0.00764286
R6133 VSS.n1713 VSS.n1502 0.00764286
R6134 VSS.n1693 VSS.n1532 0.00764286
R6135 VSS.n1673 VSS.n1579 0.00764286
R6136 VSS.n1634 VSS.n1595 0.00764286
R6137 VSS.n1635 VSS.n1634 0.00764286
R6138 VSS.n1518 VSS.n1517 0.00764286
R6139 VSS.n1518 VSS.n1507 0.00764286
R6140 VSS.n1522 VSS.n1508 0.00764286
R6141 VSS.n1712 VSS.n1504 0.00764286
R6142 VSS.n1696 VSS.n1533 0.00764286
R6143 VSS.n1695 VSS.n1694 0.00764286
R6144 VSS.n1588 VSS.n1577 0.00764286
R6145 VSS.n1667 VSS.n1666 0.00764286
R6146 VSS.n1633 VSS.n1632 0.00764286
R6147 VSS.n1633 VSS.n1631 0.00764286
R6148 VSS.n1444 VSS.n1441 0.00675
R6149 VSS.n1754 VSS.n1753 0.00675
R6150 VSS.n1471 VSS.n1468 0.00675
R6151 VSS.n1443 VSS.n1442 0.00675
R6152 VSS.n1755 VSS.n1375 0.00675
R6153 VSS.n1743 VSS.n1387 0.00675
R6154 VSS.n1470 VSS.n1469 0.00675
R6155 VSS.n1739 VSS.n1391 0.00675
R6156 VSS.n1832 VSS.n232 0.00675
R6157 VSS.n1867 VSS.n1866 0.00675
R6158 VSS.n1887 VSS.n1886 0.00675
R6159 VSS.n1893 VSS.n199 0.00675
R6160 VSS.n459 VSS.n456 0.00675
R6161 VSS.n770 VSS.n769 0.00675
R6162 VSS.n486 VSS.n483 0.00675
R6163 VSS.n316 VSS.n311 0.00675
R6164 VSS.n303 VSS.n257 0.00675
R6165 VSS.n1793 VSS.n267 0.00675
R6166 VSS.n349 VSS.n348 0.00675
R6167 VSS.n259 VSS.n256 0.00675
R6168 VSS.n1792 VSS.n1791 0.00675
R6169 VSS.n351 VSS.n270 0.00675
R6170 VSS.n536 VSS.n517 0.00675
R6171 VSS.n716 VSS.n715 0.00675
R6172 VSS.n709 VSS.n548 0.00675
R6173 VSS.n581 VSS.n580 0.00675
R6174 VSS.n612 VSS.n611 0.00675
R6175 VSS.n676 VSS.n675 0.00675
R6176 VSS.n524 VSS.n523 0.00675
R6177 VSS.n717 VSS.n544 0.00675
R6178 VSS.n708 VSS.n550 0.00675
R6179 VSS.n613 VSS.n596 0.00675
R6180 VSS.n674 VSS.n628 0.00675
R6181 VSS.n670 VSS.n634 0.00675
R6182 VSS.n458 VSS.n457 0.00675
R6183 VSS.n771 VSS.n390 0.00675
R6184 VSS.n759 VSS.n402 0.00675
R6185 VSS.n485 VSS.n484 0.00675
R6186 VSS.n755 VSS.n406 0.00675
R6187 VSS.n1051 VSS.n1048 0.00675
R6188 VSS.n1343 VSS.n1342 0.00675
R6189 VSS.n1078 VSS.n1075 0.00675
R6190 VSS.n877 VSS.n856 0.00675
R6191 VSS.n848 VSS.n847 0.00675
R6192 VSS.n939 VSS.n818 0.00675
R6193 VSS.n826 VSS.n825 0.00675
R6194 VSS.n913 VSS.n912 0.00675
R6195 VSS.n940 VSS.n816 0.00675
R6196 VSS.n823 VSS.n817 0.00675
R6197 VSS.n1128 VSS.n1109 0.00675
R6198 VSS.n1289 VSS.n1288 0.00675
R6199 VSS.n1282 VSS.n1140 0.00675
R6200 VSS.n1173 VSS.n1172 0.00675
R6201 VSS.n1204 VSS.n1203 0.00675
R6202 VSS.n1249 VSS.n1248 0.00675
R6203 VSS.n1116 VSS.n1115 0.00675
R6204 VSS.n1290 VSS.n1136 0.00675
R6205 VSS.n1281 VSS.n1142 0.00675
R6206 VSS.n1205 VSS.n1188 0.00675
R6207 VSS.n1247 VSS.n1239 0.00675
R6208 VSS.n1242 VSS.n2 0.00675
R6209 VSS.n1050 VSS.n1049 0.00675
R6210 VSS.n1344 VSS.n982 0.00675
R6211 VSS.n1332 VSS.n994 0.00675
R6212 VSS.n1077 VSS.n1076 0.00675
R6213 VSS.n1328 VSS.n998 0.00675
R6214 VSS.n152 VSS.n143 0.00675
R6215 VSS.n146 VSS.n144 0.00675
R6216 VSS.n2003 VSS.n124 0.00675
R6217 VSS.n150 VSS.n145 0.00675
R6218 VSS.n1969 VSS.n147 0.00675
R6219 VSS.n131 VSS.n128 0.00675
R6220 VSS.n2002 VSS.n2001 0.00675
R6221 VSS.n2000 VSS.n1996 0.00675
R6222 VSS.n2060 VSS.n90 0.00675
R6223 VSS.n2083 VSS.n77 0.00675
R6224 VSS.n2107 VSS.n2106 0.00675
R6225 VSS.n2105 VSS.n64 0.00675
R6226 VSS.n2129 VSS.n50 0.00675
R6227 VSS.n2165 VSS.n2163 0.00675
R6228 VSS.n95 VSS.n92 0.00675
R6229 VSS.n2084 VSS.n78 0.00675
R6230 VSS.n2108 VSS.n62 0.00675
R6231 VSS.n2128 VSS.n2127 0.00675
R6232 VSS.n2166 VSS.n25 0.00675
R6233 VSS.n2167 VSS.n23 0.00675
R6234 VSS.n1861 VSS.n224 0.00675
R6235 VSS.n1888 VSS.n203 0.00675
R6236 VSS.n1897 VSS.n200 0.00675
R6237 VSS.n1520 VSS.n1502 0.00675
R6238 VSS.n1697 VSS.n1532 0.00675
R6239 VSS.n1563 VSS.n1557 0.00675
R6240 VSS.n1565 VSS.n1564 0.00675
R6241 VSS.n1675 VSS.n1578 0.00675
R6242 VSS.n1637 VSS.n1635 0.00675
R6243 VSS.n1508 VSS.n1504 0.00675
R6244 VSS.n1696 VSS.n1695 0.00675
R6245 VSS.n1562 VSS.n1561 0.00675
R6246 VSS.n1676 VSS.n1576 0.00675
R6247 VSS.n1638 VSS.n1631 0.00675
R6248 VSS.n1639 VSS.n1625 0.00675
R6249 VSS.n527 VSS.n511 0.00636816
R6250 VSS.n1119 VSS.n1103 0.00636816
R6251 VSS.n2036 VSS.n2035 0.00636816
R6252 VSS.n1511 VSS.n1496 0.00636816
R6253 VSS.n667 VSS.n635 0.00636785
R6254 VSS.n2194 VSS.n3 0.00636785
R6255 VSS.n22 VSS.n16 0.00636785
R6256 VSS.n1630 VSS.n1624 0.00636785
R6257 VSS.n725 VSS.n724 0.00620714
R6258 VSS.n724 VSS.n723 0.00620714
R6259 VSS.n688 VSS.n618 0.00620714
R6260 VSS.n631 VSS.n618 0.00620714
R6261 VSS.n1298 VSS.n1297 0.00620714
R6262 VSS.n1297 VSS.n1296 0.00620714
R6263 VSS.n1261 VSS.n1210 0.00620714
R6264 VSS.n1244 VSS.n1210 0.00620714
R6265 VSS.n2064 VSS.n80 0.00620714
R6266 VSS.n2090 VSS.n80 0.00620714
R6267 VSS.n2151 VSS.n2150 0.00620714
R6268 VSS.n2150 VSS.n2149 0.00620714
R6269 VSS.n1535 VSS.n1524 0.00620714
R6270 VSS.n1540 VSS.n1535 0.00620714
R6271 VSS.n1661 VSS.n1660 0.00620714
R6272 VSS.n1660 VSS.n1659 0.00620714
R6273 VSS.n532 VSS.n521 0.00587143
R6274 VSS.n554 VSS.n553 0.00587143
R6275 VSS.n617 VSS.n616 0.00587143
R6276 VSS.n672 VSS.n671 0.00587143
R6277 VSS.n1124 VSS.n1113 0.00587143
R6278 VSS.n1146 VSS.n1145 0.00587143
R6279 VSS.n1209 VSS.n1208 0.00587143
R6280 VSS.n1245 VSS.n1 0.00587143
R6281 VSS.n2056 VSS.n93 0.00587143
R6282 VSS.n2091 VSS.n60 0.00587143
R6283 VSS.n2125 VSS.n33 0.00587143
R6284 VSS.n2170 VSS.n2169 0.00587143
R6285 VSS.n1516 VSS.n1506 0.00587143
R6286 VSS.n1559 VSS.n1558 0.00587143
R6287 VSS.n1590 VSS.n1575 0.00587143
R6288 VSS.n1642 VSS.n1641 0.00587143
R6289 VSS.n1433 VSS.n1428 0.00585714
R6290 VSS.n1420 VSS.n1376 0.00585714
R6291 VSS.n1744 VSS.n1385 0.00585714
R6292 VSS.n1472 VSS.n1465 0.00585714
R6293 VSS.n1482 VSS.n1407 0.00585714
R6294 VSS.n1759 VSS.n1369 0.00585714
R6295 VSS.n1378 VSS.n1375 0.00585714
R6296 VSS.n1743 VSS.n1742 0.00585714
R6297 VSS.n1856 VSS.n220 0.00585714
R6298 VSS.n223 VSS.n221 0.00585714
R6299 VSS.n448 VSS.n443 0.00585714
R6300 VSS.n435 VSS.n391 0.00585714
R6301 VSS.n760 VSS.n400 0.00585714
R6302 VSS.n487 VSS.n480 0.00585714
R6303 VSS.n497 VSS.n422 0.00585714
R6304 VSS.n325 VSS.n324 0.00585714
R6305 VSS.n1803 VSS.n1802 0.00585714
R6306 VSS.n323 VSS.n253 0.00585714
R6307 VSS.n1804 VSS.n256 0.00585714
R6308 VSS.n1792 VSS.n269 0.00585714
R6309 VSS.n1787 VSS.n274 0.00585714
R6310 VSS.n719 VSS.n543 0.00585714
R6311 VSS.n610 VSS.n609 0.00585714
R6312 VSS.n646 VSS.n592 0.00585714
R6313 VSS.n650 VSS.n649 0.00585714
R6314 VSS.n647 VSS.n594 0.00585714
R6315 VSS.n775 VSS.n384 0.00585714
R6316 VSS.n393 VSS.n390 0.00585714
R6317 VSS.n759 VSS.n758 0.00585714
R6318 VSS.n1040 VSS.n1035 0.00585714
R6319 VSS.n1027 VSS.n983 0.00585714
R6320 VSS.n1333 VSS.n992 0.00585714
R6321 VSS.n1079 VSS.n1072 0.00585714
R6322 VSS.n1089 VSS.n1014 0.00585714
R6323 VSS.n906 VSS.n905 0.00585714
R6324 VSS.n914 VSS.n840 0.00585714
R6325 VSS.n907 VSS.n844 0.00585714
R6326 VSS.n913 VSS.n841 0.00585714
R6327 VSS.n919 VSS.n816 0.00585714
R6328 VSS.n944 VSS.n812 0.00585714
R6329 VSS.n1292 VSS.n1135 0.00585714
R6330 VSS.n1202 VSS.n1201 0.00585714
R6331 VSS.n1223 VSS.n1184 0.00585714
R6332 VSS.n1227 VSS.n1226 0.00585714
R6333 VSS.n1224 VSS.n1186 0.00585714
R6334 VSS.n1348 VSS.n976 0.00585714
R6335 VSS.n985 VSS.n982 0.00585714
R6336 VSS.n1332 VSS.n1331 0.00585714
R6337 VSS.n1937 VSS.n157 0.00585714
R6338 VSS.n1972 VSS.n1971 0.00585714
R6339 VSS.n1992 VSS.n1991 0.00585714
R6340 VSS.n2004 VSS.n123 0.00585714
R6341 VSS.n114 VSS.n107 0.00585714
R6342 VSS.n161 VSS.n149 0.00585714
R6343 VSS.n1966 VSS.n147 0.00585714
R6344 VSS.n1993 VSS.n128 0.00585714
R6345 VSS.n2086 VSS.n2082 0.00585714
R6346 VSS.n2130 VSS.n49 0.00585714
R6347 VSS.n2145 VSS.n38 0.00585714
R6348 VSS.n43 VSS.n42 0.00585714
R6349 VSS.n40 VSS.n35 0.00585714
R6350 VSS.n1857 VSS.n222 0.00585714
R6351 VSS.n1864 VSS.n224 0.00585714
R6352 VSS.n206 VSS.n203 0.00585714
R6353 VSS.n201 VSS.n186 0.00585714
R6354 VSS.n1698 VSS.n1531 0.00585714
R6355 VSS.n1607 VSS.n1606 0.00585714
R6356 VSS.n1669 VSS.n1582 0.00585714
R6357 VSS.n1665 VSS.n1585 0.00585714
R6358 VSS.n1668 VSS.n1667 0.00585714
R6359 VSS.n1931 VSS.n176 0.00565497
R6360 VSS.n1779 VSS.n282 0.00565497
R6361 VSS.n969 VSS.n796 0.00565497
R6362 VSS.n1730 VSS.n1400 0.00511752
R6363 VSS.n746 VSS.n415 0.00511752
R6364 VSS.n1319 VSS.n1007 0.00511752
R6365 VSS.n2052 VSS.n101 0.00511752
R6366 VSS.n1766 VSS.n1366 0.00496429
R6367 VSS.n1762 VSS.n1369 0.00496429
R6368 VSS.n1738 VSS.n1392 0.00496429
R6369 VSS.n1735 VSS.n1392 0.00496429
R6370 VSS.n1732 VSS.n1398 0.00496429
R6371 VSS.n1899 VSS.n198 0.00496429
R6372 VSS.n189 VSS.n182 0.00496429
R6373 VSS.n353 VSS.n346 0.00496429
R6374 VSS.n364 VSS.n289 0.00496429
R6375 VSS.n1815 VSS.n247 0.00496429
R6376 VSS.n1811 VSS.n250 0.00496429
R6377 VSS.n1808 VSS.n250 0.00496429
R6378 VSS.n1784 VSS.n274 0.00496429
R6379 VSS.n1781 VSS.n280 0.00496429
R6380 VSS.n681 VSS.n625 0.00496429
R6381 VSS.n705 VSS.n704 0.00496429
R6382 VSS.n680 VSS.n627 0.00496429
R6383 VSS.n782 VSS.n381 0.00496429
R6384 VSS.n778 VSS.n384 0.00496429
R6385 VSS.n754 VSS.n407 0.00496429
R6386 VSS.n751 VSS.n407 0.00496429
R6387 VSS.n748 VSS.n413 0.00496429
R6388 VSS.n938 VSS.n937 0.00496429
R6389 VSS.n806 VSS.n803 0.00496429
R6390 VSS.n885 VSS.n863 0.00496429
R6391 VSS.n888 VSS.n861 0.00496429
R6392 VSS.n861 VSS.n843 0.00496429
R6393 VSS.n947 VSS.n812 0.00496429
R6394 VSS.n950 VSS.n794 0.00496429
R6395 VSS.n1254 VSS.n1236 0.00496429
R6396 VSS.n1278 VSS.n1277 0.00496429
R6397 VSS.n1253 VSS.n1238 0.00496429
R6398 VSS.n1355 VSS.n973 0.00496429
R6399 VSS.n1351 VSS.n976 0.00496429
R6400 VSS.n1327 VSS.n999 0.00496429
R6401 VSS.n1324 VSS.n999 0.00496429
R6402 VSS.n1321 VSS.n1005 0.00496429
R6403 VSS.n1945 VSS.n163 0.00496429
R6404 VSS.n1948 VSS.n161 0.00496429
R6405 VSS.n126 VSS.n111 0.00496429
R6406 VSS.n2016 VSS.n111 0.00496429
R6407 VSS.n2019 VSS.n99 0.00496429
R6408 VSS.n2158 VSS.n28 0.00496429
R6409 VSS.n2112 VSS.n2111 0.00496429
R6410 VSS.n2159 VSS.n27 0.00496429
R6411 VSS.n1840 VSS.n238 0.00496429
R6412 VSS.n1843 VSS.n236 0.00496429
R6413 VSS.n236 VSS.n226 0.00496429
R6414 VSS.n1912 VSS.n186 0.00496429
R6415 VSS.n1915 VSS.n174 0.00496429
R6416 VSS.n1657 VSS.n1656 0.00496429
R6417 VSS.n1572 VSS.n1571 0.00496429
R6418 VSS.n1658 VSS.n1593 0.00496429
R6419 VSS.n1805 VSS.n254 0.00486429
R6420 VSS.n1798 VSS.n262 0.00486429
R6421 VSS.n1797 VSS.n263 0.00486429
R6422 VSS.n1790 VSS.n271 0.00486429
R6423 VSS.n772 VSS.n388 0.00486429
R6424 VSS.n765 VSS.n396 0.00486429
R6425 VSS.n764 VSS.n397 0.00486429
R6426 VSS.n757 VSS.n404 0.00486429
R6427 VSS.n911 VSS.n910 0.00486429
R6428 VSS.n918 VSS.n838 0.00486429
R6429 VSS.n922 VSS.n921 0.00486429
R6430 VSS.n941 VSS.n815 0.00486429
R6431 VSS.n1345 VSS.n980 0.00486429
R6432 VSS.n1338 VSS.n988 0.00486429
R6433 VSS.n1337 VSS.n989 0.00486429
R6434 VSS.n1330 VSS.n996 0.00486429
R6435 VSS.n1863 VSS.n1862 0.00486429
R6436 VSS.n1880 VSS.n207 0.00486429
R6437 VSS.n1882 VSS.n1881 0.00486429
R6438 VSS.n1889 VSS.n202 0.00486429
R6439 VSS.n1968 VSS.n1967 0.00486429
R6440 VSS.n1985 VSS.n132 0.00486429
R6441 VSS.n1987 VSS.n1986 0.00486429
R6442 VSS.n1994 VSS.n127 0.00486429
R6443 VSS.n1756 VSS.n1373 0.00486429
R6444 VSS.n1749 VSS.n1381 0.00486429
R6445 VSS.n1748 VSS.n1382 0.00486429
R6446 VSS.n1741 VSS.n1389 0.00486429
R6447 VSS.n632 VSS 0.00452857
R6448 VSS.n2198 VSS 0.00452857
R6449 VSS.n2171 VSS 0.00452857
R6450 VSS VSS.n2200 0.00452857
R6451 VSS.n1855 VSS.n227 0.00407143
R6452 VSS.n326 VSS.n252 0.00407143
R6453 VSS.n528 VSS.n526 0.00407143
R6454 VSS.n728 VSS.n519 0.00407143
R6455 VSS.n721 VSS.n720 0.00407143
R6456 VSS.n668 VSS.n637 0.00407143
R6457 VSS.n727 VSS.n726 0.00407143
R6458 VSS.n722 VSS.n541 0.00407143
R6459 VSS.n603 VSS.n602 0.00407143
R6460 VSS.n858 VSS.n845 0.00407143
R6461 VSS.n1120 VSS.n1118 0.00407143
R6462 VSS.n1301 VSS.n1111 0.00407143
R6463 VSS.n1294 VSS.n1293 0.00407143
R6464 VSS.n2195 VSS.n4 0.00407143
R6465 VSS.n1300 VSS.n1299 0.00407143
R6466 VSS.n1295 VSS.n1133 0.00407143
R6467 VSS.n1195 VSS.n1194 0.00407143
R6468 VSS.n2034 VSS.n96 0.00407143
R6469 VSS.n2068 VSS.n91 0.00407143
R6470 VSS.n2088 VSS.n2087 0.00407143
R6471 VSS.n2175 VSS.n2174 0.00407143
R6472 VSS.n2070 VSS.n2069 0.00407143
R6473 VSS.n2089 VSS.n82 0.00407143
R6474 VSS.n2122 VSS.n55 0.00407143
R6475 VSS.n1512 VSS.n1510 0.00407143
R6476 VSS.n1709 VSS.n1503 0.00407143
R6477 VSS.n1538 VSS.n1537 0.00407143
R6478 VSS.n1646 VSS.n1645 0.00407143
R6479 VSS.n1711 VSS.n1710 0.00407143
R6480 VSS.n1539 VSS.n1536 0.00407143
R6481 VSS.n1680 VSS.n1679 0.00407143
R6482 VSS.n532 VSS.n531 0.00352143
R6483 VSS.n539 VSS.n521 0.00352143
R6484 VSS.n553 VSS.n540 0.00352143
R6485 VSS.n707 VSS.n554 0.00352143
R6486 VSS.n616 VSS.n595 0.00352143
R6487 VSS.n689 VSS.n617 0.00352143
R6488 VSS.n673 VSS.n672 0.00352143
R6489 VSS.n671 VSS.n633 0.00352143
R6490 VSS.n1124 VSS.n1123 0.00352143
R6491 VSS.n1131 VSS.n1113 0.00352143
R6492 VSS.n1145 VSS.n1132 0.00352143
R6493 VSS.n1280 VSS.n1146 0.00352143
R6494 VSS.n1208 VSS.n1187 0.00352143
R6495 VSS.n1262 VSS.n1209 0.00352143
R6496 VSS.n1246 VSS.n1245 0.00352143
R6497 VSS.n2197 VSS.n1 0.00352143
R6498 VSS.n2056 VSS.n2055 0.00352143
R6499 VSS.n2063 VSS.n93 0.00352143
R6500 VSS.n2092 VSS.n2091 0.00352143
R6501 VSS.n2109 VSS.n60 0.00352143
R6502 VSS.n2126 VSS.n2125 0.00352143
R6503 VSS.n2148 VSS.n33 0.00352143
R6504 VSS.n2169 VSS.n24 0.00352143
R6505 VSS.n2172 VSS.n2170 0.00352143
R6506 VSS.n1516 VSS.n1515 0.00352143
R6507 VSS.n1523 VSS.n1506 0.00352143
R6508 VSS.n1558 VSS.n1541 0.00352143
R6509 VSS.n1559 VSS.n1554 0.00352143
R6510 VSS.n1677 VSS.n1575 0.00352143
R6511 VSS.n1591 VSS.n1590 0.00352143
R6512 VSS.n1641 VSS.n1592 0.00352143
R6513 VSS.n1643 VSS.n1642 0.00352143
R6514 VSS.n262 VSS.n254 0.00318571
R6515 VSS.n271 VSS.n263 0.00318571
R6516 VSS.n396 VSS.n388 0.00318571
R6517 VSS.n404 VSS.n397 0.00318571
R6518 VSS.n911 VSS.n838 0.00318571
R6519 VSS.n921 VSS.n815 0.00318571
R6520 VSS.n988 VSS.n980 0.00318571
R6521 VSS.n996 VSS.n989 0.00318571
R6522 VSS.n1862 VSS.n207 0.00318571
R6523 VSS.n1882 VSS.n202 0.00318571
R6524 VSS.n1967 VSS.n132 0.00318571
R6525 VSS.n1987 VSS.n127 0.00318571
R6526 VSS.n1381 VSS.n1373 0.00318571
R6527 VSS.n1389 VSS.n1382 0.00318571
R6528 VSS.n1431 VSS.n1364 0.00317857
R6529 VSS.n1761 VSS.n1370 0.00317857
R6530 VSS.n1746 VSS.n1745 0.00317857
R6531 VSS.n1467 VSS.n1393 0.00317857
R6532 VSS.n1736 VSS.n1394 0.00317857
R6533 VSS.n1731 VSS.n1399 0.00317857
R6534 VSS.n1430 VSS.n1366 0.00317857
R6535 VSS.n1762 VSS.n1368 0.00317857
R6536 VSS.n1747 VSS.n1383 0.00317857
R6537 VSS.n1735 VSS.n1395 0.00317857
R6538 VSS.n1732 VSS.n1397 0.00317857
R6539 VSS.n1839 VSS.n1838 0.00317857
R6540 VSS.n1845 VSS.n235 0.00317857
R6541 VSS.n1878 VSS.n210 0.00317857
R6542 VSS.n1894 VSS.n1893 0.00317857
R6543 VSS.n1911 VSS.n1910 0.00317857
R6544 VSS.n1916 VSS.n175 0.00317857
R6545 VSS.n446 VSS.n378 0.00317857
R6546 VSS.n777 VSS.n385 0.00317857
R6547 VSS.n762 VSS.n761 0.00317857
R6548 VSS.n482 VSS.n408 0.00317857
R6549 VSS.n752 VSS.n409 0.00317857
R6550 VSS.n747 VSS.n414 0.00317857
R6551 VSS.n314 VSS.n245 0.00317857
R6552 VSS.n1810 VSS.n251 0.00317857
R6553 VSS.n1801 VSS.n258 0.00317857
R6554 VSS.n348 VSS.n275 0.00317857
R6555 VSS.n1785 VSS.n276 0.00317857
R6556 VSS.n1780 VSS.n281 0.00317857
R6557 VSS.n313 VSS.n247 0.00317857
R6558 VSS.n1811 VSS.n249 0.00317857
R6559 VSS.n1800 VSS.n1799 0.00317857
R6560 VSS.n1784 VSS.n277 0.00317857
R6561 VSS.n1781 VSS.n279 0.00317857
R6562 VSS.n528 VSS.n527 0.00317857
R6563 VSS.n579 VSS.n558 0.00317857
R6564 VSS.n606 VSS.n605 0.00317857
R6565 VSS.n686 VSS.n621 0.00317857
R6566 VSS.n675 VSS.n629 0.00317857
R6567 VSS.n668 VSS.n667 0.00317857
R6568 VSS.n687 VSS.n619 0.00317857
R6569 VSS.n445 VSS.n381 0.00317857
R6570 VSS.n778 VSS.n383 0.00317857
R6571 VSS.n763 VSS.n398 0.00317857
R6572 VSS.n751 VSS.n410 0.00317857
R6573 VSS.n748 VSS.n412 0.00317857
R6574 VSS.n1038 VSS.n792 0.00317857
R6575 VSS.n1350 VSS.n977 0.00317857
R6576 VSS.n1335 VSS.n1334 0.00317857
R6577 VSS.n1074 VSS.n1000 0.00317857
R6578 VSS.n1325 VSS.n1001 0.00317857
R6579 VSS.n1320 VSS.n1006 0.00317857
R6580 VSS.n884 VSS.n883 0.00317857
R6581 VSS.n890 VSS.n860 0.00317857
R6582 VSS.n915 VSS.n833 0.00317857
R6583 VSS.n826 VSS.n813 0.00317857
R6584 VSS.n946 VSS.n802 0.00317857
R6585 VSS.n952 VSS.n795 0.00317857
R6586 VSS.n885 VSS.n864 0.00317857
R6587 VSS.n889 VSS.n888 0.00317857
R6588 VSS.n917 VSS.n916 0.00317857
R6589 VSS.n947 VSS.n804 0.00317857
R6590 VSS.n951 VSS.n950 0.00317857
R6591 VSS.n1120 VSS.n1119 0.00317857
R6592 VSS.n1171 VSS.n1150 0.00317857
R6593 VSS.n1198 VSS.n1197 0.00317857
R6594 VSS.n1259 VSS.n1213 0.00317857
R6595 VSS.n1248 VSS.n1240 0.00317857
R6596 VSS.n2195 VSS.n2194 0.00317857
R6597 VSS.n1260 VSS.n1211 0.00317857
R6598 VSS.n1037 VSS.n973 0.00317857
R6599 VSS.n1351 VSS.n975 0.00317857
R6600 VSS.n1336 VSS.n990 0.00317857
R6601 VSS.n1324 VSS.n1002 0.00317857
R6602 VSS.n1321 VSS.n1004 0.00317857
R6603 VSS.n1944 VSS.n1943 0.00317857
R6604 VSS.n1950 VSS.n160 0.00317857
R6605 VSS.n1990 VSS.n129 0.00317857
R6606 VSS.n1999 VSS.n1998 0.00317857
R6607 VSS.n2015 VSS.n2014 0.00317857
R6608 VSS.n2020 VSS.n100 0.00317857
R6609 VSS.n1945 VSS.n164 0.00317857
R6610 VSS.n1949 VSS.n1948 0.00317857
R6611 VSS.n1989 VSS.n130 0.00317857
R6612 VSS.n2016 VSS.n112 0.00317857
R6613 VSS.n2021 VSS.n2019 0.00317857
R6614 VSS.n2035 VSS.n2034 0.00317857
R6615 VSS.n69 VSS.n68 0.00317857
R6616 VSS.n2119 VSS.n56 0.00317857
R6617 VSS.n2153 VSS.n30 0.00317857
R6618 VSS.n2165 VSS.n2164 0.00317857
R6619 VSS.n2174 VSS.n22 0.00317857
R6620 VSS.n2152 VSS.n31 0.00317857
R6621 VSS.n1840 VSS.n239 0.00317857
R6622 VSS.n1844 VSS.n1843 0.00317857
R6623 VSS.n1879 VSS.n208 0.00317857
R6624 VSS.n1912 VSS.n187 0.00317857
R6625 VSS.n1917 VSS.n1915 0.00317857
R6626 VSS.n1512 VSS.n1511 0.00317857
R6627 VSS.n1569 VSS.n1556 0.00317857
R6628 VSS.n1603 VSS.n1551 0.00317857
R6629 VSS.n1664 VSS.n1663 0.00317857
R6630 VSS.n1637 VSS.n1636 0.00317857
R6631 VSS.n1645 VSS.n1624 0.00317857
R6632 VSS.n1662 VSS.n1584 0.00317857
R6633 VSS.n1440 VSS.n1371 0.00228571
R6634 VSS.n1445 VSS.n1440 0.00228571
R6635 VSS.n1441 VSS.n1420 0.00228571
R6636 VSS.n1752 VSS.n1377 0.00228571
R6637 VSS.n1472 VSS.n1471 0.00228571
R6638 VSS.n1751 VSS.n1750 0.00228571
R6639 VSS.n1867 VSS.n220 0.00228571
R6640 VSS.n1885 VSS.n204 0.00228571
R6641 VSS.n1899 VSS.n1898 0.00228571
R6642 VSS.n455 VSS.n386 0.00228571
R6643 VSS.n460 VSS.n455 0.00228571
R6644 VSS.n456 VSS.n435 0.00228571
R6645 VSS.n768 VSS.n392 0.00228571
R6646 VSS.n487 VSS.n486 0.00228571
R6647 VSS.n324 VSS.n303 0.00228571
R6648 VSS.n1795 VSS.n1794 0.00228571
R6649 VSS.n353 VSS.n352 0.00228571
R6650 VSS.n1796 VSS.n265 0.00228571
R6651 VSS.n566 VSS.n519 0.00228571
R6652 VSS.n716 VSS.n543 0.00228571
R6653 VSS.n710 VSS.n709 0.00228571
R6654 VSS.n650 VSS.n646 0.00228571
R6655 VSS.n625 VSS.n622 0.00228571
R6656 VSS.n767 VSS.n766 0.00228571
R6657 VSS.n1047 VSS.n978 0.00228571
R6658 VSS.n1052 VSS.n1047 0.00228571
R6659 VSS.n1048 VSS.n1027 0.00228571
R6660 VSS.n1341 VSS.n984 0.00228571
R6661 VSS.n1079 VSS.n1078 0.00228571
R6662 VSS.n905 VSS.n848 0.00228571
R6663 VSS.n836 VSS.n835 0.00228571
R6664 VSS.n937 VSS.n819 0.00228571
R6665 VSS.n923 VSS.n837 0.00228571
R6666 VSS.n1158 VSS.n1111 0.00228571
R6667 VSS.n1289 VSS.n1135 0.00228571
R6668 VSS.n1283 VSS.n1282 0.00228571
R6669 VSS.n1227 VSS.n1223 0.00228571
R6670 VSS.n1236 VSS.n1214 0.00228571
R6671 VSS.n1340 VSS.n1339 0.00228571
R6672 VSS.n1961 VSS.n151 0.00228571
R6673 VSS.n1961 VSS.n1960 0.00228571
R6674 VSS.n1972 VSS.n143 0.00228571
R6675 VSS.n1983 VSS.n135 0.00228571
R6676 VSS.n2004 VSS.n2003 0.00228571
R6677 VSS.n1984 VSS.n133 0.00228571
R6678 VSS.n2068 VSS.n2067 0.00228571
R6679 VSS.n2083 VSS.n2082 0.00228571
R6680 VSS.n2107 VSS.n63 0.00228571
R6681 VSS.n43 VSS.n38 0.00228571
R6682 VSS.n2155 VSS.n28 0.00228571
R6683 VSS.n1884 VSS.n205 0.00228571
R6684 VSS.n1709 VSS.n1708 0.00228571
R6685 VSS.n1698 VSS.n1697 0.00228571
R6686 VSS.n1557 VSS.n1543 0.00228571
R6687 VSS.n1585 VSS.n1582 0.00228571
R6688 VSS.n1657 VSS.n1594 0.00228571
R6689 VSS.n1814 VSS.n1813 0.00217857
R6690 VSS.n1812 VSS.n248 0.00217857
R6691 VSS.n1783 VSS.n272 0.00217857
R6692 VSS.n1782 VSS.n278 0.00217857
R6693 VSS.n781 VSS.n780 0.00217857
R6694 VSS.n779 VSS.n382 0.00217857
R6695 VSS.n750 VSS.n405 0.00217857
R6696 VSS.n749 VSS.n411 0.00217857
R6697 VSS.n886 VSS.n862 0.00217857
R6698 VSS.n887 VSS.n842 0.00217857
R6699 VSS.n948 VSS.n811 0.00217857
R6700 VSS.n949 VSS.n793 0.00217857
R6701 VSS.n1354 VSS.n1353 0.00217857
R6702 VSS.n1352 VSS.n974 0.00217857
R6703 VSS.n1323 VSS.n997 0.00217857
R6704 VSS.n1322 VSS.n1003 0.00217857
R6705 VSS.n1841 VSS.n237 0.00217857
R6706 VSS.n1842 VSS.n225 0.00217857
R6707 VSS.n1913 VSS.n185 0.00217857
R6708 VSS.n1914 VSS.n173 0.00217857
R6709 VSS.n1946 VSS.n162 0.00217857
R6710 VSS.n1947 VSS.n148 0.00217857
R6711 VSS.n2017 VSS.n110 0.00217857
R6712 VSS.n2018 VSS.n98 0.00217857
R6713 VSS.n1765 VSS.n1764 0.00217857
R6714 VSS.n1763 VSS.n1367 0.00217857
R6715 VSS.n1734 VSS.n1390 0.00217857
R6716 VSS.n1733 VSS.n1396 0.00217857
R6717 VSS.n1481 VSS.n1410 0.00139286
R6718 VSS.n1487 VSS.n1407 0.00139286
R6719 VSS.n1877 VSS.n212 0.00139286
R6720 VSS.n1909 VSS.n191 0.00139286
R6721 VSS.n1921 VSS.n182 0.00139286
R6722 VSS.n496 VSS.n425 0.00139286
R6723 VSS.n502 VSS.n422 0.00139286
R6724 VSS.n297 VSS.n266 0.00139286
R6725 VSS.n363 VSS.n292 0.00139286
R6726 VSS.n369 VSS.n289 0.00139286
R6727 VSS.n264 VSS.n261 0.00139286
R6728 VSS.n609 VSS.n597 0.00139286
R6729 VSS.n612 VSS.n591 0.00139286
R6730 VSS.n600 VSS.n598 0.00139286
R6731 VSS.n614 VSS.n613 0.00139286
R6732 VSS.n1088 VSS.n1017 0.00139286
R6733 VSS.n1094 VSS.n1014 0.00139286
R6734 VSS.n926 VSS.n925 0.00139286
R6735 VSS.n959 VSS.n958 0.00139286
R6736 VSS.n810 VSS.n806 0.00139286
R6737 VSS.n924 VSS.n834 0.00139286
R6738 VSS.n1201 VSS.n1189 0.00139286
R6739 VSS.n1204 VSS.n1183 0.00139286
R6740 VSS.n1192 VSS.n1190 0.00139286
R6741 VSS.n1206 VSS.n1205 0.00139286
R6742 VSS.n2013 VSS.n116 0.00139286
R6743 VSS.n2025 VSS.n107 0.00139286
R6744 VSS.n2120 VSS.n49 0.00139286
R6745 VSS.n52 VSS.n50 0.00139286
R6746 VSS.n2121 VSS.n51 0.00139286
R6747 VSS.n2127 VSS.n53 0.00139286
R6748 VSS.n211 VSS.n209 0.00139286
R6749 VSS.n1606 VSS.n1604 0.00139286
R6750 VSS.n1675 VSS.n1674 0.00139286
R6751 VSS.n1605 VSS.n1553 0.00139286
R6752 VSS.n1676 VSS.n1577 0.00139286
R6753 VSS.n2199 VSS.n2198 0.00054824
R6754 VSS.n632 VSS.n0 0.00054824
R6755 D2 D2.n0 125.046
R6756 D2.n0 D2.t0 77.1205
R6757 D2.n0 D2.t1 61.6965
R6758 D2_BUF.n2 D2_BUF.n1 173.293
R6759 D2_BUF.n1 D2_BUF.t3 84.3505
R6760 D2_BUF.n1 D2_BUF.t2 53.5025
R6761 D2_BUF.n0 D2_BUF.t0 46.9077
R6762 D2_BUF.n0 D2_BUF.t1 35.0239
R6763 D2_BUF D2_BUF.n2 3.75226
R6764 D2_BUF.n2 D2_BUF.n0 0.204238
R6765 D3_BUF.n2 D3_BUF.n1 173.293
R6766 D3_BUF.n1 D3_BUF.t2 84.3505
R6767 D3_BUF.n1 D3_BUF.t3 53.5025
R6768 D3_BUF.n0 D3_BUF.t0 46.9077
R6769 D3_BUF.n0 D3_BUF.t1 35.0239
R6770 D3_BUF D3_BUF.n2 3.75099
R6771 D3_BUF.n2 D3_BUF.n0 0.204238
R6772 D0 D0.n0 115.853
R6773 D0.n0 D0.t0 81.9405
R6774 D0.n0 D0.t1 56.8765
R6775 VOUT.n0 VOUT.t1 46.8495
R6776 VOUT.n0 VOUT.t2 46.5654
R6777 VOUT.n5 VOUT.t0 34.887
R6778 VOUT.n10 VOUT.t3 27.6955
R6779 VOUT.n4 VOUT.n3 13.362
R6780 VOUT.n2 VOUT.n1 9.3005
R6781 VOUT.n7 VOUT.n6 9.3005
R6782 VOUT.n9 VOUT.n8 9.3005
R6783 VOUT.n12 VOUT.n11 9.3005
R6784 VOUT.n11 VOUT.n10 9.02061
R6785 VOUT.n5 VOUT.n4 4.55875
R6786 VOUT.n0 VOUT 3.09322
R6787 VOUT VOUT.n12 0.815717
R6788 VOUT.n2 VOUT.n0 0.613
R6789 VOUT.n12 VOUT.n9 0.0439783
R6790 VOUT.n7 VOUT.n5 0.0439783
R6791 VOUT.n5 VOUT.n2 0.014087
R6792 VOUT.n9 VOUT.n7 0.00321739
R6793 D3 D3.n0 125.046
R6794 D3.n0 D3.t1 77.1205
R6795 D3.n0 D3.t0 61.6965
R6796 D1.n1 D1.n0 127.099
R6797 D1.n0 D1.t1 77.6025
R6798 D1.n0 D1.t0 61.2145
R6799 D1.n1 D1 0.0485769
R6800 D1 D1.n1 0.0365577
R6801 D1_BUF.n2 D1_BUF.n1 169.566
R6802 D1_BUF.n1 D1_BUF.t2 84.8325
R6803 D1_BUF.n1 D1_BUF.t3 53.0205
R6804 D1_BUF.n0 D1_BUF.t0 46.9158
R6805 D1_BUF.n0 D1_BUF.t1 35.0302
R6806 D1_BUF.n3 D1_BUF.n2 3.65455
R6807 D1_BUF D1_BUF.n3 2.60341
R6808 D1_BUF.n2 D1_BUF.n0 0.199588
R6809 D1_BUF.n3 D1_BUF 0.0389615
R6810 VREFL.n1 VREFL.t1 99.7169
R6811 VREFL.n0 VREFL.t2 44.9543
R6812 VREFL.n0 VREFL.t0 37.5373
R6813 VREFL.n1 VREFL.n0 2.88557
R6814 VREFL VREFL.n1 1.84958
R6815 VREFH VREFH.t0 98.071
C778 switch_n_3v3_0.D7 VSS 0.701f
C779 switch_n_3v3_0.D6 VSS 0.295f
C780 switch_n_3v3_0.D5 VSS 0.29f
C781 switch_n_3v3_0.D4 VSS 0.289f
C782 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS 0.667f 
C783 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS 1.53f 
C784 D1_BUF VSS 1.17f
C785 3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS 1.13f 
C786 D0_BUF VSS 2.53f
C787 a_1556_406# VSS 1.22f 
C788 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS 0.676f 
C789 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS 0.519f 
C790 VREFH VSS 0.29f
C791 3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH VSS 0.544f 
C792 3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS 1.32f 
C793 3_bit_dac_0[0].2_bit_dac_0[1].VOUT VSS 1.08f 
C794 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS 0.627f 
C795 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS 1.07f 
C796 D2_BUF VSS 1.14f
C797 3_bit_dac_0[0].switch_n_3v3_1.DX_ VSS 1.14f 
C798 3_bit_dac_0[0].2_bit_dac_0[0].D1 VSS 1.63f 
C799 3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS 1.06f 
C800 3_bit_dac_0[0].2_bit_dac_0[0].D0 VSS 3.26f 
C801 a_1556_1634# VSS 1.16f 
C802 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS 0.663f 
C803 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS 0.467f 
C804 3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS 1.5f 
C805 3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH VSS 0.543f 
C806 3_bit_dac_0[0].VOUT VSS 0.951f 
C807 VOUT VSS 0.378f
C808 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS 0.633f 
C809 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS 1.07f 
C810 D3_BUF VSS 1.17f
C811 switch_n_3v3_0.DX_ VSS 1.09f 
C812 D3 VSS 0.641f
C813 3_bit_dac_0[0].D1 VSS 1.61f 
C814 3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS 1.06f 
C815 3_bit_dac_0[0].D0 VSS 3.25f 
C816 a_1556_2862# VSS 1.16f 
C817 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS 0.663f 
C818 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS 0.467f 
C819 3_bit_dac_0[1].VREFH VSS 1.42f 
C820 3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH VSS 0.543f 
C821 3_bit_dac_0[1].2_bit_dac_0[0].VOUT VSS 0.984f 
C822 3_bit_dac_0[1].VOUT VSS 0.944f 
C823 3_bit_dac_0[1].2_bit_dac_0[1].VOUT VSS 1.36f 
C824 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS 0.905f 
C825 VREFL VSS 1.15f
C826 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS 1.11f 
C827 switch_n_3v3_0.D2 VSS 1.87f 
C828 3_bit_dac_0[1].switch_n_3v3_1.DX_ VSS 1.1f 
C829 D2 VSS 0.59f
C830 3_bit_dac_0[1].2_bit_dac_0[0].D1 VSS 1.61f 
C831 3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS 1.08f 
C832 D1 VSS 0.48f
C833 3_bit_dac_0[1].2_bit_dac_0[0].D0 VSS 3.35f 
C834 a_1556_4090# VSS 1.18f 
C835 D0 VSS 0.729f
C836 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS 0.68f 
C837 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS 0.521f 
C838 3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS 1.42f 
C839 3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH VSS 0.714f 
C840 VCC VSS 43.8f
.ends

X1 D0 VREFL D0_BUF VREFH D1 D1_BUF D2 D3 D2_BUF D3_BUF VOUT VSS VCC x4_bit_dac


.param mc_mm_switch=0
.param mc_pr_switch=0
.lib "/foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice.tt.red" tt

V1 VSS 0 dc 0
V2 VCC 0 dc 3.3

V3 VREFL 0 dc 0
V4 VREFH 0 dc 3.3

V5  D0 0 PULSE(0 1.8 4n 1p 1p 4n 8n)
V6  D1 0 PULSE(0 1.8 8n 1p 1p 8n 16n)
V7  D2 0 PULSE(0 1.8 16n 1p 1p 16n 32n)
V8  D3 0 PULSE(0 1.8 32n 1p 1p 32n 64n)


.tran 0.1n 128n uic


.control
run

set xbrushwidth=3
set hcopydevtype = svg

plot D0 D1 D2 D3 VOUT

hardcopy 4_bit_dac_RCX.svg D0 D1 D2 D3 VOUT

.endc
.end
