* SPICE3 file created from 3_bit_dac.ext - technology: sky130A

.subckt x3_bit_dac D0 VREFL D0_BUF VREFH D1 D1_BUF D2 D2_BUF VOUT VSS VCC
X0 2_bit_dac_0[1].switch2n_3v3_0.VREFH 2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t21 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X1 a_1438_1634# D0.t0 VSS.t27 VSS.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2 a_1438_406# 2_bit_dac_0[0].D0 VCC.t33 VCC.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X3 D0_BUF.t0 a_1438_406# VCC.t12 VCC.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X4 2_bit_dac_0[0].switch2n_3v3_0.VOUTH 2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 2_bit_dac_0[0].VOUT VCC.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X5 2_bit_dac_0[0].D0 a_1438_1634# VSS.t25 VSS.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6 2_bit_dac_0[1].VREFH D0_BUF.t2 2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X7 2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1438_406# 2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8 2_bit_dac_0[1].switch2n_3v3_0.R_L VREFL.t1 VSS.t15 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X9 2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ D1.t0 VCC.t1 VCC.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X10 2_bit_dac_0[1].VOUT 2_bit_dac_0[0].D1 2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X11 2_bit_dac_0[1].VOUT switch_n_3v3_1.DX_ VOUT.t1 VSS.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X12 2_bit_dac_0[0].switch2n_3v3_0.R_H D0_BUF.t3 2_bit_dac_0[0].switch2n_3v3_0.VOUTH VCC.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X13 2_bit_dac_0[1].switch2n_3v3_0.VOUTH 2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 2_bit_dac_0[1].VOUT VCC.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X14 2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1438_406# 2_bit_dac_0[1].VREFH VSS.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X15 2_bit_dac_0[1].switch2n_3v3_0.VREFH 2_bit_dac_0[0].D0 2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X16 2_bit_dac_0[0].switch2n_3v3_0.VOUTL 2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 2_bit_dac_0[0].VOUT VSS.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X17 VREFL.t2 2_bit_dac_0[0].D0 2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X18 2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 2_bit_dac_0[0].D1 VSS.t5 VSS.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X19 2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1438_1634# 2_bit_dac_0[1].switch2n_3v3_0.VREFH VCC.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X20 2_bit_dac_0[0].D1 2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VCC.t28 VCC.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X21 2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 2_bit_dac_0[1].VOUT VSS.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X22 D2_BUF.t1 switch_n_3v3_1.DX_ VSS.t1 VSS.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X23 D1_BUF.t0 2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VCC.t17 VCC.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X24 switch_n_3v3_1.DX_ D2.t0 VCC.t26 VCC.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X25 2_bit_dac_0[0].switch2n_3v3_0.VREFH 2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t21 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X26 2_bit_dac_0[0].switch2n_3v3_0.R_H 2_bit_dac_0[0].switch2n_3v3_0.R_L VSS.t19 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X27 2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1438_1634# 2_bit_dac_0[1].switch2n_3v3_0.R_L VCC.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X28 a_1438_1634# D0.t1 VCC.t14 VCC.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X29 VOUT.t2 D2_BUF.t2 2_bit_dac_0[1].VOUT VCC.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X30 2_bit_dac_0[0].switch2n_3v3_0.R_L 2_bit_dac_0[1].VREFH VSS.t15 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X31 a_1438_406# 2_bit_dac_0[0].D0 VSS.t34 VSS.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X32 D0_BUF.t1 a_1438_406# VSS.t9 VSS.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X33 2_bit_dac_0[0].VOUT D1_BUF.t2 2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X34 2_bit_dac_0[0].D0 a_1438_1634# VCC.t21 VCC.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X35 2_bit_dac_0[0].switch2n_3v3_0.R_L D0_BUF.t4 2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X36 2_bit_dac_0[1].switch2n_3v3_0.R_H 2_bit_dac_0[1].switch2n_3v3_0.R_L VSS.t19 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X37 2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ D1.t1 VSS.t14 VSS.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X38 2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1438_406# 2_bit_dac_0[0].switch2n_3v3_0.VREFH VCC.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X39 VOUT.t3 D2_BUF.t3 2_bit_dac_0[0].VOUT VSS.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X40 2_bit_dac_0[0].switch2n_3v3_0.VREFH D0_BUF.t5 2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X41 2_bit_dac_0[0].switch2n_3v3_0.VREFH VREFH.t0 VSS.t12 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X42 2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1438_406# 2_bit_dac_0[0].switch2n_3v3_0.R_L VCC.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X43 2_bit_dac_0[1].switch2n_3v3_0.VREFH 2_bit_dac_0[1].VREFH VSS.t12 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X44 2_bit_dac_0[0].VOUT D1_BUF.t3 2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X45 2_bit_dac_0[1].switch2n_3v3_0.R_H 2_bit_dac_0[0].D0 2_bit_dac_0[1].switch2n_3v3_0.VOUTH VCC.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X46 2_bit_dac_0[1].switch2n_3v3_0.R_L 2_bit_dac_0[0].D0 2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X47 2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1438_1634# 2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X48 2_bit_dac_0[0].D1 2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS.t30 VSS.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X49 2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 2_bit_dac_0[0].D1 VCC.t8 VCC.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X50 D2_BUF.t0 switch_n_3v3_1.DX_ VCC.t4 VCC.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X51 D1_BUF.t1 2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS.t17 VSS.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X52 switch_n_3v3_1.DX_ D2.t1 VSS.t37 VSS.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X53 2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1438_1634# VREFL.t0 VSS.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X54 2_bit_dac_0[1].VOUT 2_bit_dac_0[0].D1 2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X55 2_bit_dac_0[0].VOUT switch_n_3v3_1.DX_ VOUT.t0 VCC.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
C0 2_bit_dac_0[0].switch2n_3v3_0.VOUTH 2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00123f
C1 2_bit_dac_0[0].switch2n_3v3_0.R_H 2_bit_dac_0[1].switch2n_3v3_0.VOUTH 1.68e-19
C2 switch_n_3v3_1.DX_ switch_n_3v3_1.D7 0.0268f
C3 switch_n_3v3_1.D3 2_bit_dac_0[0].D1 2.79e-20
C4 switch_n_3v3_1.DX_ D2_BUF 0.219f
C5 D1_BUF 2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.176f
C6 D1_BUF 2_bit_dac_0[0].switch2n_3v3_0.R_H 0.00237f
C7 VCC 2_bit_dac_0[0].VOUT 0.379f
C8 D0_BUF VCC 0.732f
C9 D1 2_bit_dac_0[0].D0 0.0179f
C10 D2_BUF D1 1.48e-19
C11 D1_BUF 2_bit_dac_0[1].VREFH 3.54e-19
C12 switch_n_3v3_1.DX_ 2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00394f
C13 2_bit_dac_0[1].switch2n_3v3_0.R_H 2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.00832f
C14 D2_BUF switch_n_3v3_1.D3 0.302f
C15 D1 2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.007f
C16 D1 VREFL 1.7e-19
C17 2_bit_dac_0[1].switch2n_3v3_0.VOUTH 2_bit_dac_0[0].VOUT 0.00114f
C18 2_bit_dac_0[0].D1 2_bit_dac_0[1].switch2n_3v3_0.R_H 0.00237f
C19 switch_n_3v3_1.D3 2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0269f
C20 D1_BUF 2_bit_dac_0[0].VOUT 0.0757f
C21 D1 2_bit_dac_0[1].switch2n_3v3_0.R_L 0.00319f
C22 D0_BUF 2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00164f
C23 D2 VCC 0.331f
C24 D0_BUF D1_BUF 0.00262f
C25 2_bit_dac_0[1].VOUT switch_n_3v3_1.D6 0.0234f
C26 2_bit_dac_0[1].switch2n_3v3_0.R_H 2_bit_dac_0[0].D0 0.24f
C27 2_bit_dac_0[0].D1 switch_n_3v3_1.D5 2.05e-20
C28 D1 2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.00491f
C29 switch_n_3v3_1.DX_ switch_n_3v3_1.D4 1.33e-19
C30 2_bit_dac_0[0].D1 2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.00491f
C31 2_bit_dac_0[1].switch2n_3v3_0.R_H VREFL 0.138f
C32 2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2_bit_dac_0[1].switch2n_3v3_0.R_H 0.115f
C33 2_bit_dac_0[1].switch2n_3v3_0.R_H D0 0.117f
C34 D2 2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00872f
C35 switch_n_3v3_1.DX_ 2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 1.79e-20
C36 2_bit_dac_0[0].switch2n_3v3_0.VOUTL 2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.322f
C37 D1 switch_n_3v3_1.D4 1.41e-21
C38 D2_BUF switch_n_3v3_1.D5 0.0293f
C39 2_bit_dac_0[1].switch2n_3v3_0.R_H 2_bit_dac_0[1].switch2n_3v3_0.R_L 0.805f
C40 2_bit_dac_0[0].D1 2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00805f
C41 D1 2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.111f
C42 2_bit_dac_0[0].switch2n_3v3_0.VREFH 2_bit_dac_0[0].D0 0.0824f
C43 switch_n_3v3_1.D3 switch_n_3v3_1.D4 0.625f
C44 2_bit_dac_0[1].switch2n_3v3_0.VOUTL switch_n_3v3_1.D5 0.00306f
C45 D1 2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3.53e-19
C46 switch_n_3v3_1.D3 2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.00213f
C47 2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 2_bit_dac_0[0].switch2n_3v3_0.VREFH 5.89e-20
C48 2_bit_dac_0[0].D1 switch_n_3v3_1.D7 1.57e-20
C49 2_bit_dac_0[0].switch2n_3v3_0.R_L VCC 0.29f
C50 2_bit_dac_0[0].D1 2_bit_dac_0[0].D0 0.00262f
C51 D2_BUF 2_bit_dac_0[0].D1 0.00779f
C52 2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0102f
C53 VREFL 2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0551f
C54 switch_n_3v3_1.DX_ VOUT 0.236f
C55 D0 2_bit_dac_0[0].switch2n_3v3_0.VREFH 1.9e-19
C56 switch_n_3v3_1.D3 2_bit_dac_0[0].switch2n_3v3_0.VOUTH 1.15e-19
C57 2_bit_dac_0[0].switch2n_3v3_0.VOUTL 2_bit_dac_0[0].D0 2.38e-19
C58 2_bit_dac_0[1].switch2n_3v3_0.R_H 2_bit_dac_0[1].switch2n_3v3_0.VREFH 1.39f
C59 2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 2_bit_dac_0[0].D1 0.111f
C60 2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2_bit_dac_0[0].D1 0.635f
C61 2_bit_dac_0[0].D1 VREFL 3.54e-19
C62 2_bit_dac_0[1].switch2n_3v3_0.R_L 2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.00577f
C63 2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.128f
C64 switch_n_3v3_1.DX_ 2_bit_dac_0[0].VOUT 0.088f
C65 2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.0107f
C66 2_bit_dac_0[0].switch2n_3v3_0.VOUTL VREFL 2.66e-20
C67 D2_BUF switch_n_3v3_1.D7 0.0399f
C68 a_1438_406# 2_bit_dac_0[1].switch2n_3v3_0.R_H 4.83e-19
C69 switch_n_3v3_1.D3 VOUT 1.41e-20
C70 2_bit_dac_0[0].D1 2_bit_dac_0[1].switch2n_3v3_0.R_L 2.51e-20
C71 2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 2_bit_dac_0[1].switch2n_3v3_0.R_H 0.00819f
C72 2_bit_dac_0[0].switch2n_3v3_0.R_L D1_BUF 2.51e-20
C73 2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2_bit_dac_0[0].D0 0.38f
C74 VREFL 2_bit_dac_0[0].D0 0.544f
C75 2_bit_dac_0[1].switch2n_3v3_0.VOUTL switch_n_3v3_1.D7 0.00143f
C76 D2_BUF 2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0668f
C77 D0 2_bit_dac_0[0].D0 0.0255f
C78 2_bit_dac_0[1].switch2n_3v3_0.R_H 2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5.59e-19
C79 2_bit_dac_0[1].switch2n_3v3_0.VREFH 2_bit_dac_0[0].switch2n_3v3_0.VREFH 3.82e-19
C80 VREFH 2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0124f
C81 2_bit_dac_0[0].switch2n_3v3_0.R_H 2_bit_dac_0[1].switch2n_3v3_0.R_H 0.0261f
C82 switch_n_3v3_1.D3 2_bit_dac_0[0].VOUT 0.0201f
C83 VCC 2_bit_dac_0[1].VOUT 0.77f
C84 switch_n_3v3_1.D4 switch_n_3v3_1.D5 0.67f
C85 2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 2_bit_dac_0[1].switch2n_3v3_0.VOUTL 7.75e-19
C86 2_bit_dac_0[1].switch2n_3v3_0.VOUTL VREFL 0.404f
C87 2_bit_dac_0[1].switch2n_3v3_0.R_H 2_bit_dac_0[1].VREFH 0.0579f
C88 2_bit_dac_0[1].switch2n_3v3_0.R_L 2_bit_dac_0[0].D0 0.315f
C89 2_bit_dac_0[1].switch2n_3v3_0.VOUTL D0 8.97e-20
C90 VREFL D0 0.77f
C91 2_bit_dac_0[0].D1 2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.00375f
C92 2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ switch_n_3v3_1.D5 2.07e-19
C93 switch_n_3v3_1.DX_ D2 0.0904f
C94 a_1438_406# 2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.175f
C95 2_bit_dac_0[0].switch2n_3v3_0.VOUTH switch_n_3v3_1.D5 5.19e-20
C96 2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2_bit_dac_0[1].switch2n_3v3_0.R_L 0.189f
C97 VREFL 2_bit_dac_0[1].switch2n_3v3_0.R_L 0.482f
C98 2_bit_dac_0[1].switch2n_3v3_0.R_L D0 0.253f
C99 VCC a_1438_1634# 0.713f
C100 2_bit_dac_0[0].D1 switch_n_3v3_1.D4 2.38e-20
C101 VCC switch_n_3v3_1.D6 0.0601f
C102 D1 D2 0.00881f
C103 a_1438_406# 2_bit_dac_0[0].D1 0.003f
C104 2_bit_dac_0[0].switch2n_3v3_0.VOUTH 2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.236f
C105 2_bit_dac_0[1].VOUT 2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.514f
C106 2_bit_dac_0[0].switch2n_3v3_0.R_H 2_bit_dac_0[0].switch2n_3v3_0.VREFH 1.39f
C107 2_bit_dac_0[1].switch2n_3v3_0.VREFH 2_bit_dac_0[0].D0 0.472f
C108 2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 2_bit_dac_0[0].D1 0.219f
C109 VREFH 2_bit_dac_0[0].D0 0.0104f
C110 D1_BUF 2_bit_dac_0[1].VOUT 1.81e-20
C111 a_1438_406# 2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.296f
C112 switch_n_3v3_1.D3 D2 0.348f
C113 2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.0172f
C114 D0_BUF 2_bit_dac_0[1].switch2n_3v3_0.R_H 0.00379f
C115 2_bit_dac_0[1].VREFH 2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.205f
C116 VOUT switch_n_3v3_1.D5 1.98e-20
C117 2_bit_dac_0[0].D1 2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0801f
C118 2_bit_dac_0[0].switch2n_3v3_0.R_H 2_bit_dac_0[0].D1 0.037f
C119 2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.322f
C120 2_bit_dac_0[1].switch2n_3v3_0.VREFH VREFL 0.201f
C121 2_bit_dac_0[1].switch2n_3v3_0.VREFH D0 0.0572f
C122 D2_BUF switch_n_3v3_1.D4 0.0295f
C123 2_bit_dac_0[0].switch2n_3v3_0.VOUTH 2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.579f
C124 a_1438_406# 2_bit_dac_0[0].D0 0.0981f
C125 2_bit_dac_0[0].switch2n_3v3_0.R_H 2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.115f
C126 2_bit_dac_0[0].D1 2_bit_dac_0[1].VREFH 1.7e-19
C127 2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1438_1634# 0.0892f
C128 2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 2_bit_dac_0[0].D0 5.84e-19
C129 2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ switch_n_3v3_1.D7 1.45e-19
C130 D2_BUF 2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.00132f
C131 2_bit_dac_0[1].switch2n_3v3_0.VOUTH switch_n_3v3_1.D6 6.1e-19
C132 switch_n_3v3_1.D5 2_bit_dac_0[0].VOUT 0.0199f
C133 2_bit_dac_0[1].switch2n_3v3_0.VREFH 2_bit_dac_0[1].switch2n_3v3_0.R_L 0.0923f
C134 2_bit_dac_0[1].VREFH 2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.404f
C135 2_bit_dac_0[1].switch2n_3v3_0.VOUTL switch_n_3v3_1.D4 0.00517f
C136 a_1438_406# 2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 1.21e-20
C137 2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.0104f
C138 2_bit_dac_0[0].switch2n_3v3_0.VOUTH switch_n_3v3_1.D7 2.94e-20
C139 a_1438_406# VREFL 1.97e-19
C140 2_bit_dac_0[0].switch2n_3v3_0.VOUTH 2_bit_dac_0[0].D0 3.36e-19
C141 a_1438_406# 2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00538f
C142 D2_BUF 2_bit_dac_0[0].switch2n_3v3_0.VOUTH 1.98e-19
C143 2_bit_dac_0[0].switch2n_3v3_0.R_H 2_bit_dac_0[0].D0 0.13f
C144 2_bit_dac_0[0].VOUT 2_bit_dac_0[0].switch2n_3v3_0.VREFH 2.34e-21
C145 2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.128f
C146 D0_BUF 2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.472f
C147 2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0927f
C148 2_bit_dac_0[1].VREFH 2_bit_dac_0[0].D0 1.06f
C149 2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 2_bit_dac_0[0].switch2n_3v3_0.R_H 0.00819f
C150 2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.511f
C151 2_bit_dac_0[0].D1 2_bit_dac_0[0].VOUT 0.00692f
C152 a_1438_406# 2_bit_dac_0[1].switch2n_3v3_0.R_L 1.29e-19
C153 2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2_bit_dac_0[0].switch2n_3v3_0.R_H 8.92e-19
C154 2_bit_dac_0[0].switch2n_3v3_0.R_H VREFL 3.7e-20
C155 2_bit_dac_0[0].switch2n_3v3_0.R_H D0 1.48e-19
C156 2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 2_bit_dac_0[1].switch2n_3v3_0.R_L 4.25e-19
C157 D0_BUF 2_bit_dac_0[0].D1 0.0179f
C158 VOUT switch_n_3v3_1.D7 0.00684f
C159 D2_BUF VOUT 0.0718f
C160 2_bit_dac_0[0].switch2n_3v3_0.VOUTL 2_bit_dac_0[0].VOUT 0.302f
C161 2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2_bit_dac_0[1].VREFH 3.38e-20
C162 2_bit_dac_0[1].VREFH VREFL 0.0988f
C163 2_bit_dac_0[1].VREFH D0 0.00555f
C164 D0_BUF 2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.38f
C165 2_bit_dac_0[0].switch2n_3v3_0.R_H 2_bit_dac_0[1].switch2n_3v3_0.R_L 0.00368f
C166 D2 switch_n_3v3_1.D5 0.0322f
C167 switch_n_3v3_1.D7 2_bit_dac_0[0].VOUT 0.0265f
C168 D2_BUF 2_bit_dac_0[0].VOUT 0.546f
C169 2_bit_dac_0[1].VREFH 2_bit_dac_0[1].switch2n_3v3_0.R_L 0.00183f
C170 a_1438_406# 2_bit_dac_0[1].switch2n_3v3_0.VREFH 9.57e-20
C171 a_1438_406# VREFH 2.68e-20
C172 2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 2_bit_dac_0[1].switch2n_3v3_0.VREFH 5.89e-20
C173 D0_BUF 2_bit_dac_0[0].D0 0.124f
C174 2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 2_bit_dac_0[0].VOUT 0.229f
C175 2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2_bit_dac_0[0].VOUT 0.051f
C176 switch_n_3v3_1.DX_ 2_bit_dac_0[1].VOUT 0.125f
C177 2_bit_dac_0[0].switch2n_3v3_0.VOUTH 2_bit_dac_0[1].switch2n_3v3_0.VREFH 5.55e-20
C178 2_bit_dac_0[0].D1 D2 0.0026f
C179 D0_BUF 2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5.84e-19
C180 2_bit_dac_0[0].switch2n_3v3_0.R_H 2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.0018f
C181 VREFH 2_bit_dac_0[0].switch2n_3v3_0.R_H 0.0579f
C182 D0_BUF VREFL 4.97e-19
C183 D0_BUF 2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00349f
C184 2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ switch_n_3v3_1.D4 2.51e-19
C185 2_bit_dac_0[1].switch2n_3v3_0.VREFH 2_bit_dac_0[1].VREFH 0.0124f
C186 VREFH 2_bit_dac_0[1].VREFH 0.0988f
C187 D1 2_bit_dac_0[1].VOUT 0.0057f
C188 2_bit_dac_0[0].switch2n_3v3_0.VOUTH switch_n_3v3_1.D4 7.43e-20
C189 a_1438_406# 2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0892f
C190 D0_BUF 2_bit_dac_0[1].switch2n_3v3_0.R_L 1.9e-19
C191 a_1438_406# 2_bit_dac_0[0].switch2n_3v3_0.R_H 0.397f
C192 2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.00143f
C193 D2 switch_n_3v3_1.D7 0.0518f
C194 switch_n_3v3_1.D3 2_bit_dac_0[1].VOUT 0.0121f
C195 D2_BUF D2 0.0694f
C196 switch_n_3v3_1.DX_ switch_n_3v3_1.D6 2.54e-19
C197 VCC 2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.622f
C198 a_1438_406# 2_bit_dac_0[1].VREFH 0.337f
C199 D1_BUF VCC 0.317f
C200 2_bit_dac_0[0].switch2n_3v3_0.R_H 2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.394f
C201 switch_n_3v3_1.D4 VOUT 1.74e-20
C202 2_bit_dac_0[1].switch2n_3v3_0.VOUTL D2 0.0701f
C203 D1 a_1438_1634# 0.003f
C204 D0_BUF 2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.00105f
C205 D0_BUF VREFH 0.281f
C206 2_bit_dac_0[0].switch2n_3v3_0.R_H 2_bit_dac_0[1].VREFH 0.138f
C207 2_bit_dac_0[0].switch2n_3v3_0.R_L 2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0923f
C208 switch_n_3v3_1.D4 2_bit_dac_0[0].VOUT 0.02f
C209 2_bit_dac_0[1].switch2n_3v3_0.R_H 2_bit_dac_0[1].VOUT 3.62e-20
C210 2_bit_dac_0[0].switch2n_3v3_0.R_L 2_bit_dac_0[0].D1 0.00319f
C211 2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 2_bit_dac_0[0].VOUT 0.0035f
C212 D1_BUF 2_bit_dac_0[1].switch2n_3v3_0.VOUTH 1.85e-19
C213 a_1438_406# D0_BUF 0.325f
C214 2_bit_dac_0[0].switch2n_3v3_0.R_L 2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.189f
C215 2_bit_dac_0[0].switch2n_3v3_0.VOUTH 2_bit_dac_0[0].VOUT 0.504f
C216 2_bit_dac_0[0].switch2n_3v3_0.R_H 2_bit_dac_0[0].VOUT 3.62e-20
C217 D0_BUF 2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.347f
C218 D0_BUF 2_bit_dac_0[0].switch2n_3v3_0.R_H 0.24f
C219 2_bit_dac_0[1].VOUT switch_n_3v3_1.D5 0.0234f
C220 2_bit_dac_0[1].switch2n_3v3_0.R_H a_1438_1634# 0.397f
C221 2_bit_dac_0[0].switch2n_3v3_0.R_L 2_bit_dac_0[0].D0 0.265f
C222 D0_BUF 2_bit_dac_0[1].VREFH 0.538f
C223 VOUT 2_bit_dac_0[0].VOUT 0.314f
C224 D2 switch_n_3v3_1.D4 0.0568f
C225 2_bit_dac_0[0].switch2n_3v3_0.R_L 2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 4.25e-19
C226 2_bit_dac_0[0].switch2n_3v3_0.R_L VREFL 0.005f
C227 2_bit_dac_0[0].switch2n_3v3_0.R_L D0 9.68e-20
C228 2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ D2 0.0222f
C229 2_bit_dac_0[0].D1 2_bit_dac_0[1].VOUT 0.0757f
C230 switch_n_3v3_1.D5 switch_n_3v3_1.D6 0.67f
C231 2_bit_dac_0[1].VOUT 2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00473f
C232 D0_BUF 2_bit_dac_0[0].VOUT 2.29e-20
C233 switch_n_3v3_1.DX_ VCC 0.698f
C234 2_bit_dac_0[0].switch2n_3v3_0.VREFH a_1438_1634# 0.0331f
C235 2_bit_dac_0[1].VOUT 2_bit_dac_0[0].D0 2.29e-20
C236 2_bit_dac_0[1].VOUT switch_n_3v3_1.D7 0.036f
C237 D2_BUF 2_bit_dac_0[1].VOUT 0.177f
C238 D1 VCC 0.459f
C239 2_bit_dac_0[0].D1 a_1438_1634# 6.04e-19
C240 2_bit_dac_0[0].D1 switch_n_3v3_1.D6 1.79e-20
C241 D2 VOUT 1.75e-20
C242 2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1438_1634# 2.93e-19
C243 2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 2_bit_dac_0[1].VOUT 1.06e-19
C244 2_bit_dac_0[0].switch2n_3v3_0.R_L VREFH 7.62e-19
C245 switch_n_3v3_1.D3 VCC 0.0539f
C246 2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2_bit_dac_0[1].VOUT 0.303f
C247 switch_n_3v3_1.DX_ 2_bit_dac_0[1].switch2n_3v3_0.VOUTH 9.82e-21
C248 D2 2_bit_dac_0[0].VOUT 2.96e-19
C249 a_1438_1634# 2_bit_dac_0[0].D0 0.325f
C250 switch_n_3v3_1.D6 switch_n_3v3_1.D7 0.67f
C251 D2_BUF switch_n_3v3_1.D6 0.0293f
C252 2_bit_dac_0[0].switch2n_3v3_0.R_L a_1438_406# 0.403f
C253 D1 2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0778f
C254 2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1438_1634# 0.296f
C255 VREFL a_1438_1634# 0.337f
C256 2_bit_dac_0[1].switch2n_3v3_0.VOUTL switch_n_3v3_1.D6 0.00202f
C257 D0 a_1438_1634# 0.0975f
C258 switch_n_3v3_1.D3 2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00189f
C259 2_bit_dac_0[0].switch2n_3v3_0.R_L 2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0018f
C260 2_bit_dac_0[0].switch2n_3v3_0.R_L 2_bit_dac_0[0].switch2n_3v3_0.R_H 0.805f
C261 2_bit_dac_0[1].switch2n_3v3_0.R_H VCC 0.312f
C262 2_bit_dac_0[1].VOUT 2_bit_dac_0[1].switch2n_3v3_0.VREFH 2.34e-21
C263 2_bit_dac_0[0].switch2n_3v3_0.R_L 2_bit_dac_0[1].VREFH 0.482f
C264 2_bit_dac_0[1].switch2n_3v3_0.R_L a_1438_1634# 0.403f
C265 switch_n_3v3_1.D4 2_bit_dac_0[1].VOUT 0.0268f
C266 VCC switch_n_3v3_1.D5 0.0583f
C267 2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 2_bit_dac_0[1].VOUT 0.229f
C268 2_bit_dac_0[1].switch2n_3v3_0.R_H 2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.394f
C269 2_bit_dac_0[1].switch2n_3v3_0.VREFH a_1438_1634# 0.175f
C270 VCC 2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.835f
C271 2_bit_dac_0[0].switch2n_3v3_0.VOUTH 2_bit_dac_0[1].VOUT 6.14e-19
C272 2_bit_dac_0[0].switch2n_3v3_0.R_L D0_BUF 0.315f
C273 2_bit_dac_0[0].D1 VCC 0.793f
C274 a_1438_406# a_1438_1634# 0.00981f
C275 VCC 2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.243f
C276 2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ switch_n_3v3_1.D6 1.72e-19
C277 2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ a_1438_1634# 1.21e-20
C278 2_bit_dac_0[1].switch2n_3v3_0.VOUTH switch_n_3v3_1.D5 8.21e-19
C279 2_bit_dac_0[1].VOUT VOUT 0.537f
C280 2_bit_dac_0[0].switch2n_3v3_0.VOUTH switch_n_3v3_1.D6 3.83e-20
C281 2_bit_dac_0[0].switch2n_3v3_0.R_H a_1438_1634# 4.09e-19
C282 VCC 2_bit_dac_0[0].D0 1.18f
C283 VCC switch_n_3v3_1.D7 0.145f
C284 D1_BUF 2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.00375f
C285 D2_BUF VCC 0.337f
C286 2_bit_dac_0[0].D1 2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.176f
C287 2_bit_dac_0[1].VREFH a_1438_1634# 2.68e-20
C288 2_bit_dac_0[1].VOUT 2_bit_dac_0[0].VOUT 0.349f
C289 2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VCC 0.697f
C290 D1_BUF 2_bit_dac_0[0].D1 0.0392f
C291 switch_n_3v3_1.DX_ switch_n_3v3_1.D3 1.03e-19
C292 2_bit_dac_0[0].switch2n_3v3_0.VOUTL 2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00163f
C293 2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC 0.312f
C294 VCC VREFL 0.144f
C295 VCC D0 0.407f
C296 VOUT switch_n_3v3_1.D6 2.29e-20
C297 D1_BUF 2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.632f
C298 switch_n_3v3_1.D3 D1 2.93e-21
C299 VCC 2_bit_dac_0[1].switch2n_3v3_0.R_L 0.291f
C300 2_bit_dac_0[1].switch2n_3v3_0.VOUTH 2_bit_dac_0[0].D0 0.347f
C301 2_bit_dac_0[1].switch2n_3v3_0.VOUTH switch_n_3v3_1.D7 4.71e-19
C302 D2_BUF 2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00476f
C303 switch_n_3v3_1.D6 2_bit_dac_0[0].VOUT 0.0199f
C304 D0_BUF a_1438_1634# 0.00365f
C305 2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 2_bit_dac_0[1].switch2n_3v3_0.VOUTH 1.46e-19
C306 2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.579f
C307 2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ D1_BUF 0.219f
C308 D2 2_bit_dac_0[1].VOUT 0.137f
C309 D1_BUF 2_bit_dac_0[1].switch2n_3v3_0.VOUTL 4.15e-19
C310 VCC 2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.836f
C311 VREFH VCC 0.0022f
C312 2_bit_dac_0[1].switch2n_3v3_0.VOUTH 2_bit_dac_0[1].switch2n_3v3_0.R_L 0.0018f
C313 D1 2_bit_dac_0[1].switch2n_3v3_0.R_H 0.037f
C314 VCC switch_n_3v3_1.D4 0.0574f
C315 D2 switch_n_3v3_1.D6 0.0325f
C316 a_1438_406# VCC 0.706f
C317 switch_n_3v3_1.DX_ switch_n_3v3_1.D5 1.8e-19
C318 2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VCC 0.714f
C319 2_bit_dac_0[1].switch2n_3v3_0.VREFH 2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.236f
C320 VCC 2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.603f
C321 2_bit_dac_0[0].switch2n_3v3_0.R_H VCC 0.307f
C322 switch_n_3v3_1.DX_ 2_bit_dac_0[0].D1 1.34e-20
C323 VCC 2_bit_dac_0[1].VREFH 0.135f
C324 switch_n_3v3_1.D4 2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00116f
C325 2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0927f
C326 VCC VOUT 0.282f
C327 a_1438_406# D1_BUF 6.04e-19
C328 D1 2_bit_dac_0[0].D1 0.0384f
C329 2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ D1_BUF 6.11e-19
R0 VSS.n982 VSS.n981 12274.8
R1 VSS.n981 VSS.n980 12232.2
R2 VSS.n841 VSS.t35 4305.17
R3 VSS.n524 VSS.t3 2804.58
R4 VSS.n523 VSS.t28 2770.93
R5 VSS.n525 VSS.n524 2671.38
R6 VSS.n841 VSS.n840 2406.66
R7 VSS.t7 VSS.n622 2349.66
R8 VSS.t18 VSS.t7 2304.76
R9 VSS.t6 VSS.n673 1937.11
R10 VSS.n842 VSS.n841 1896.55
R11 VSS.t31 VSS.t6 1892.74
R12 VSS.t32 VSS.n842 1791.5
R13 VSS.t22 VSS.t32 1683.22
R14 VSS.n45 VSS.t10 1560.55
R15 VSS.n674 VSS.t18 1331.97
R16 VSS.n674 VSS.t31 1093.85
R17 VSS.n843 VSS.t22 1045.79
R18 VSS.n676 VSS.n675 1017.62
R19 VSS.n675 VSS.n674 772.908
R20 VSS.n354 VSS.t20 758.37
R21 VSS.t20 VSS.t2 746.255
R22 VSS.n981 VSS.t15 447.884
R23 VSS.n933 VSS.n930 332.558
R24 VSS.n129 VSS.n128 292.5
R25 VSS.t15 VSS.t19 275.897
R26 VSS.n523 VSS.t11 269.807
R27 VSS.t21 VSS.t12 261.565
R28 VSS.t19 VSS.t21 257.981
R29 VSS.n609 VSS.t16 239.457
R30 VSS.n660 VSS.t29 198.87
R31 VSS.n842 VSS.t23 188.758
R32 VSS.n106 VSS.n105 121.799
R33 VSS.n134 VSS.n133 121.799
R34 VSS.n590 VSS.n589 112.246
R35 VSS.n561 VSS.n560 112.246
R36 VSS.n87 VSS.n86 106.575
R37 VSS.n150 VSS.t33 106.575
R38 VSS.n910 VSS.n909 102.326
R39 VSS.n933 VSS.n932 102.326
R40 VSS.n85 VSS.t8 98.9624
R41 VSS.n608 VSS.n607 97.2794
R42 VSS.t4 VSS.n541 97.2794
R43 VSS.n640 VSS.n639 93.2208
R44 VSS.n814 VSS.n813 93.2208
R45 VSS.n66 VSS.n65 91.35
R46 VSS.n181 VSS.n180 91.35
R47 VSS.n891 VSS.n890 89.5354
R48 VSS.n203 VSS.t26 89.5354
R49 VSS.n889 VSS.t24 83.14
R50 VSS.n425 VSS.n424 82.3134
R51 VSS.n522 VSS.n521 82.3134
R52 VSS.n659 VSS.n658 80.7915
R53 VSS.t13 VSS.n285 80.7915
R54 VSS.n135 VSS.n129 80.0317
R55 VSS.n934 VSS.n927 80.0317
R56 VSS.n261 VSS.n260 76.7447
R57 VSS.n224 VSS.n223 76.7447
R58 VSS.n47 VSS.n46 76.1251
R59 VSS.n984 VSS.n983 76.1251
R60 VSS.n373 VSS.t0 75.1106
R61 VSS.n624 VSS.n623 68.3621
R62 VSS.n278 VSS.n277 68.3621
R63 VSS.n845 VSS.n844 63.954
R64 VSS.n979 VSS.n978 63.954
R65 VSS.n46 VSS.n45 53.2877
R66 VSS.n983 VSS.n982 53.2877
R67 VSS.n679 VSS.t37 46.866
R68 VSS.n837 VSS.t14 46.863
R69 VSS.n528 VSS.t5 46.863
R70 VSS.n649 VSS.t30 46.8459
R71 VSS.n599 VSS.t17 46.8459
R72 VSS.n380 VSS.t1 46.8455
R73 VSS.n168 VSS.t34 46.8085
R74 VSS.n233 VSS.t27 46.8085
R75 VSS.n96 VSS.t9 46.808
R76 VSS.n900 VSS.t25 46.808
R77 VSS.n622 VSS.n425 44.8985
R78 VSS.n525 VSS.n522 44.8985
R79 VSS.n844 VSS.n843 44.7679
R80 VSS.n980 VSS.n979 44.7679
R81 VSS.n65 VSS.n64 38.0628
R82 VSS.n180 VSS.n179 38.0628
R83 VSS.n673 VSS.n624 37.2886
R84 VSS.n840 VSS.n278 37.2886
R85 VSS.n389 VSS.n388 36.3441
R86 VSS.n701 VSS.n700 36.3441
R87 VSS.n524 VSS.n523 33.5883
R88 VSS.n260 VSS.n259 31.9772
R89 VSS.n223 VSS.n222 31.9772
R90 VSS.n372 VSS.n371 31.4983
R91 VSS.n410 VSS.n409 31.4983
R92 VSS.n609 VSS.n608 29.9325
R93 VSS.n542 VSS.t4 29.9325
R94 VSS.n353 VSS.n352 26.6525
R95 VSS.n423 VSS.n422 26.6525
R96 VSS.n660 VSS.n659 24.8593
R97 VSS.n286 VSS.t13 24.8593
R98 VSS.n107 VSS.n103 24.6255
R99 VSS.n135 VSS.n131 24.6255
R100 VSS.n911 VSS.n907 24.6255
R101 VSS.n934 VSS.n929 24.6255
R102 VSS.n86 VSS.n85 22.8379
R103 VSS.t33 VSS.n149 22.8379
R104 VSS.n88 VSS.n84 21.5474
R105 VSS.n151 VSS.n148 21.5474
R106 VSS.n892 VSS.n888 21.5474
R107 VSS.n204 VSS.n201 21.5474
R108 VSS.n638 VSS.n637 21.1076
R109 VSS.n812 VSS.n811 21.1076
R110 VSS.n387 VSS.n386 21.1076
R111 VSS.n699 VSS.n698 21.1076
R112 VSS.n588 VSS.n587 21.1076
R113 VSS.n559 VSS.n558 21.1076
R114 VSS.n890 VSS.n889 19.1865
R115 VSS.t26 VSS.n202 19.1865
R116 VSS.n67 VSS.n63 18.4693
R117 VSS.n182 VSS.n178 18.4693
R118 VSS.n262 VSS.n258 18.4693
R119 VSS.n225 VSS.n221 18.4693
R120 VSS.n657 VSS.n656 18.2934
R121 VSS.n284 VSS.n283 18.2934
R122 VSS.n370 VSS.n369 18.2934
R123 VSS.n408 VSS.n407 18.2934
R124 VSS.n606 VSS.n605 18.2934
R125 VSS.n540 VSS.n539 18.2934
R126 VSS.n626 VSS.n625 15.4791
R127 VSS.n280 VSS.n279 15.4791
R128 VSS.n351 VSS.n350 15.4791
R129 VSS.n421 VSS.n420 15.4791
R130 VSS.n427 VSS.n426 15.4791
R131 VSS.n520 VSS.n519 15.4791
R132 VSS.n48 VSS.n44 15.3911
R133 VSS.n985 VSS.n188 15.3911
R134 VSS.n846 VSS.n276 15.3911
R135 VSS.n977 VSS.n190 15.3911
R136 VSS.n591 VSS.n590 14.9665
R137 VSS.n562 VSS.n561 14.9665
R138 VSS.n354 VSS.n353 14.5379
R139 VSS.n676 VSS.n423 14.5379
R140 VSS.n641 VSS.n640 12.4299
R141 VSS.n815 VSS.n814 12.4299
R142 VSS.n373 VSS.n372 9.69213
R143 VSS.n672 VSS.n671 9.38145
R144 VSS.n358 VSS.n355 9.38145
R145 VSS.n621 VSS.n620 9.38145
R146 VSS.n564 VSS.n563 9.3005
R147 VSS.n563 VSS.n562 9.3005
R148 VSS.n593 VSS.n592 9.3005
R149 VSS.n592 VSS.n591 9.3005
R150 VSS.n611 VSS.n610 9.3005
R151 VSS.n610 VSS.n609 9.3005
R152 VSS.n544 VSS.n543 9.3005
R153 VSS.n543 VSS.n542 9.3005
R154 VSS.n527 VSS.n526 9.3005
R155 VSS.n526 VSS.n525 9.3005
R156 VSS.n622 VSS.n621 9.3005
R157 VSS.n183 VSS.n182 9.3005
R158 VSS.n182 VSS.n181 9.3005
R159 VSS.n152 VSS.n151 9.3005
R160 VSS.n151 VSS.n150 9.3005
R161 VSS.n136 VSS.n135 9.3005
R162 VSS.n135 VSS.n134 9.3005
R163 VSS.n89 VSS.n88 9.3005
R164 VSS.n88 VSS.n87 9.3005
R165 VSS.n108 VSS.n107 9.3005
R166 VSS.n107 VSS.n106 9.3005
R167 VSS.n986 VSS.n985 9.3005
R168 VSS.n985 VSS.n984 9.3005
R169 VSS.n49 VSS.n48 9.3005
R170 VSS.n48 VSS.n47 9.3005
R171 VSS.n68 VSS.n67 9.3005
R172 VSS.n67 VSS.n66 9.3005
R173 VSS.n704 VSS.n703 9.3005
R174 VSS.n703 VSS.n702 9.3005
R175 VSS.n392 VSS.n391 9.3005
R176 VSS.n391 VSS.n390 9.3005
R177 VSS.n375 VSS.n374 9.3005
R178 VSS.n374 VSS.n373 9.3005
R179 VSS.n413 VSS.n412 9.3005
R180 VSS.n412 VSS.n411 9.3005
R181 VSS.n678 VSS.n677 9.3005
R182 VSS.n677 VSS.n676 9.3005
R183 VSS.n355 VSS.n354 9.3005
R184 VSS.n817 VSS.n816 9.3005
R185 VSS.n816 VSS.n815 9.3005
R186 VSS.n643 VSS.n642 9.3005
R187 VSS.n642 VSS.n641 9.3005
R188 VSS.n662 VSS.n661 9.3005
R189 VSS.n661 VSS.n660 9.3005
R190 VSS.n288 VSS.n287 9.3005
R191 VSS.n287 VSS.n286 9.3005
R192 VSS.n839 VSS.n838 9.3005
R193 VSS.n840 VSS.n839 9.3005
R194 VSS.n673 VSS.n672 9.3005
R195 VSS.n847 VSS.n846 9.3005
R196 VSS.n846 VSS.n845 9.3005
R197 VSS.n263 VSS.n262 9.3005
R198 VSS.n262 VSS.n261 9.3005
R199 VSS.n893 VSS.n892 9.3005
R200 VSS.n892 VSS.n891 9.3005
R201 VSS.n912 VSS.n911 9.3005
R202 VSS.n911 VSS.n910 9.3005
R203 VSS.n935 VSS.n934 9.3005
R204 VSS.n934 VSS.n933 9.3005
R205 VSS.n205 VSS.n204 9.3005
R206 VSS.n204 VSS.n203 9.3005
R207 VSS.n226 VSS.n225 9.3005
R208 VSS.n225 VSS.n224 9.3005
R209 VSS.n977 VSS.n976 9.3005
R210 VSS.n978 VSS.n977 9.3005
R211 VSS.n576 VSS.n575 9.15497
R212 VSS.n575 VSS.n574 9.15497
R213 VSS.n403 VSS.n402 9.15497
R214 VSS.n402 VSS.n401 9.15497
R215 VSS.n801 VSS.n800 9.15497
R216 VSS.n800 VSS.n799 9.15497
R217 VSS.n672 VSS.n626 8.44336
R218 VSS.n839 VSS.n280 8.44336
R219 VSS.n355 VSS.n351 8.44336
R220 VSS.n677 VSS.n421 8.44336
R221 VSS.n621 VSS.n427 8.44336
R222 VSS.n526 VSS.n520 8.44336
R223 VSS.n63 VSS.n62 7.69581
R224 VSS.n178 VSS.n177 7.69581
R225 VSS.n258 VSS.n257 7.69581
R226 VSS.n221 VSS.n220 7.69581
R227 VSS.n105 VSS.n104 7.61296
R228 VSS.n133 VSS.n132 7.61296
R229 VSS.n411 VSS.t36 7.26922
R230 VSS.n909 VSS.n908 6.39585
R231 VSS.n932 VSS.n931 6.39585
R232 VSS.n661 VSS.n657 5.62907
R233 VSS.n287 VSS.n284 5.62907
R234 VSS.n374 VSS.n370 5.62907
R235 VSS.n412 VSS.n408 5.62907
R236 VSS.n610 VSS.n606 5.62907
R237 VSS.n543 VSS.n540 5.62907
R238 VSS.n188 VSS.n187 5.33568
R239 VSS.n44 VSS.n43 5.33568
R240 VSS.n276 VSS.n275 5.33568
R241 VSS.n190 VSS.n189 5.33568
R242 VSS.n390 VSS.n389 4.84631
R243 VSS.n702 VSS.n701 4.84631
R244 VSS.n84 VSS.n83 4.61769
R245 VSS.n148 VSS.n147 4.61769
R246 VSS.n888 VSS.n887 4.61769
R247 VSS.n201 VSS.n200 4.61769
R248 VSS.n645 VSS.n644 4.5005
R249 VSS.n820 VSS.n819 4.5005
R250 VSS.n394 VSS.n393 4.5005
R251 VSS.n707 VSS.n706 4.5005
R252 VSS.n52 VSS.n51 4.5005
R253 VSS.n72 VSS.n71 4.5005
R254 VSS.n111 VSS.n110 4.5005
R255 VSS.n93 VSS.n92 4.5005
R256 VSS.n154 VSS.n153 4.5005
R257 VSS.n138 VSS.n137 4.5005
R258 VSS.n117 VSS.n116 4.5005
R259 VSS.n121 VSS.n120 4.5005
R260 VSS.n988 VSS.n987 4.5005
R261 VSS.n548 VSS.n547 4.5005
R262 VSS.n595 VSS.n594 4.5005
R263 VSS.n567 VSS.n566 4.5005
R264 VSS.n897 VSS.n896 4.5005
R265 VSS.n850 VSS.n849 4.5005
R266 VSS.n267 VSS.n266 4.5005
R267 VSS.n915 VSS.n914 4.5005
R268 VSS.n921 VSS.n920 4.5005
R269 VSS.n943 VSS.n942 4.5005
R270 VSS.n937 VSS.n936 4.5005
R271 VSS.n207 VSS.n206 4.5005
R272 VSS.n228 VSS.n227 4.5005
R273 VSS.n975 VSS.n974 4.5005
R274 VSS.n528 VSS.n527 3.69976
R275 VSS.n838 VSS.n837 3.69976
R276 VSS.n679 VSS.n678 3.69922
R277 VSS.n186 VSS.n185 3.29193
R278 VSS.n429 VSS.n428 3.29193
R279 VSS.n292 VSS.n291 3.2005
R280 VSS.n417 VSS.n416 3.2005
R281 VSS.n577 VSS.n576 3.03311
R282 VSS.n612 VSS.n611 3.03311
R283 VSS.n404 VSS.n403 3.03311
R284 VSS.n376 VSS.n375 3.03311
R285 VSS.n802 VSS.n801 3.03311
R286 VSS.n663 VSS.n662 3.03311
R287 VSS.n642 VSS.n638 2.81479
R288 VSS.n816 VSS.n812 2.81479
R289 VSS.n391 VSS.n387 2.81479
R290 VSS.n703 VSS.n699 2.81479
R291 VSS.n592 VSS.n588 2.81479
R292 VSS.n563 VSS.n559 2.81479
R293 VSS.t36 VSS.n410 2.42341
R294 VSS.n174 VSS.n173 2.37764
R295 VSS.n1008 VSS.n1007 2.27266
R296 VSS.n116 VSS.n115 2.01193
R297 VSS.n920 VSS.n919 2.01193
R298 VSS.n671 VSS.n670 1.98071
R299 VSS.n359 VSS.n358 1.98071
R300 VSS.n620 VSS.n619 1.98071
R301 VSS.n662 VSS.n653 1.55479
R302 VSS.n375 VSS.n366 1.55479
R303 VSS.n103 VSS.n102 1.53956
R304 VSS.n131 VSS.n130 1.53956
R305 VSS.n907 VSS.n906 1.53956
R306 VSS.n929 VSS.n928 1.53956
R307 VSS.n715 VSS.n714 1.5005
R308 VSS.n290 VSS.n289 1.46336
R309 VSS.n415 VSS.n414 1.46336
R310 VSS.n108 VSS.n101 1.46336
R311 VSS.n136 VSS.n127 1.46336
R312 VSS.n547 VSS.n546 1.46336
R313 VSS.n912 VSS.n905 1.46336
R314 VSS.n935 VSS.n926 1.46336
R315 VSS.n644 VSS.n634 1.37193
R316 VSS.n636 VSS.n635 1.37193
R317 VSS.n810 VSS.n809 1.37193
R318 VSS.n819 VSS.n818 1.37193
R319 VSS.n393 VSS.n383 1.37193
R320 VSS.n385 VSS.n384 1.37193
R321 VSS.n697 VSS.n696 1.37193
R322 VSS.n706 VSS.n705 1.37193
R323 VSS.n594 VSS.n584 1.37193
R324 VSS.n586 VSS.n585 1.37193
R325 VSS.n557 VSS.n556 1.37193
R326 VSS.n566 VSS.n565 1.37193
R327 VSS.n89 VSS.n82 1.2805
R328 VSS.n893 VSS.n886 1.2805
R329 VSS.n205 VSS.n199 1.2805
R330 VSS.n655 VSS.n654 1.18907
R331 VSS.n282 VSS.n281 1.18907
R332 VSS.n368 VSS.n367 1.18907
R333 VSS.n406 VSS.n405 1.18907
R334 VSS.n604 VSS.n603 1.18907
R335 VSS.n538 VSS.n537 1.18907
R336 VSS.n460 VSS.n459 1.13717
R337 VSS.n511 VSS.n510 1.13717
R338 VSS.n345 VSS.n344 1.13717
R339 VSS.n739 VSS.n738 1.13717
R340 VSS.n757 VSS.n756 1.13717
R341 VSS.n794 VSS.n793 1.13717
R342 VSS.n802 VSS.n798 1.1255
R343 VSS.n577 VSS.n515 1.1255
R344 VSS.n68 VSS.n61 1.09764
R345 VSS.n184 VSS.n183 1.09764
R346 VSS.n263 VSS.n256 1.09764
R347 VSS.n226 VSS.n219 1.09764
R348 VSS.n949 VSS.n944 1.04225
R349 VSS.n628 VSS.n627 1.00621
R350 VSS.n293 VSS.n292 1.00621
R351 VSS.n357 VSS.n356 1.00621
R352 VSS.n418 VSS.n417 1.00621
R353 VSS.n71 VSS.n68 1.00621
R354 VSS.n70 VSS.n69 1.00621
R355 VSS.n137 VSS.n125 1.00621
R356 VSS.n430 VSS.n429 1.00621
R357 VSS.n517 VSS.n516 1.00621
R358 VSS.n266 VSS.n263 1.00621
R359 VSS.n265 VSS.n264 1.00621
R360 VSS.n936 VSS.n924 1.00621
R361 VSS.n51 VSS.n49 0.914786
R362 VSS.n110 VSS.n109 0.914786
R363 VSS.n116 VSS.n114 0.914786
R364 VSS.n175 VSS.n174 0.914786
R365 VSS.n183 VSS.n176 0.914786
R366 VSS.n987 VSS.n986 0.914786
R367 VSS.n849 VSS.n847 0.914786
R368 VSS.n914 VSS.n913 0.914786
R369 VSS.n920 VSS.n918 0.914786
R370 VSS.n217 VSS.n216 0.914786
R371 VSS.n227 VSS.n226 0.914786
R372 VSS.n976 VSS.n975 0.914786
R373 VSS.n990 VSS.n989 0.908949
R374 VSS.n973 VSS.n972 0.908949
R375 VSS.n42 VSS.n41 0.908879
R376 VSS.n852 VSS.n851 0.908879
R377 VSS.n1001 VSS.n1000 0.853
R378 VSS.n868 VSS.n867 0.853
R379 VSS.n950 VSS.n949 0.853
R380 VSS.n962 VSS.n961 0.853
R381 VSS.n92 VSS.n89 0.823357
R382 VSS.n91 VSS.n90 0.823357
R383 VSS.n120 VSS.n119 0.823357
R384 VSS.n153 VSS.n146 0.823357
R385 VSS.n896 VSS.n893 0.823357
R386 VSS.n895 VSS.n894 0.823357
R387 VSS.n942 VSS.n941 0.823357
R388 VSS.n206 VSS.n197 0.823357
R389 VSS.n92 VSS.n91 0.731929
R390 VSS.n146 VSS.n145 0.731929
R391 VSS.n153 VSS.n152 0.731929
R392 VSS.n896 VSS.n895 0.731929
R393 VSS.n197 VSS.n196 0.731929
R394 VSS.n206 VSS.n205 0.731929
R395 VSS.n51 VSS.n50 0.6405
R396 VSS.n110 VSS.n108 0.6405
R397 VSS.n176 VSS.n175 0.6405
R398 VSS.n987 VSS.n186 0.6405
R399 VSS.n849 VSS.n848 0.6405
R400 VSS.n914 VSS.n912 0.6405
R401 VSS.n227 VSS.n217 0.6405
R402 VSS.n975 VSS.n191 0.6405
R403 VSS.n71 VSS.n70 0.549071
R404 VSS.n137 VSS.n136 0.549071
R405 VSS.n266 VSS.n265 0.549071
R406 VSS.n936 VSS.n935 0.549071
R407 VSS VSS.n502 0.517836
R408 VSS VSS.n785 0.517836
R409 VSS.n671 VSS.n628 0.465127
R410 VSS.n358 VSS.n357 0.465127
R411 VSS.n620 VSS.n430 0.465127
R412 VSS.n294 VSS.n293 0.457643
R413 VSS.n419 VSS.n418 0.457643
R414 VSS.n61 VSS.n60 0.457643
R415 VSS.n185 VSS.n184 0.457643
R416 VSS.n518 VSS.n517 0.457643
R417 VSS.n256 VSS.n255 0.457643
R418 VSS.n219 VSS.n218 0.457643
R419 VSS.n662 VSS.n655 0.366214
R420 VSS.n288 VSS.n282 0.366214
R421 VSS.n375 VSS.n368 0.366214
R422 VSS.n413 VSS.n406 0.366214
R423 VSS.n611 VSS.n604 0.366214
R424 VSS.n544 VSS.n538 0.366214
R425 VSS.n450 VSS 0.301636
R426 VSS.n335 VSS 0.301636
R427 VSS VSS.n1006 0.300964
R428 VSS VSS.n0 0.300964
R429 VSS.n747 VSS 0.29425
R430 VSS.n82 VSS.n81 0.274786
R431 VSS.n173 VSS.n172 0.274786
R432 VSS.n886 VSS.n885 0.274786
R433 VSS.n199 VSS.n198 0.274786
R434 VSS VSS.n746 0.206964
R435 VSS.n644 VSS.n643 0.183357
R436 VSS.n643 VSS.n636 0.183357
R437 VSS.n817 VSS.n810 0.183357
R438 VSS.n819 VSS.n817 0.183357
R439 VSS.n393 VSS.n392 0.183357
R440 VSS.n392 VSS.n385 0.183357
R441 VSS.n704 VSS.n697 0.183357
R442 VSS.n706 VSS.n704 0.183357
R443 VSS.n594 VSS.n593 0.183357
R444 VSS.n593 VSS.n586 0.183357
R445 VSS.n564 VSS.n557 0.183357
R446 VSS.n566 VSS.n564 0.183357
R447 VSS.n1007 VSS 0.107929
R448 VSS VSS.n1008 0.107929
R449 VSS.n503 VSS 0.107593
R450 VSS.n786 VSS 0.107593
R451 VSS.n289 VSS.n288 0.0919286
R452 VSS.n291 VSS.n290 0.0919286
R453 VSS.n838 VSS.n294 0.0919286
R454 VSS.n414 VSS.n413 0.0919286
R455 VSS.n416 VSS.n415 0.0919286
R456 VSS.n678 VSS.n419 0.0919286
R457 VSS.n101 VSS.n100 0.0919286
R458 VSS.n127 VSS.n126 0.0919286
R459 VSS.n547 VSS.n544 0.0919286
R460 VSS.n546 VSS.n545 0.0919286
R461 VSS.n527 VSS.n518 0.0919286
R462 VSS.n905 VSS.n904 0.0919286
R463 VSS.n926 VSS.n925 0.0919286
R464 VSS.n453 VSS.n452 0.024
R465 VSS.n506 VSS.n505 0.024
R466 VSS.n338 VSS.n337 0.024
R467 VSS.n744 VSS.n743 0.024
R468 VSS.n750 VSS.n749 0.024
R469 VSS.n789 VSS.n788 0.024
R470 VSS.n630 VSS.n629 0.0228214
R471 VSS.n805 VSS.n804 0.0228214
R472 VSS.n824 VSS.n823 0.0228214
R473 VSS.n399 VSS.n398 0.0228214
R474 VSS.n712 VSS.n711 0.0228214
R475 VSS.n693 VSS.n692 0.0228214
R476 VSS.n580 VSS.n579 0.0228214
R477 VSS.n572 VSS.n571 0.0228214
R478 VSS.n553 VSS.n552 0.0228214
R479 VSS.n143 VSS.n142 0.0228214
R480 VSS.n194 VSS.n193 0.0228214
R481 VSS.n650 VSS.n649 0.0210357
R482 VSS.n380 VSS.n379 0.0210357
R483 VSS.n600 VSS.n599 0.0210357
R484 VSS.n96 VSS.n95 0.0210357
R485 VSS.n121 VSS.n118 0.0210357
R486 VSS.n26 VSS.n25 0.0210357
R487 VSS.n900 VSS.n899 0.0210357
R488 VSS.n944 VSS.n943 0.0210357
R489 VSS.n949 VSS.n948 0.0210357
R490 VSS.n118 VSS.n117 0.0201429
R491 VSS.n160 VSS.n159 0.0201429
R492 VSS.n25 VSS.n24 0.0201429
R493 VSS.n944 VSS.n921 0.0201429
R494 VSS.n213 VSS.n212 0.0201429
R495 VSS.n949 VSS.n882 0.0201429
R496 VSS.n76 VSS.n75 0.01925
R497 VSS.n252 VSS.n251 0.01925
R498 VSS.n802 VSS.n295 0.0174643
R499 VSS.n803 VSS.n802 0.0174643
R500 VSS.n798 VSS.n760 0.0174643
R501 VSS.n798 VSS.n797 0.0174643
R502 VSS.n714 VSS.n713 0.0174643
R503 VSS.n716 VSS.n715 0.0174643
R504 VSS.n578 VSS.n577 0.0174643
R505 VSS.n577 VSS.n573 0.0174643
R506 VSS.n22 VSS.n21 0.0174643
R507 VSS.n515 VSS.n463 0.0174643
R508 VSS.n515 VSS.n514 0.0174643
R509 VSS.n880 VSS.n879 0.0174643
R510 VSS.n302 VSS.n301 0.0165714
R511 VSS.n773 VSS.n772 0.0165714
R512 VSS.n767 VSS.n766 0.0165714
R513 VSS.n404 VSS.n400 0.0165714
R514 VSS.n323 VSS.n322 0.0165714
R515 VSS.n329 VSS.n328 0.0165714
R516 VSS.n330 VSS.n329 0.0165714
R517 VSS.n349 VSS.n348 0.0165714
R518 VSS.n725 VSS.n724 0.0165714
R519 VSS.n23 VSS.n22 0.0165714
R520 VSS.n28 VSS.n27 0.0165714
R521 VSS.n30 VSS.n29 0.0165714
R522 VSS.n437 VSS.n436 0.0165714
R523 VSS.n476 VSS.n475 0.0165714
R524 VSS.n470 VSS.n469 0.0165714
R525 VSS.n881 VSS.n880 0.0165714
R526 VSS.n947 VSS.n946 0.0165714
R527 VSS.n308 VSS.n307 0.0156786
R528 VSS.n731 VSS.n730 0.0156786
R529 VSS.n56 VSS.n55 0.0156786
R530 VSS.n11 VSS.n10 0.0156786
R531 VSS.n12 VSS.n11 0.0156786
R532 VSS.n1000 VSS.n40 0.0156786
R533 VSS.n1000 VSS.n999 0.0156786
R534 VSS.n443 VSS.n442 0.0156786
R535 VSS.n272 VSS.n271 0.0156786
R536 VSS.n867 VSS.n861 0.0156786
R537 VSS.n867 VSS.n866 0.0156786
R538 VSS.n962 VSS.n247 0.0156786
R539 VSS.n963 VSS.n962 0.0156786
R540 VSS.n456 VSS.n455 0.0152714
R541 VSS.n509 VSS.n508 0.0152714
R542 VSS.n492 VSS.n491 0.0152714
R543 VSS.n489 VSS.n488 0.0152714
R544 VSS.n341 VSS.n340 0.0152714
R545 VSS.n741 VSS.n740 0.0152714
R546 VSS.n753 VSS.n752 0.0152714
R547 VSS.n792 VSS.n791 0.0152714
R548 VSS.n874 VSS.n873 0.0152714
R549 VSS.n952 VSS.n951 0.0152714
R550 VSS.n19 VSS.n18 0.0147857
R551 VSS.n34 VSS.n33 0.0147857
R552 VSS.n877 VSS.n876 0.0147857
R553 VSS.n241 VSS.n240 0.0147857
R554 VSS.n169 VSS.n168 0.0138929
R555 VSS.n234 VSS.n233 0.0138929
R556 VSS.n499 VSS.n498 0.0132571
R557 VSS.n496 VSS.n495 0.0132571
R558 VSS.n485 VSS.n1 0.0132571
R559 VSS.n1003 VSS.n1002 0.0132571
R560 VSS.n782 VSS.n248 0.0132571
R561 VSS.n870 VSS.n869 0.0132571
R562 VSS.n956 VSS.n955 0.0132571
R563 VSS.n960 VSS.n959 0.0132571
R564 VSS.n833 VSS.n832 0.013
R565 VSS.n836 VSS.n835 0.013
R566 VSS.n766 VSS.n765 0.013
R567 VSS.n360 VSS.n359 0.013
R568 VSS.n363 VSS.n362 0.013
R569 VSS.n322 VSS.n321 0.013
R570 VSS.n533 VSS.n532 0.013
R571 VSS.n530 VSS.n529 0.013
R572 VSS.n469 VSS.n468 0.013
R573 VSS.n670 VSS.n669 0.0121071
R574 VSS.n667 VSS.n666 0.0121071
R575 VSS.n301 VSS.n300 0.0121071
R576 VSS.n769 VSS.n768 0.0121071
R577 VSS.n377 VSS.n376 0.0121071
R578 VSS.n684 VSS.n683 0.0121071
R579 VSS.n681 VSS.n680 0.0121071
R580 VSS.n325 VSS.n324 0.0121071
R581 VSS.n724 VSS.n723 0.0121071
R582 VSS.n619 VSS.n618 0.0121071
R583 VSS.n616 VSS.n615 0.0121071
R584 VSS.n55 VSS.n54 0.0121071
R585 VSS.n436 VSS.n435 0.0121071
R586 VSS.n472 VSS.n471 0.0121071
R587 VSS.n273 VSS.n272 0.0121071
R588 VSS.n666 VSS.n665 0.0112143
R589 VSS.n663 VSS.n652 0.0112143
R590 VSS.n827 VSS.n826 0.0112143
R591 VSS.n304 VSS.n303 0.0112143
R592 VSS.n685 VSS.n684 0.0112143
R593 VSS.n727 VSS.n726 0.0112143
R594 VSS.n615 VSS.n614 0.0112143
R595 VSS.n612 VSS.n602 0.0112143
R596 VSS.n550 VSS.n549 0.0112143
R597 VSS.n99 VSS.n98 0.0112143
R598 VSS.n140 VSS.n139 0.0112143
R599 VSS.n158 VSS.n157 0.0112143
R600 VSS.n170 VSS.n169 0.0112143
R601 VSS.n39 VSS.n38 0.0112143
R602 VSS.n439 VSS.n438 0.0112143
R603 VSS.n903 VSS.n902 0.0112143
R604 VSS.n923 VSS.n922 0.0112143
R605 VSS.n211 VSS.n210 0.0112143
R606 VSS.n235 VSS.n234 0.0112143
R607 VSS.n246 VSS.n245 0.0112143
R608 VSS.n664 VSS.n663 0.0103214
R609 VSS.n651 VSS.n650 0.0103214
R610 VSS.n632 VSS.n631 0.0103214
R611 VSS.n807 VSS.n806 0.0103214
R612 VSS.n832 VSS.n831 0.0103214
R613 VSS.n303 VSS.n302 0.0103214
R614 VSS.n313 VSS.n312 0.0103214
R615 VSS.n759 VSS.n758 0.0103214
R616 VSS.n778 VSS.n777 0.0103214
R617 VSS.n775 VSS.n774 0.0103214
R618 VSS.n364 VSS.n363 0.0103214
R619 VSS.n397 VSS.n396 0.0103214
R620 VSS.n710 VSS.n709 0.0103214
R621 VSS.n692 VSS.n691 0.0103214
R622 VSS.n690 VSS.n689 0.0103214
R623 VSS.n688 VSS.n687 0.0103214
R624 VSS.n333 VSS.n332 0.0103214
R625 VSS.n718 VSS.n717 0.0103214
R626 VSS.n736 VSS.n735 0.0103214
R627 VSS.n726 VSS.n725 0.0103214
R628 VSS.n613 VSS.n612 0.0103214
R629 VSS.n601 VSS.n600 0.0103214
R630 VSS.n582 VSS.n581 0.0103214
R631 VSS.n570 VSS.n569 0.0103214
R632 VSS.n534 VSS.n533 0.0103214
R633 VSS.n72 VSS.n59 0.0103214
R634 VSS.n75 VSS.n74 0.0103214
R635 VSS.n78 VSS.n77 0.0103214
R636 VSS.n9 VSS.n8 0.0103214
R637 VSS.n14 VSS.n13 0.0103214
R638 VSS.n438 VSS.n437 0.0103214
R639 VSS.n448 VSS.n447 0.0103214
R640 VSS.n462 VSS.n461 0.0103214
R641 VSS.n481 VSS.n480 0.0103214
R642 VSS.n478 VSS.n477 0.0103214
R643 VSS.n268 VSS.n267 0.0103214
R644 VSS.n253 VSS.n252 0.0103214
R645 VSS.n250 VSS.n249 0.0103214
R646 VSS.n860 VSS.n859 0.0103214
R647 VSS.n865 VSS.n864 0.0103214
R648 VSS.n491 VSS.n490 0.00956429
R649 VSS.n490 VSS.n489 0.00956429
R650 VSS.n950 VSS.n874 0.00956429
R651 VSS.n951 VSS.n950 0.00956429
R652 VSS.n668 VSS.n667 0.00942857
R653 VSS.n825 VSS.n824 0.00942857
R654 VSS.n829 VSS.n828 0.00942857
R655 VSS.n300 VSS.n299 0.00942857
R656 VSS.n310 VSS.n309 0.00942857
R657 VSS.n796 VSS.n795 0.00942857
R658 VSS.n768 VSS.n767 0.00942857
R659 VSS.n376 VSS.n365 0.00942857
R660 VSS.n379 VSS.n378 0.00942857
R661 VSS.n683 VSS.n682 0.00942857
R662 VSS.n324 VSS.n323 0.00942857
R663 VSS.n347 VSS.n346 0.00942857
R664 VSS.n733 VSS.n732 0.00942857
R665 VSS.n723 VSS.n722 0.00942857
R666 VSS.n617 VSS.n616 0.00942857
R667 VSS.n552 VSS.n551 0.00942857
R668 VSS.n548 VSS.n536 0.00942857
R669 VSS.n112 VSS.n111 0.00942857
R670 VSS.n117 VSS.n113 0.00942857
R671 VSS.n124 VSS.n123 0.00942857
R672 VSS.n161 VSS.n160 0.00942857
R673 VSS.n164 VSS.n163 0.00942857
R674 VSS.n998 VSS.n997 0.00942857
R675 VSS.n435 VSS.n434 0.00942857
R676 VSS.n445 VSS.n444 0.00942857
R677 VSS.n513 VSS.n512 0.00942857
R678 VSS.n471 VSS.n470 0.00942857
R679 VSS.n916 VSS.n915 0.00942857
R680 VSS.n921 VSS.n917 0.00942857
R681 VSS.n939 VSS.n938 0.00942857
R682 VSS.n214 VSS.n213 0.00942857
R683 VSS.n229 VSS.n228 0.00942857
R684 VSS.n965 VSS.n964 0.00942857
R685 VSS.n834 VSS.n833 0.00853571
R686 VSS.n765 VSS.n764 0.00853571
R687 VSS.n762 VSS.n761 0.00853571
R688 VSS.n362 VSS.n361 0.00853571
R689 VSS.n382 VSS.n381 0.00853571
R690 VSS.n318 VSS.n317 0.00853571
R691 VSS.n321 VSS.n320 0.00853571
R692 VSS.n332 VSS.n331 0.00853571
R693 VSS.n532 VSS.n531 0.00853571
R694 VSS.n95 VSS.n94 0.00853571
R695 VSS.n122 VSS.n121 0.00853571
R696 VSS.n154 VSS.n144 0.00853571
R697 VSS.n5 VSS.n4 0.00853571
R698 VSS.n18 VSS.n17 0.00853571
R699 VSS.n20 VSS.n19 0.00853571
R700 VSS.n35 VSS.n34 0.00853571
R701 VSS.n36 VSS.n35 0.00853571
R702 VSS.n994 VSS.n993 0.00853571
R703 VSS.n993 VSS.n992 0.00853571
R704 VSS.n991 VSS.n990 0.00853571
R705 VSS.n468 VSS.n467 0.00853571
R706 VSS.n465 VSS.n464 0.00853571
R707 VSS.n899 VSS.n898 0.00853571
R708 VSS.n943 VSS.n940 0.00853571
R709 VSS.n207 VSS.n195 0.00853571
R710 VSS.n853 VSS.n852 0.00853571
R711 VSS.n856 VSS.n855 0.00853571
R712 VSS.n876 VSS.n875 0.00853571
R713 VSS.n878 VSS.n877 0.00853571
R714 VSS.n242 VSS.n241 0.00853571
R715 VSS.n243 VSS.n242 0.00853571
R716 VSS.n969 VSS.n968 0.00853571
R717 VSS.n970 VSS.n969 0.00853571
R718 VSS.n972 VSS.n971 0.00853571
R719 VSS.n451 VSS.n450 0.00822143
R720 VSS.n455 VSS.n454 0.00822143
R721 VSS.n508 VSS.n507 0.00822143
R722 VSS.n504 VSS.n503 0.00822143
R723 VSS.n336 VSS.n335 0.00822143
R724 VSS.n340 VSS.n339 0.00822143
R725 VSS.n742 VSS.n741 0.00822143
R726 VSS.n746 VSS.n745 0.00822143
R727 VSS.n748 VSS.n747 0.00822143
R728 VSS.n752 VSS.n751 0.00822143
R729 VSS.n791 VSS.n790 0.00822143
R730 VSS.n787 VSS.n786 0.00822143
R731 VSS.n647 VSS.n646 0.00764286
R732 VSS.n822 VSS.n821 0.00764286
R733 VSS.n297 VSS.n296 0.00764286
R734 VSS.n309 VSS.n308 0.00764286
R735 VSS.n312 VSS.n311 0.00764286
R736 VSS.n758 VSS.n757 0.00764286
R737 VSS.n795 VSS.n794 0.00764286
R738 VSS.n777 VSS.n776 0.00764286
R739 VSS.n707 VSS.n695 0.00764286
R740 VSS.n346 VSS.n345 0.00764286
R741 VSS.n738 VSS.n718 0.00764286
R742 VSS.n734 VSS.n733 0.00764286
R743 VSS.n732 VSS.n731 0.00764286
R744 VSS.n720 VSS.n719 0.00764286
R745 VSS.n597 VSS.n596 0.00764286
R746 VSS.n555 VSS.n554 0.00764286
R747 VSS.n57 VSS.n56 0.00764286
R748 VSS.n59 VSS.n58 0.00764286
R749 VSS.n94 VSS.n93 0.00764286
R750 VSS.n144 VSS.n143 0.00764286
R751 VSS.n165 VSS.n164 0.00764286
R752 VSS.n166 VSS.n165 0.00764286
R753 VSS.n3 VSS.n2 0.00764286
R754 VSS.n4 VSS.n3 0.00764286
R755 VSS.n6 VSS.n5 0.00764286
R756 VSS.n8 VSS.n7 0.00764286
R757 VSS.n15 VSS.n14 0.00764286
R758 VSS.n17 VSS.n16 0.00764286
R759 VSS.n33 VSS.n32 0.00764286
R760 VSS.n38 VSS.n37 0.00764286
R761 VSS.n997 VSS.n996 0.00764286
R762 VSS.n996 VSS.n995 0.00764286
R763 VSS.n432 VSS.n431 0.00764286
R764 VSS.n444 VSS.n443 0.00764286
R765 VSS.n447 VSS.n446 0.00764286
R766 VSS.n461 VSS.n460 0.00764286
R767 VSS.n512 VSS.n511 0.00764286
R768 VSS.n480 VSS.n479 0.00764286
R769 VSS.n271 VSS.n270 0.00764286
R770 VSS.n269 VSS.n268 0.00764286
R771 VSS.n898 VSS.n897 0.00764286
R772 VSS.n195 VSS.n194 0.00764286
R773 VSS.n230 VSS.n229 0.00764286
R774 VSS.n231 VSS.n230 0.00764286
R775 VSS.n854 VSS.n853 0.00764286
R776 VSS.n855 VSS.n854 0.00764286
R777 VSS.n857 VSS.n856 0.00764286
R778 VSS.n859 VSS.n858 0.00764286
R779 VSS.n864 VSS.n863 0.00764286
R780 VSS.n240 VSS.n239 0.00764286
R781 VSS.n245 VSS.n244 0.00764286
R782 VSS.n966 VSS.n965 0.00764286
R783 VSS.n967 VSS.n966 0.00764286
R784 VSS.n646 VSS.n645 0.00675
R785 VSS.n631 VSS.n630 0.00675
R786 VSS.n821 VSS.n820 0.00675
R787 VSS.n311 VSS.n310 0.00675
R788 VSS.n314 VSS.n313 0.00675
R789 VSS.n794 VSS.n779 0.00675
R790 VSS.n776 VSS.n775 0.00675
R791 VSS.n774 VSS.n773 0.00675
R792 VSS.n365 VSS.n364 0.00675
R793 VSS.n396 VSS.n395 0.00675
R794 VSS.n711 VSS.n710 0.00675
R795 VSS.n695 VSS.n694 0.00675
R796 VSS.n345 VSS.n334 0.00675
R797 VSS.n737 VSS.n736 0.00675
R798 VSS.n735 VSS.n734 0.00675
R799 VSS.n596 VSS.n595 0.00675
R800 VSS.n581 VSS.n580 0.00675
R801 VSS.n567 VSS.n555 0.00675
R802 VSS.n58 VSS.n57 0.00675
R803 VSS.n93 VSS.n80 0.00675
R804 VSS.n98 VSS.n97 0.00675
R805 VSS.n111 VSS.n99 0.00675
R806 VSS.n141 VSS.n140 0.00675
R807 VSS.n167 VSS.n166 0.00675
R808 VSS.n7 VSS.n6 0.00675
R809 VSS.n16 VSS.n15 0.00675
R810 VSS.n21 VSS.n20 0.00675
R811 VSS.n31 VSS.n30 0.00675
R812 VSS.n995 VSS.n994 0.00675
R813 VSS.n992 VSS.n991 0.00675
R814 VSS.n446 VSS.n445 0.00675
R815 VSS.n449 VSS.n448 0.00675
R816 VSS.n511 VSS.n482 0.00675
R817 VSS.n479 VSS.n478 0.00675
R818 VSS.n477 VSS.n476 0.00675
R819 VSS.n270 VSS.n269 0.00675
R820 VSS.n897 VSS.n884 0.00675
R821 VSS.n902 VSS.n901 0.00675
R822 VSS.n915 VSS.n903 0.00675
R823 VSS.n232 VSS.n231 0.00675
R824 VSS.n858 VSS.n857 0.00675
R825 VSS.n863 VSS.n862 0.00675
R826 VSS.n879 VSS.n878 0.00675
R827 VSS.n238 VSS.n237 0.00675
R828 VSS.n968 VSS.n967 0.00675
R829 VSS.n971 VSS.n970 0.00675
R830 VSS.n52 VSS.n42 0.00636816
R831 VSS.n851 VSS.n850 0.00636816
R832 VSS.n989 VSS.n988 0.00636785
R833 VSS.n974 VSS.n973 0.00636785
R834 VSS.n498 VSS.n497 0.00620714
R835 VSS.n497 VSS.n496 0.00620714
R836 VSS.n1001 VSS.n1 0.00620714
R837 VSS.n1002 VSS.n1001 0.00620714
R838 VSS.n868 VSS.n248 0.00620714
R839 VSS.n869 VSS.n868 0.00620714
R840 VSS.n961 VSS.n956 0.00620714
R841 VSS.n961 VSS.n960 0.00620714
R842 VSS.n501 VSS.n500 0.00587143
R843 VSS.n494 VSS.n493 0.00587143
R844 VSS.n487 VSS.n486 0.00587143
R845 VSS.n1005 VSS.n1004 0.00587143
R846 VSS.n784 VSS.n783 0.00587143
R847 VSS.n872 VSS.n871 0.00587143
R848 VSS.n954 VSS.n953 0.00587143
R849 VSS.n958 VSS.n957 0.00587143
R850 VSS.n665 VSS.n664 0.00585714
R851 VSS.n633 VSS.n632 0.00585714
R852 VSS.n806 VSS.n805 0.00585714
R853 VSS.n808 VSS.n807 0.00585714
R854 VSS.n830 VSS.n829 0.00585714
R855 VSS.n307 VSS.n306 0.00585714
R856 VSS.n757 VSS.n314 0.00585714
R857 VSS.n779 VSS.n778 0.00585714
R858 VSS.n394 VSS.n382 0.00585714
R859 VSS.n398 VSS.n397 0.00585714
R860 VSS.n331 VSS.n330 0.00585714
R861 VSS.n334 VSS.n333 0.00585714
R862 VSS.n738 VSS.n737 0.00585714
R863 VSS.n730 VSS.n729 0.00585714
R864 VSS.n614 VSS.n613 0.00585714
R865 VSS.n583 VSS.n582 0.00585714
R866 VSS.n571 VSS.n570 0.00585714
R867 VSS.n569 VSS.n568 0.00585714
R868 VSS.n536 VSS.n535 0.00585714
R869 VSS.n79 VSS.n78 0.00585714
R870 VSS.n139 VSS.n138 0.00585714
R871 VSS.n155 VSS.n154 0.00585714
R872 VSS.n157 VSS.n156 0.00585714
R873 VSS.n37 VSS.n36 0.00585714
R874 VSS.n442 VSS.n441 0.00585714
R875 VSS.n460 VSS.n449 0.00585714
R876 VSS.n482 VSS.n481 0.00585714
R877 VSS.n937 VSS.n923 0.00585714
R878 VSS.n208 VSS.n207 0.00585714
R879 VSS.n210 VSS.n209 0.00585714
R880 VSS.n244 VSS.n243 0.00585714
R881 VSS.n680 VSS.n679 0.00565497
R882 VSS.n837 VSS.n836 0.00511752
R883 VSS.n529 VSS.n528 0.00511752
R884 VSS.n298 VSS.n297 0.00496429
R885 VSS.n306 VSS.n305 0.00496429
R886 VSS.n772 VSS.n771 0.00496429
R887 VSS.n771 VSS.n770 0.00496429
R888 VSS.n763 VSS.n762 0.00496429
R889 VSS.n709 VSS.n708 0.00496429
R890 VSS.n687 VSS.n686 0.00496429
R891 VSS.n319 VSS.n318 0.00496429
R892 VSS.n327 VSS.n326 0.00496429
R893 VSS.n328 VSS.n327 0.00496429
R894 VSS.n729 VSS.n728 0.00496429
R895 VSS.n721 VSS.n720 0.00496429
R896 VSS.n163 VSS.n162 0.00496429
R897 VSS.n24 VSS.n23 0.00496429
R898 VSS.n999 VSS.n998 0.00496429
R899 VSS.n433 VSS.n432 0.00496429
R900 VSS.n441 VSS.n440 0.00496429
R901 VSS.n475 VSS.n474 0.00496429
R902 VSS.n474 VSS.n473 0.00496429
R903 VSS.n466 VSS.n465 0.00496429
R904 VSS.n228 VSS.n215 0.00496429
R905 VSS.n882 VSS.n881 0.00496429
R906 VSS.n964 VSS.n963 0.00496429
R907 VSS.n459 VSS.n456 0.00486429
R908 VSS.n458 VSS.n457 0.00486429
R909 VSS.n484 VSS.n483 0.00486429
R910 VSS.n510 VSS.n509 0.00486429
R911 VSS.n344 VSS.n341 0.00486429
R912 VSS.n343 VSS.n342 0.00486429
R913 VSS.n316 VSS.n315 0.00486429
R914 VSS.n740 VSS.n739 0.00486429
R915 VSS.n756 VSS.n753 0.00486429
R916 VSS.n755 VSS.n754 0.00486429
R917 VSS.n781 VSS.n780 0.00486429
R918 VSS.n793 VSS.n792 0.00486429
R919 VSS.n1007 VSS 0.00452857
R920 VSS.n1008 VSS 0.00452857
R921 VSS.n381 VSS.n380 0.00407143
R922 VSS.n54 VSS.n53 0.00407143
R923 VSS.n73 VSS.n72 0.00407143
R924 VSS.n77 VSS.n76 0.00407143
R925 VSS.n171 VSS.n170 0.00407143
R926 VSS.n10 VSS.n9 0.00407143
R927 VSS.n13 VSS.n12 0.00407143
R928 VSS.n27 VSS.n26 0.00407143
R929 VSS.n274 VSS.n273 0.00407143
R930 VSS.n267 VSS.n254 0.00407143
R931 VSS.n251 VSS.n250 0.00407143
R932 VSS.n236 VSS.n235 0.00407143
R933 VSS.n861 VSS.n860 0.00407143
R934 VSS.n866 VSS.n865 0.00407143
R935 VSS.n948 VSS.n947 0.00407143
R936 VSS.n502 VSS.n501 0.00352143
R937 VSS.n500 VSS.n499 0.00352143
R938 VSS.n495 VSS.n494 0.00352143
R939 VSS.n493 VSS.n492 0.00352143
R940 VSS.n488 VSS.n487 0.00352143
R941 VSS.n486 VSS.n485 0.00352143
R942 VSS.n1004 VSS.n1003 0.00352143
R943 VSS.n1006 VSS.n1005 0.00352143
R944 VSS.n785 VSS.n784 0.00352143
R945 VSS.n783 VSS.n782 0.00352143
R946 VSS.n871 VSS.n870 0.00352143
R947 VSS.n873 VSS.n872 0.00352143
R948 VSS.n953 VSS.n952 0.00352143
R949 VSS.n955 VSS.n954 0.00352143
R950 VSS.n959 VSS.n958 0.00352143
R951 VSS.n957 VSS.n0 0.00352143
R952 VSS.n459 VSS.n458 0.00318571
R953 VSS.n510 VSS.n484 0.00318571
R954 VSS.n344 VSS.n343 0.00318571
R955 VSS.n739 VSS.n316 0.00318571
R956 VSS.n756 VSS.n755 0.00318571
R957 VSS.n793 VSS.n781 0.00318571
R958 VSS.n669 VSS.n668 0.00317857
R959 VSS.n652 VSS.n651 0.00317857
R960 VSS.n804 VSS.n803 0.00317857
R961 VSS.n823 VSS.n822 0.00317857
R962 VSS.n826 VSS.n825 0.00317857
R963 VSS.n835 VSS.n834 0.00317857
R964 VSS.n299 VSS.n298 0.00317857
R965 VSS.n305 VSS.n304 0.00317857
R966 VSS.n797 VSS.n796 0.00317857
R967 VSS.n770 VSS.n769 0.00317857
R968 VSS.n764 VSS.n763 0.00317857
R969 VSS.n361 VSS.n360 0.00317857
R970 VSS.n378 VSS.n377 0.00317857
R971 VSS.n400 VSS.n399 0.00317857
R972 VSS.n694 VSS.n693 0.00317857
R973 VSS.n691 VSS.n690 0.00317857
R974 VSS.n682 VSS.n681 0.00317857
R975 VSS.n320 VSS.n319 0.00317857
R976 VSS.n326 VSS.n325 0.00317857
R977 VSS.n348 VSS.n347 0.00317857
R978 VSS.n728 VSS.n727 0.00317857
R979 VSS.n722 VSS.n721 0.00317857
R980 VSS.n618 VSS.n617 0.00317857
R981 VSS.n602 VSS.n601 0.00317857
R982 VSS.n573 VSS.n572 0.00317857
R983 VSS.n554 VSS.n553 0.00317857
R984 VSS.n551 VSS.n550 0.00317857
R985 VSS.n531 VSS.n530 0.00317857
R986 VSS.n53 VSS.n52 0.00317857
R987 VSS.n113 VSS.n112 0.00317857
R988 VSS.n123 VSS.n122 0.00317857
R989 VSS.n159 VSS.n158 0.00317857
R990 VSS.n168 VSS.n167 0.00317857
R991 VSS.n988 VSS.n171 0.00317857
R992 VSS.n40 VSS.n39 0.00317857
R993 VSS.n434 VSS.n433 0.00317857
R994 VSS.n440 VSS.n439 0.00317857
R995 VSS.n514 VSS.n513 0.00317857
R996 VSS.n473 VSS.n472 0.00317857
R997 VSS.n467 VSS.n466 0.00317857
R998 VSS.n850 VSS.n274 0.00317857
R999 VSS.n917 VSS.n916 0.00317857
R1000 VSS.n940 VSS.n939 0.00317857
R1001 VSS.n212 VSS.n211 0.00317857
R1002 VSS.n233 VSS.n232 0.00317857
R1003 VSS.n974 VSS.n236 0.00317857
R1004 VSS.n247 VSS.n246 0.00317857
R1005 VSS.n649 VSS.n648 0.00228571
R1006 VSS.n648 VSS.n647 0.00228571
R1007 VSS.n645 VSS.n633 0.00228571
R1008 VSS.n629 VSS.n295 0.00228571
R1009 VSS.n820 VSS.n808 0.00228571
R1010 VSS.n760 VSS.n759 0.00228571
R1011 VSS.n395 VSS.n394 0.00228571
R1012 VSS.n713 VSS.n712 0.00228571
R1013 VSS.n708 VSS.n707 0.00228571
R1014 VSS.n717 VSS.n716 0.00228571
R1015 VSS.n599 VSS.n598 0.00228571
R1016 VSS.n598 VSS.n597 0.00228571
R1017 VSS.n595 VSS.n583 0.00228571
R1018 VSS.n579 VSS.n578 0.00228571
R1019 VSS.n568 VSS.n567 0.00228571
R1020 VSS.n74 VSS.n73 0.00228571
R1021 VSS.n80 VSS.n79 0.00228571
R1022 VSS.n97 VSS.n96 0.00228571
R1023 VSS.n156 VSS.n155 0.00228571
R1024 VSS.n162 VSS.n161 0.00228571
R1025 VSS.n463 VSS.n462 0.00228571
R1026 VSS.n254 VSS.n253 0.00228571
R1027 VSS.n884 VSS.n883 0.00228571
R1028 VSS.n901 VSS.n900 0.00228571
R1029 VSS.n209 VSS.n208 0.00228571
R1030 VSS.n215 VSS.n214 0.00228571
R1031 VSS.n452 VSS.n451 0.00217857
R1032 VSS.n454 VSS.n453 0.00217857
R1033 VSS.n507 VSS.n506 0.00217857
R1034 VSS.n505 VSS.n504 0.00217857
R1035 VSS.n337 VSS.n336 0.00217857
R1036 VSS.n339 VSS.n338 0.00217857
R1037 VSS.n743 VSS.n742 0.00217857
R1038 VSS.n745 VSS.n744 0.00217857
R1039 VSS.n749 VSS.n748 0.00217857
R1040 VSS.n751 VSS.n750 0.00217857
R1041 VSS.n790 VSS.n789 0.00217857
R1042 VSS.n788 VSS.n787 0.00217857
R1043 VSS.n828 VSS.n827 0.00139286
R1044 VSS.n831 VSS.n830 0.00139286
R1045 VSS.n714 VSS.n404 0.00139286
R1046 VSS.n689 VSS.n688 0.00139286
R1047 VSS.n686 VSS.n685 0.00139286
R1048 VSS.n715 VSS.n349 0.00139286
R1049 VSS.n549 VSS.n548 0.00139286
R1050 VSS.n535 VSS.n534 0.00139286
R1051 VSS.n138 VSS.n124 0.00139286
R1052 VSS.n142 VSS.n141 0.00139286
R1053 VSS.n29 VSS.n28 0.00139286
R1054 VSS.n32 VSS.n31 0.00139286
R1055 VSS.n938 VSS.n937 0.00139286
R1056 VSS.n193 VSS.n192 0.00139286
R1057 VSS.n946 VSS.n945 0.00139286
R1058 VSS.n239 VSS.n238 0.00139286
R1059 D0 D0.n0 115.853
R1060 D0.n0 D0.t1 81.9405
R1061 D0.n0 D0.t0 56.8765
R1062 VCC.n498 VCC.t15 4282.54
R1063 VCC.n672 VCC.t30 4282.54
R1064 VCC.t10 VCC.t24 1149.1
R1065 VCC.t23 VCC.t31 1149.1
R1066 VCC.t15 VCC.t10 978.443
R1067 VCC.t30 VCC.t23 978.443
R1068 VCC.t24 VCC.t9 972.755
R1069 VCC.t31 VCC.t22 972.755
R1070 VCC.t9 VCC.n497 723.087
R1071 VCC.t22 VCC.n671 723.087
R1072 VCC.t5 VCC.t2 571.485
R1073 VCC.t19 VCC.t18 571.485
R1074 VCC.t6 VCC.t29 571.485
R1075 VCC.n381 VCC.t19 544.823
R1076 VCC.n21 VCC.t6 544.823
R1077 VCC.n775 VCC.t5 542.996
R1078 VCC.n382 VCC.n381 187.349
R1079 VCC.n498 VCC.n338 187.349
R1080 VCC.n22 VCC.n21 187.349
R1081 VCC.n673 VCC.n672 187.349
R1082 VCC.n431 VCC.n430 185
R1083 VCC.n432 VCC.n431 185
R1084 VCC.n351 VCC.n350 185
R1085 VCC.n467 VCC.n351 185
R1086 VCC.n488 VCC.n487 185
R1087 VCC.n489 VCC.n488 185
R1088 VCC.n486 VCC.n339 185
R1089 VCC.n490 VCC.n339 185
R1090 VCC.n470 VCC.n469 185
R1091 VCC.n469 VCC.n468 185
R1092 VCC.n499 VCC.n340 185
R1093 VCC.n380 VCC.n379 185
R1094 VCC.n378 VCC.n377 185
R1095 VCC.n408 VCC.n378 185
R1096 VCC.n411 VCC.n410 185
R1097 VCC.n410 VCC.n409 185
R1098 VCC.n366 VCC.n365 185
R1099 VCC.n433 VCC.n366 185
R1100 VCC.n493 VCC.n315 185
R1101 VCC.n491 VCC.n315 185
R1102 VCC.n314 VCC.n313 185
R1103 VCC.n543 VCC.n314 185
R1104 VCC.n564 VCC.n563 185
R1105 VCC.n564 VCC.n300 185
R1106 VCC.n283 VCC.n282 185
R1107 VCC.n282 VCC.n281 185
R1108 VCC.n601 VCC.n600 185
R1109 VCC.n600 VCC.n599 185
R1110 VCC.n620 VCC.n619 185
R1111 VCC.n621 VCC.n620 185
R1112 VCC.n570 VCC.n569 185
R1113 VCC.n569 VCC.n568 185
R1114 VCC.n547 VCC.n546 185
R1115 VCC.n546 VCC.n545 185
R1116 VCC.n565 VCC.n298 185
R1117 VCC.n566 VCC.n565 185
R1118 VCC.n280 VCC.n279 185
R1119 VCC.n598 VCC.n280 185
R1120 VCC.n265 VCC.n264 185
R1121 VCC.n495 VCC.n494 185
R1122 VCC.n495 VCC.n492 185
R1123 VCC.n39 VCC.n12 185
R1124 VCC.n720 VCC.n12 185
R1125 VCC.n99 VCC.n98 185
R1126 VCC.n100 VCC.n99 185
R1127 VCC.n77 VCC.n75 185
R1128 VCC.n685 VCC.n77 185
R1129 VCC.n683 VCC.n682 185
R1130 VCC.n684 VCC.n683 185
R1131 VCC.n97 VCC.n76 185
R1132 VCC.n101 VCC.n76 185
R1133 VCC.n111 VCC.n109 185
R1134 VCC.n20 VCC.n18 185
R1135 VCC.n34 VCC.n33 185
R1136 VCC.n35 VCC.n34 185
R1137 VCC.n11 VCC.n9 185
R1138 VCC.n36 VCC.n11 185
R1139 VCC.n718 VCC.n717 185
R1140 VCC.n719 VCC.n718 185
R1141 VCC.n257 VCC.n256 185
R1142 VCC.n258 VCC.n257 185
R1143 VCC.n192 VCC.n191 185
R1144 VCC.n191 VCC.n190 185
R1145 VCC.n223 VCC.n222 185
R1146 VCC.n224 VCC.n223 185
R1147 VCC.n178 VCC.n177 185
R1148 VCC.n242 VCC.n178 185
R1149 VCC.n245 VCC.n244 185
R1150 VCC.n244 VCC.n243 185
R1151 VCC.n229 VCC.n180 185
R1152 VCC.n180 VCC.n179 185
R1153 VCC.n228 VCC.n227 185
R1154 VCC.n227 VCC.n226 185
R1155 VCC.n221 VCC.n184 185
R1156 VCC.n184 VCC.n183 185
R1157 VCC.n213 VCC.n187 185
R1158 VCC.n217 VCC.n187 185
R1159 VCC.n215 VCC.n214 185
R1160 VCC.n216 VCC.n215 185
R1161 VCC.n114 VCC.n113 185
R1162 VCC.n113 VCC.n112 185
R1163 VCC.n168 VCC.n167 185
R1164 VCC.n432 VCC.n367 96.8274
R1165 VCC.n468 VCC.n341 96.8274
R1166 VCC.n721 VCC.n720 96.8274
R1167 VCC.n686 VCC.n101 96.8274
R1168 VCC.n879 VCC.n876 95.0005
R1169 VCC.n434 VCC.n352 95.0005
R1170 VCC.n466 VCC.n352 95.0005
R1171 VCC.n85 VCC.n37 95.0005
R1172 VCC.n85 VCC.n78 95.0005
R1173 VCC.n545 VCC.n544 93.2412
R1174 VCC.n567 VCC.n566 93.2412
R1175 VCC.n568 VCC.n567 93.2412
R1176 VCC.n621 VCC.n266 93.2412
R1177 VCC.n218 VCC.n217 93.2412
R1178 VCC.n225 VCC.n224 93.2412
R1179 VCC.n226 VCC.n225 93.2412
R1180 VCC.n258 VCC.n169 93.2412
R1181 VCC.n405 VCC.n382 92.5398
R1182 VCC.n502 VCC.n338 92.5398
R1183 VCC.n23 VCC.n22 92.5398
R1184 VCC.n674 VCC.n673 92.5398
R1185 VCC.n457 VCC.n353 92.5005
R1186 VCC.n353 VCC.n352 92.5005
R1187 VCC.n87 VCC.n86 92.5005
R1188 VCC.n86 VCC.n85 92.5005
R1189 VCC.t16 VCC.n407 73.0774
R1190 VCC.n19 VCC.t27 73.0774
R1191 VCC.n838 VCC.t25 72.544
R1192 VCC.t32 VCC.n597 70.3709
R1193 VCC.t13 VCC.n241 70.3709
R1194 VCC.n542 VCC.t11 66.8524
R1195 VCC.t20 VCC.n188 66.8524
R1196 VCC.n500 VCC.t7 65.7697
R1197 VCC.n110 VCC.t0 65.7697
R1198 VCC.n406 VCC.n378 50.3505
R1199 VCC.n431 VCC.n368 50.3505
R1200 VCC.n469 VCC.n342 50.3505
R1201 VCC.n501 VCC.n339 50.3505
R1202 VCC.n34 VCC.n13 50.3505
R1203 VCC.n722 VCC.n12 50.3505
R1204 VCC.n687 VCC.n76 50.3505
R1205 VCC.n683 VCC.n102 50.3505
R1206 VCC.n880 VCC.n873 49.4005
R1207 VCC.n435 VCC.n353 49.4005
R1208 VCC.n465 VCC.n353 49.4005
R1209 VCC.n86 VCC.n38 49.4005
R1210 VCC.n86 VCC.n79 49.4005
R1211 VCC.n541 VCC.n315 43.1576
R1212 VCC.n546 VCC.n301 43.1576
R1213 VCC.n565 VCC.n299 43.1576
R1214 VCC.n569 VCC.n299 43.1576
R1215 VCC.n596 VCC.n280 43.1576
R1216 VCC.n620 VCC.n267 43.1576
R1217 VCC.n191 VCC.n189 43.1576
R1218 VCC.n219 VCC.n187 43.1576
R1219 VCC.n223 VCC.n182 43.1576
R1220 VCC.n227 VCC.n182 43.1576
R1221 VCC.n240 VCC.n178 43.1576
R1222 VCC.n257 VCC.n170 43.1576
R1223 VCC.n622 VCC.n621 36.8662
R1224 VCC.n259 VCC.n258 36.8662
R1225 VCC.n518 VCC.t8 35.5869
R1226 VCC.n129 VCC.t1 35.5869
R1227 VCC.n611 VCC.t33 34.994
R1228 VCC.n173 VCC.t14 34.994
R1229 VCC.n311 VCC.t12 34.9892
R1230 VCC.n138 VCC.t21 34.9892
R1231 VCC.n832 VCC.t26 34.9619
R1232 VCC.n371 VCC.t17 34.945
R1233 VCC.n54 VCC.t28 34.945
R1234 VCC.n808 VCC.t4 34.9423
R1235 VCC.t7 VCC.n490 31.0582
R1236 VCC.n684 VCC.t0 31.0582
R1237 VCC.n818 VCC.n817 29.2313
R1238 VCC.n879 VCC.n878 29.2313
R1239 VCC.n434 VCC.n433 29.2313
R1240 VCC.n467 VCC.n466 29.2313
R1241 VCC.n719 VCC.n37 29.2313
R1242 VCC.n100 VCC.n78 29.2313
R1243 VCC.n491 VCC.t11 26.3894
R1244 VCC.n566 VCC.n300 26.3894
R1245 VCC.n568 VCC.n281 26.3894
R1246 VCC.n190 VCC.t20 26.3894
R1247 VCC.n224 VCC.n183 26.3894
R1248 VCC.n226 VCC.n179 26.3894
R1249 VCC.n798 VCC.n797 25.5774
R1250 VCC.n858 VCC.n857 25.5774
R1251 VCC.n409 VCC.n367 25.5774
R1252 VCC.n489 VCC.n341 25.5774
R1253 VCC.n721 VCC.n36 25.5774
R1254 VCC.n686 VCC.n685 25.5774
R1255 VCC.n408 VCC.t16 23.7505
R1256 VCC.n35 VCC.t27 23.7505
R1257 VCC.n545 VCC.n543 22.8709
R1258 VCC.n598 VCC.t32 22.8709
R1259 VCC.n599 VCC.n598 22.8709
R1260 VCC.n217 VCC.n216 22.8709
R1261 VCC.n242 VCC.t13 22.8709
R1262 VCC.n243 VCC.n242 22.8709
R1263 VCC.n777 VCC.n776 21.9236
R1264 VCC.n796 VCC.t3 21.9236
R1265 VCC.n407 VCC.n379 21.9236
R1266 VCC.n500 VCC.n499 21.9236
R1267 VCC.n20 VCC.n19 21.9236
R1268 VCC.n111 VCC.n110 21.9236
R1269 VCC.n492 VCC.n491 19.3524
R1270 VCC.n190 VCC.n112 19.3524
R1271 VCC.n819 VCC.n815 15.2005
R1272 VCC.n880 VCC.n875 15.2005
R1273 VCC.n435 VCC.n366 15.2005
R1274 VCC.n465 VCC.n351 15.2005
R1275 VCC.n718 VCC.n38 15.2005
R1276 VCC.n99 VCC.n79 15.2005
R1277 VCC.n799 VCC.n795 13.3005
R1278 VCC.n859 VCC.n855 13.3005
R1279 VCC.n410 VCC.n368 13.3005
R1280 VCC.n488 VCC.n342 13.3005
R1281 VCC.n722 VCC.n11 13.3005
R1282 VCC.n687 VCC.n77 13.3005
R1283 VCC.n565 VCC.n564 12.2148
R1284 VCC.n569 VCC.n282 12.2148
R1285 VCC.n223 VCC.n184 12.2148
R1286 VCC.n227 VCC.n180 12.2148
R1287 VCC.n778 VCC.n774 11.4005
R1288 VCC.n406 VCC.n380 11.4005
R1289 VCC.n501 VCC.n340 11.4005
R1290 VCC.n18 VCC.n13 11.4005
R1291 VCC.n109 VCC.n102 11.4005
R1292 VCC.n546 VCC.n314 10.5862
R1293 VCC.n600 VCC.n280 10.5862
R1294 VCC.n215 VCC.n187 10.5862
R1295 VCC.n244 VCC.n178 10.5862
R1296 VCC.n497 VCC.n492 10.5561
R1297 VCC.n671 VCC.n112 10.5561
R1298 VCC.n623 VCC.n622 9.80483
R1299 VCC.n260 VCC.n259 9.80483
R1300 VCC.n496 VCC.n324 9.38146
R1301 VCC.n670 VCC.n669 9.38146
R1302 VCC.n881 VCC.n880 9.3005
R1303 VCC.n880 VCC.n879 9.3005
R1304 VCC.n860 VCC.n859 9.3005
R1305 VCC.n859 VCC.n858 9.3005
R1306 VCC.n779 VCC.n778 9.3005
R1307 VCC.n778 VCC.n777 9.3005
R1308 VCC.n800 VCC.n799 9.3005
R1309 VCC.n799 VCC.n798 9.3005
R1310 VCC.n820 VCC.n819 9.3005
R1311 VCC.n819 VCC.n818 9.3005
R1312 VCC.n429 VCC.n428 9.3005
R1313 VCC.n399 VCC.n398 9.3005
R1314 VCC.n505 VCC.n504 9.3005
R1315 VCC.n472 VCC.n471 9.3005
R1316 VCC.n461 VCC.n354 9.3005
R1317 VCC.n460 VCC.n459 9.3005
R1318 VCC.n344 VCC.n343 9.3005
R1319 VCC.n337 VCC.n335 9.3005
R1320 VCC.n370 VCC.n369 9.3005
R1321 VCC.n397 VCC.n392 9.3005
R1322 VCC.n437 VCC.n364 9.3005
R1323 VCC.n357 VCC.n356 9.3005
R1324 VCC.n464 VCC.n349 9.3005
R1325 VCC.n465 VCC.n464 9.3005
R1326 VCC.n466 VCC.n465 9.3005
R1327 VCC.n485 VCC.n332 9.3005
R1328 VCC.n485 VCC.n342 9.3005
R1329 VCC.n342 VCC.n341 9.3005
R1330 VCC.n502 VCC.n327 9.3005
R1331 VCC.n502 VCC.n501 9.3005
R1332 VCC.n501 VCC.n500 9.3005
R1333 VCC.n405 VCC.n404 9.3005
R1334 VCC.n406 VCC.n405 9.3005
R1335 VCC.n407 VCC.n406 9.3005
R1336 VCC.n414 VCC.n413 9.3005
R1337 VCC.n413 VCC.n368 9.3005
R1338 VCC.n368 VCC.n367 9.3005
R1339 VCC.n436 VCC.n363 9.3005
R1340 VCC.n436 VCC.n435 9.3005
R1341 VCC.n435 VCC.n434 9.3005
R1342 VCC.n595 VCC.n594 9.3005
R1343 VCC.n596 VCC.n595 9.3005
R1344 VCC.n597 VCC.n596 9.3005
R1345 VCC.n541 VCC.n540 9.3005
R1346 VCC.n542 VCC.n541 9.3005
R1347 VCC.n549 VCC.n548 9.3005
R1348 VCC.n562 VCC.n561 9.3005
R1349 VCC.n562 VCC.n301 9.3005
R1350 VCC.n544 VCC.n301 9.3005
R1351 VCC.n588 VCC.n587 9.3005
R1352 VCC.n604 VCC.n603 9.3005
R1353 VCC.n603 VCC.n267 9.3005
R1354 VCC.n267 VCC.n266 9.3005
R1355 VCC.n269 VCC.n268 9.3005
R1356 VCC.n618 VCC.n617 9.3005
R1357 VCC.n497 VCC.n496 9.3005
R1358 VCC.n50 VCC.n49 9.3005
R1359 VCC.n32 VCC.n31 9.3005
R1360 VCC.n105 VCC.n103 9.3005
R1361 VCC.n96 VCC.n95 9.3005
R1362 VCC.n91 VCC.n80 9.3005
R1363 VCC.n90 VCC.n89 9.3005
R1364 VCC.n74 VCC.n72 9.3005
R1365 VCC.n681 VCC.n680 9.3005
R1366 VCC.n48 VCC.n47 9.3005
R1367 VCC.n17 VCC.n14 9.3005
R1368 VCC.n81 VCC.n42 9.3005
R1369 VCC.n83 VCC.n82 9.3005
R1370 VCC.n94 VCC.n69 9.3005
R1371 VCC.n94 VCC.n79 9.3005
R1372 VCC.n79 VCC.n78 9.3005
R1373 VCC.n688 VCC.n73 9.3005
R1374 VCC.n688 VCC.n687 9.3005
R1375 VCC.n687 VCC.n686 9.3005
R1376 VCC.n674 VCC.n108 9.3005
R1377 VCC.n674 VCC.n102 9.3005
R1378 VCC.n110 VCC.n102 9.3005
R1379 VCC.n23 VCC.n2 9.3005
R1380 VCC.n23 VCC.n13 9.3005
R1381 VCC.n19 VCC.n13 9.3005
R1382 VCC.n724 VCC.n723 9.3005
R1383 VCC.n723 VCC.n722 9.3005
R1384 VCC.n722 VCC.n721 9.3005
R1385 VCC.n716 VCC.n715 9.3005
R1386 VCC.n716 VCC.n38 9.3005
R1387 VCC.n38 VCC.n37 9.3005
R1388 VCC.n212 VCC.n211 9.3005
R1389 VCC.n239 VCC.n238 9.3005
R1390 VCC.n240 VCC.n239 9.3005
R1391 VCC.n241 VCC.n240 9.3005
R1392 VCC.n172 VCC.n171 9.3005
R1393 VCC.n233 VCC.n232 9.3005
R1394 VCC.n255 VCC.n254 9.3005
R1395 VCC.n246 VCC.n176 9.3005
R1396 VCC.n246 VCC.n170 9.3005
R1397 VCC.n170 VCC.n169 9.3005
R1398 VCC.n220 VCC.n186 9.3005
R1399 VCC.n220 VCC.n219 9.3005
R1400 VCC.n219 VCC.n218 9.3005
R1401 VCC.n205 VCC.n189 9.3005
R1402 VCC.n189 VCC.n188 9.3005
R1403 VCC.n671 VCC.n670 9.3005
R1404 VCC.n776 VCC.n775 9.13511
R1405 VCC.n381 VCC.n379 9.13511
R1406 VCC.n499 VCC.n498 9.13511
R1407 VCC.n21 VCC.n20 9.13511
R1408 VCC.n672 VCC.n111 9.13511
R1409 VCC.n495 VCC.n315 8.95764
R1410 VCC.n620 VCC.n265 8.95764
R1411 VCC.n191 VCC.n113 8.95764
R1412 VCC.n257 VCC.n168 8.95764
R1413 VCC.n571 VCC.n299 8.85536
R1414 VCC.n567 VCC.n299 8.85536
R1415 VCC.n182 VCC.n181 8.85536
R1416 VCC.n225 VCC.n182 8.85536
R1417 VCC.n839 VCC.n838 8.47776
R1418 VCC.n543 VCC.n542 7.03754
R1419 VCC.n599 VCC.n266 7.03754
R1420 VCC.n216 VCC.n188 7.03754
R1421 VCC.n243 VCC.n169 7.03754
R1422 VCC.n797 VCC.n796 5.48127
R1423 VCC.n857 VCC.n856 5.48127
R1424 VCC.n409 VCC.n408 5.48127
R1425 VCC.n490 VCC.n489 5.48127
R1426 VCC.n36 VCC.n35 5.48127
R1427 VCC.n685 VCC.n684 5.48127
R1428 VCC.n496 VCC.n495 4.88621
R1429 VCC.n670 VCC.n113 4.88621
R1430 VCC.n571 VCC.n298 4.84621
R1431 VCC.n571 VCC.n570 4.84621
R1432 VCC.n222 VCC.n181 4.84621
R1433 VCC.n228 VCC.n181 4.84621
R1434 VCC.n524 VCC.n316 4.6505
R1435 VCC.n199 VCC.n193 4.6505
R1436 VCC.n386 VCC.n384 4.51121
R1437 VCC.n731 VCC.n730 4.51121
R1438 VCC.n823 VCC.n822 4.5005
R1439 VCC.n804 VCC.n803 4.5005
R1440 VCC.n783 VCC.n782 4.5005
R1441 VCC.n829 VCC.n828 4.5005
R1442 VCC.n888 VCC.n887 4.5005
R1443 VCC.n883 VCC.n882 4.5005
R1444 VCC.n862 VCC.n861 4.5005
R1445 VCC.n841 VCC.n840 4.5005
R1446 VCC.n508 VCC.n333 4.5005
R1447 VCC.n507 VCC.n506 4.5005
R1448 VCC.n401 VCC.n400 4.5005
R1449 VCC.n396 VCC.n393 4.5005
R1450 VCC.n425 VCC.n424 4.5005
R1451 VCC.n395 VCC.n394 4.5005
R1452 VCC.n519 VCC.n518 4.5005
R1453 VCC.n475 VCC.n474 4.5005
R1454 VCC.n473 VCC.n345 4.5005
R1455 VCC.n510 VCC.n509 4.5005
R1456 VCC.n427 VCC.n426 4.5005
R1457 VCC.n440 VCC.n439 4.5005
R1458 VCC.n439 VCC.n438 4.5005
R1459 VCC.n376 VCC.n372 4.5005
R1460 VCC.n412 VCC.n376 4.5005
R1461 VCC.n403 VCC.n402 4.5005
R1462 VCC.n403 VCC.n383 4.5005
R1463 VCC.n455 VCC.n454 4.5005
R1464 VCC.n456 VCC.n455 4.5005
R1465 VCC.n447 VCC.n355 4.5005
R1466 VCC.n458 VCC.n355 4.5005
R1467 VCC.n462 VCC.n347 4.5005
R1468 VCC.n463 VCC.n462 4.5005
R1469 VCC.n483 VCC.n482 4.5005
R1470 VCC.n484 VCC.n483 4.5005
R1471 VCC.n336 VCC.n334 4.5005
R1472 VCC.n503 VCC.n336 4.5005
R1473 VCC.n276 VCC.n271 4.5005
R1474 VCC.n616 VCC.n615 4.5005
R1475 VCC.n526 VCC.n525 4.5005
R1476 VCC.n319 VCC.n317 4.5005
R1477 VCC.n551 VCC.n550 4.5005
R1478 VCC.n305 VCC.n303 4.5005
R1479 VCC.n303 VCC.n302 4.5005
R1480 VCC.n307 VCC.n306 4.5005
R1481 VCC.n534 VCC.n309 4.5005
R1482 VCC.n539 VCC.n538 4.5005
R1483 VCC.n523 VCC.n522 4.5005
R1484 VCC.n528 VCC.n527 4.5005
R1485 VCC.n278 VCC.n277 4.5005
R1486 VCC.n602 VCC.n278 4.5005
R1487 VCC.n590 VCC.n589 4.5005
R1488 VCC.n288 VCC.n275 4.5005
R1489 VCC.n580 VCC.n579 4.5005
R1490 VCC.n297 VCC.n295 4.5005
R1491 VCC.n581 VCC.n290 4.5005
R1492 VCC.n591 VCC.n286 4.5005
R1493 VCC.n593 VCC.n592 4.5005
R1494 VCC.n593 VCC.n284 4.5005
R1495 VCC.n614 VCC.n270 4.5005
R1496 VCC.n625 VCC.n624 4.5005
R1497 VCC.n312 VCC.n310 4.5005
R1498 VCC.n106 VCC.n104 4.5005
R1499 VCC.n679 VCC.n678 4.5005
R1500 VCC.n27 VCC.n15 4.5005
R1501 VCC.n30 VCC.n29 4.5005
R1502 VCC.n53 VCC.n46 4.5005
R1503 VCC.n28 VCC.n16 4.5005
R1504 VCC.n130 VCC.n129 4.5005
R1505 VCC.n695 VCC.n694 4.5005
R1506 VCC.n693 VCC.n70 4.5005
R1507 VCC.n121 VCC.n120 4.5005
R1508 VCC.n56 VCC.n55 4.5005
R1509 VCC.n714 VCC.n713 4.5005
R1510 VCC.n714 VCC.n40 4.5005
R1511 VCC.n45 VCC.n8 4.5005
R1512 VCC.n10 VCC.n8 4.5005
R1513 VCC.n26 VCC.n25 4.5005
R1514 VCC.n25 VCC.n24 4.5005
R1515 VCC.n63 VCC.n61 4.5005
R1516 VCC.n84 VCC.n63 4.5005
R1517 VCC.n703 VCC.n64 4.5005
R1518 VCC.n88 VCC.n64 4.5005
R1519 VCC.n92 VCC.n67 4.5005
R1520 VCC.n93 VCC.n92 4.5005
R1521 VCC.n691 VCC.n690 4.5005
R1522 VCC.n690 VCC.n689 4.5005
R1523 VCC.n677 VCC.n676 4.5005
R1524 VCC.n676 VCC.n675 4.5005
R1525 VCC.n251 VCC.n174 4.5005
R1526 VCC.n253 VCC.n252 4.5005
R1527 VCC.n235 VCC.n234 4.5005
R1528 VCC.n210 VCC.n209 4.5005
R1529 VCC.n202 VCC.n194 4.5005
R1530 VCC.n668 VCC.n667 4.5005
R1531 VCC.n198 VCC.n195 4.5005
R1532 VCC.n660 VCC.n659 4.5005
R1533 VCC.n653 VCC.n142 4.5005
R1534 VCC.n160 VCC.n158 4.5005
R1535 VCC.n644 VCC.n643 4.5005
R1536 VCC.n237 VCC.n236 4.5005
R1537 VCC.n237 VCC.n230 4.5005
R1538 VCC.n638 VCC.n637 4.5005
R1539 VCC.n250 VCC.n249 4.5005
R1540 VCC.n248 VCC.n175 4.5005
R1541 VCC.n248 VCC.n247 4.5005
R1542 VCC.n645 VCC.n150 4.5005
R1543 VCC.n652 VCC.n651 4.5005
R1544 VCC.n208 VCC.n207 4.5005
R1545 VCC.n207 VCC.n185 4.5005
R1546 VCC.n206 VCC.n139 4.5005
R1547 VCC.n204 VCC.n203 4.5005
R1548 VCC.n201 VCC.n200 4.5005
R1549 VCC.n630 VCC.n629 4.5005
R1550 VCC.n622 VCC.n265 4.31039
R1551 VCC.n259 VCC.n168 4.31039
R1552 VCC.n544 VCC.n300 3.51902
R1553 VCC.n597 VCC.n281 3.51902
R1554 VCC.n218 VCC.n183 3.51902
R1555 VCC.n241 VCC.n179 3.51902
R1556 VCC.n387 VCC.n386 3.42479
R1557 VCC.n732 VCC.n731 3.42479
R1558 VCC.n520 VCC.n519 3.42389
R1559 VCC.n522 VCC.n521 3.42389
R1560 VCC.n131 VCC.n130 3.42389
R1561 VCC.n667 VCC.n132 3.42389
R1562 VCC.n626 VCC.n625 3.423
R1563 VCC.n629 VCC.n628 3.423
R1564 VCC.n610 VCC.n609 3.4105
R1565 VCC.n610 VCC.n263 3.4105
R1566 VCC.n586 VCC.n585 3.4105
R1567 VCC.n608 VCC.n607 3.4105
R1568 VCC.n607 VCC.n606 3.4105
R1569 VCC.n576 VCC.n292 3.4105
R1570 VCC.n292 VCC.n291 3.4105
R1571 VCC.n578 VCC.n577 3.4105
R1572 VCC.n584 VCC.n583 3.4105
R1573 VCC.n583 VCC.n582 3.4105
R1574 VCC.n558 VCC.n557 3.4105
R1575 VCC.n558 VCC.n304 3.4105
R1576 VCC.n554 VCC.n294 3.4105
R1577 VCC.n575 VCC.n574 3.4105
R1578 VCC.n574 VCC.n573 3.4105
R1579 VCC.n536 VCC.n533 3.4105
R1580 VCC.n536 VCC.n535 3.4105
R1581 VCC.n553 VCC.n552 3.4105
R1582 VCC.n532 VCC.n531 3.4105
R1583 VCC.n531 VCC.n530 3.4105
R1584 VCC.n516 VCC.n515 3.4105
R1585 VCC.n517 VCC.n516 3.4105
R1586 VCC.n481 VCC.n480 3.4105
R1587 VCC.n514 VCC.n513 3.4105
R1588 VCC.n513 VCC.n512 3.4105
R1589 VCC.n451 VCC.n450 3.4105
R1590 VCC.n450 VCC.n449 3.4105
R1591 VCC.n446 VCC.n444 3.4105
R1592 VCC.n479 VCC.n478 3.4105
R1593 VCC.n478 VCC.n477 3.4105
R1594 VCC.n362 VCC.n361 3.4105
R1595 VCC.n422 VCC.n362 3.4105
R1596 VCC.n443 VCC.n359 3.4105
R1597 VCC.n453 VCC.n452 3.4105
R1598 VCC.n453 VCC.n358 3.4105
R1599 VCC.n416 VCC.n373 3.4105
R1600 VCC.n416 VCC.n415 3.4105
R1601 VCC.n420 VCC.n419 3.4105
R1602 VCC.n390 VCC.n389 3.4105
R1603 VCC.n390 VCC.n384 3.4105
R1604 VCC.n640 VCC.n639 3.4105
R1605 VCC.n635 VCC.n634 3.4105
R1606 VCC.n636 VCC.n635 3.4105
R1607 VCC.n648 VCC.n647 3.4105
R1608 VCC.n647 VCC.n646 3.4105
R1609 VCC.n153 VCC.n149 3.4105
R1610 VCC.n642 VCC.n641 3.4105
R1611 VCC.n642 VCC.n152 3.4105
R1612 VCC.n656 VCC.n655 3.4105
R1613 VCC.n655 VCC.n654 3.4105
R1614 VCC.n148 VCC.n146 3.4105
R1615 VCC.n650 VCC.n649 3.4105
R1616 VCC.n650 VCC.n144 3.4105
R1617 VCC.n663 VCC.n662 3.4105
R1618 VCC.n662 VCC.n661 3.4105
R1619 VCC.n658 VCC.n657 3.4105
R1620 VCC.n127 VCC.n126 3.4105
R1621 VCC.n128 VCC.n127 3.4105
R1622 VCC.n692 VCC.n66 3.4105
R1623 VCC.n125 VCC.n124 3.4105
R1624 VCC.n124 VCC.n123 3.4105
R1625 VCC.n704 VCC.n60 3.4105
R1626 VCC.n705 VCC.n704 3.4105
R1627 VCC.n702 VCC.n701 3.4105
R1628 VCC.n699 VCC.n698 3.4105
R1629 VCC.n698 VCC.n697 3.4105
R1630 VCC.n59 VCC.n43 3.4105
R1631 VCC.n43 VCC.n41 3.4105
R1632 VCC.n710 VCC.n44 3.4105
R1633 VCC.n709 VCC.n708 3.4105
R1634 VCC.n708 VCC.n707 3.4105
R1635 VCC.n727 VCC.n726 3.4105
R1636 VCC.n726 VCC.n725 3.4105
R1637 VCC.n58 VCC.n57 3.4105
R1638 VCC.n729 VCC.n728 3.4105
R1639 VCC.n730 VCC.n729 3.4105
R1640 VCC.n664 VCC.n133 3.4105
R1641 VCC.n133 VCC.n115 3.4105
R1642 VCC.n633 VCC.n632 3.4105
R1643 VCC.n632 VCC.n631 3.4105
R1644 VCC.n493 VCC.n316 3.29193
R1645 VCC.n548 VCC.n547 3.29193
R1646 VCC.n587 VCC.n279 3.29193
R1647 VCC.n193 VCC.n192 3.29193
R1648 VCC.n213 VCC.n212 3.29193
R1649 VCC.n232 VCC.n177 3.29193
R1650 VCC.n541 VCC.n314 3.25764
R1651 VCC.n600 VCC.n267 3.25764
R1652 VCC.n215 VCC.n189 3.25764
R1653 VCC.n244 VCC.n170 3.25764
R1654 VCC.n619 VCC.n618 3.2005
R1655 VCC.n256 VCC.n255 3.2005
R1656 VCC.n540 VCC.n539 3.03311
R1657 VCC.n572 VCC.n571 3.03311
R1658 VCC.n181 VCC.n151 3.03311
R1659 VCC.n205 VCC.n204 3.03311
R1660 VCC.n795 VCC.n794 2.8505
R1661 VCC.n855 VCC.n854 2.8505
R1662 VCC.n410 VCC.n378 2.8505
R1663 VCC.n488 VCC.n339 2.8505
R1664 VCC.n34 VCC.n11 2.8505
R1665 VCC.n683 VCC.n77 2.8505
R1666 VCC.n471 VCC.n470 2.5605
R1667 VCC.n97 VCC.n96 2.5605
R1668 VCC.n430 VCC.n429 2.46907
R1669 VCC.n49 VCC.n39 2.46907
R1670 VCC.n486 VCC.n337 2.37764
R1671 VCC.n682 VCC.n681 2.37764
R1672 VCC.n774 VCC.n773 2.34304
R1673 VCC.n340 VCC.n338 2.34304
R1674 VCC.n382 VCC.n380 2.34304
R1675 VCC.n673 VCC.n109 2.34304
R1676 VCC.n22 VCC.n18 2.34304
R1677 VCC.n398 VCC.n377 2.28621
R1678 VCC.n33 VCC.n32 2.28621
R1679 VCC.n328 VCC.n327 2.2505
R1680 VCC.n511 VCC.n331 2.2505
R1681 VCC.n476 VCC.n348 2.2505
R1682 VCC.n404 VCC.n391 2.2505
R1683 VCC.n375 VCC.n374 2.2505
R1684 VCC.n423 VCC.n421 2.2505
R1685 VCC.n613 VCC.n612 2.2505
R1686 VCC.n605 VCC.n274 2.2505
R1687 VCC.n287 VCC.n285 2.2505
R1688 VCC.n529 VCC.n323 2.2505
R1689 VCC.n537 VCC.n318 2.2505
R1690 VCC.n560 VCC.n559 2.2505
R1691 VCC.n108 VCC.n107 2.2505
R1692 VCC.n122 VCC.n119 2.2505
R1693 VCC.n696 VCC.n68 2.2505
R1694 VCC.n3 VCC.n2 2.2505
R1695 VCC.n7 VCC.n5 2.2505
R1696 VCC.n52 VCC.n51 2.2505
R1697 VCC.n166 VCC.n164 2.2505
R1698 VCC.n137 VCC.n135 2.2505
R1699 VCC.n143 VCC.n141 2.2505
R1700 VCC.n231 VCC.n155 2.2505
R1701 VCC.n162 VCC.n161 2.2505
R1702 VCC.n197 VCC.n196 2.2505
R1703 VCC.n627 VCC 2.24168
R1704 VCC.n458 VCC.n457 2.10336
R1705 VCC.n88 VCC.n87 2.10336
R1706 VCC.n828 VCC.n827 2.01193
R1707 VCC.n457 VCC.n456 2.01193
R1708 VCC.n87 VCC.n84 2.01193
R1709 VCC.n624 VCC.n623 2.00996
R1710 VCC.n630 VCC.n260 2.00996
R1711 VCC.n523 VCC.n324 1.98102
R1712 VCC.n669 VCC.n668 1.98102
R1713 VCC.n817 VCC.n816 1.82742
R1714 VCC.n878 VCC.n877 1.82742
R1715 VCC.n433 VCC.n432 1.82742
R1716 VCC.n468 VCC.n467 1.82742
R1717 VCC.n720 VCC.n719 1.82742
R1718 VCC.n101 VCC.n100 1.82742
R1719 VCC.n564 VCC.n301 1.62907
R1720 VCC.n596 VCC.n282 1.62907
R1721 VCC.n219 VCC.n184 1.62907
R1722 VCC.n240 VCC.n180 1.62907
R1723 VCC.n540 VCC.n316 1.55479
R1724 VCC.n205 VCC.n193 1.55479
R1725 VCC.n891 VCC.n890 1.5005
R1726 VCC.n820 VCC.n813 1.46336
R1727 VCC.n881 VCC.n872 1.46336
R1728 VCC.n436 VCC.n365 1.46336
R1729 VCC.n464 VCC.n350 1.46336
R1730 VCC.n602 VCC.n268 1.46336
R1731 VCC.n717 VCC.n716 1.46336
R1732 VCC.n98 VCC.n94 1.46336
R1733 VCC.n247 VCC.n171 1.46336
R1734 VCC.n548 VCC.n302 1.37193
R1735 VCC.n563 VCC.n298 1.37193
R1736 VCC.n570 VCC.n283 1.37193
R1737 VCC.n587 VCC.n284 1.37193
R1738 VCC.n212 VCC.n185 1.37193
R1739 VCC.n222 VCC.n221 1.37193
R1740 VCC.n229 VCC.n228 1.37193
R1741 VCC.n232 VCC.n230 1.37193
R1742 VCC.n800 VCC.n793 1.2805
R1743 VCC.n860 VCC.n853 1.2805
R1744 VCC.n413 VCC.n411 1.2805
R1745 VCC.n487 VCC.n485 1.2805
R1746 VCC.n723 VCC.n9 1.2805
R1747 VCC.n688 VCC.n75 1.2805
R1748 VCC.n547 VCC.n313 1.18907
R1749 VCC.n601 VCC.n279 1.18907
R1750 VCC.n214 VCC.n213 1.18907
R1751 VCC.n245 VCC.n177 1.18907
R1752 VCC.n388 VCC.n385 1.13717
R1753 VCC.n418 VCC.n417 1.13717
R1754 VCC.n442 VCC.n441 1.13717
R1755 VCC.n445 VCC.n346 1.13717
R1756 VCC.n330 VCC.n329 1.13717
R1757 VCC.n326 VCC.n325 1.13717
R1758 VCC.n322 VCC.n321 1.13717
R1759 VCC.n320 VCC.n308 1.13717
R1760 VCC.n556 VCC.n555 1.13717
R1761 VCC.n293 VCC.n289 1.13717
R1762 VCC.n273 VCC.n272 1.13717
R1763 VCC.n262 VCC.n261 1.13717
R1764 VCC.n165 VCC.n163 1.13717
R1765 VCC.n918 VCC.n917 1.13717
R1766 VCC.n908 VCC.n907 1.13717
R1767 VCC.n897 VCC.n896 1.13717
R1768 VCC.n762 VCC.n761 1.13717
R1769 VCC.n750 VCC.n749 1.13717
R1770 VCC.n739 VCC.n738 1.13717
R1771 VCC.n1 VCC.n0 1.13717
R1772 VCC.n6 VCC.n4 1.13717
R1773 VCC.n712 VCC.n711 1.13717
R1774 VCC.n700 VCC.n65 1.13717
R1775 VCC.n118 VCC.n71 1.13717
R1776 VCC.n117 VCC.n116 1.13717
R1777 VCC.n666 VCC.n665 1.13717
R1778 VCC.n136 VCC.n134 1.13717
R1779 VCC.n145 VCC.n140 1.13717
R1780 VCC.n156 VCC.n154 1.13717
R1781 VCC.n159 VCC.n157 1.13717
R1782 VCC.n448 VCC.n360 1.1255
R1783 VCC.n572 VCC.n296 1.1255
R1784 VCC.n706 VCC.n62 1.1255
R1785 VCC.n151 VCC.n147 1.1255
R1786 VCC.n782 VCC.n779 1.00621
R1787 VCC.n781 VCC.n780 1.00621
R1788 VCC.n882 VCC.n870 1.00621
R1789 VCC.n405 VCC.n383 1.00621
R1790 VCC.n398 VCC.n397 1.00621
R1791 VCC.n463 VCC.n354 1.00621
R1792 VCC.n494 VCC.n493 1.00621
R1793 VCC.n619 VCC.n264 1.00621
R1794 VCC.n24 VCC.n23 1.00621
R1795 VCC.n32 VCC.n14 1.00621
R1796 VCC.n93 VCC.n80 1.00621
R1797 VCC.n192 VCC.n114 1.00621
R1798 VCC.n256 VCC.n167 1.00621
R1799 VCC.n815 VCC.n814 0.9505
R1800 VCC.n875 VCC.n874 0.9505
R1801 VCC.n431 VCC.n366 0.9505
R1802 VCC.n469 VCC.n351 0.9505
R1803 VCC.n718 VCC.n12 0.9505
R1804 VCC.n99 VCC.n76 0.9505
R1805 VCC.n822 VCC.n821 0.914786
R1806 VCC.n887 VCC.n886 0.914786
R1807 VCC.n837 VCC.n836 0.914786
R1808 VCC.n840 VCC.n839 0.914786
R1809 VCC.n438 VCC.n437 0.914786
R1810 VCC.n456 VCC.n356 0.914786
R1811 VCC.n504 VCC.n337 0.914786
R1812 VCC.n503 VCC.n502 0.914786
R1813 VCC.n81 VCC.n40 0.914786
R1814 VCC.n84 VCC.n83 0.914786
R1815 VCC.n681 VCC.n103 0.914786
R1816 VCC.n675 VCC.n674 0.914786
R1817 VCC.n803 VCC.n800 0.823357
R1818 VCC.n802 VCC.n801 0.823357
R1819 VCC.n828 VCC.n826 0.823357
R1820 VCC.n861 VCC.n851 0.823357
R1821 VCC.n413 VCC.n412 0.823357
R1822 VCC.n429 VCC.n369 0.823357
R1823 VCC.n459 VCC.n458 0.823357
R1824 VCC.n484 VCC.n343 0.823357
R1825 VCC.n723 VCC.n10 0.823357
R1826 VCC.n49 VCC.n48 0.823357
R1827 VCC.n89 VCC.n88 0.823357
R1828 VCC.n689 VCC.n74 0.823357
R1829 VCC.n803 VCC.n802 0.731929
R1830 VCC.n851 VCC.n850 0.731929
R1831 VCC.n861 VCC.n860 0.731929
R1832 VCC.n412 VCC.n369 0.731929
R1833 VCC.n471 VCC.n343 0.731929
R1834 VCC.n485 VCC.n484 0.731929
R1835 VCC.n48 VCC.n10 0.731929
R1836 VCC.n96 VCC.n74 0.731929
R1837 VCC.n689 VCC.n688 0.731929
R1838 VCC.n822 VCC.n820 0.6405
R1839 VCC.n840 VCC.n837 0.6405
R1840 VCC.n438 VCC.n436 0.6405
R1841 VCC.n504 VCC.n503 0.6405
R1842 VCC.n716 VCC.n40 0.6405
R1843 VCC.n675 VCC.n103 0.6405
R1844 VCC.n782 VCC.n781 0.549071
R1845 VCC.n882 VCC.n881 0.549071
R1846 VCC.n397 VCC.n383 0.549071
R1847 VCC.n464 VCC.n463 0.549071
R1848 VCC.n24 VCC.n14 0.549071
R1849 VCC.n94 VCC.n93 0.549071
R1850 VCC.n521 VCC 0.535293
R1851 VCC.n132 VCC 0.535293
R1852 VCC.n623 VCC.n264 0.507747
R1853 VCC.n260 VCC.n167 0.507747
R1854 VCC.n494 VCC.n324 0.465115
R1855 VCC.n669 VCC.n114 0.465115
R1856 VCC.n540 VCC.n313 0.366214
R1857 VCC.n603 VCC.n601 0.366214
R1858 VCC.n214 VCC.n205 0.366214
R1859 VCC.n246 VCC.n245 0.366214
R1860 VCC VCC.n626 0.300964
R1861 VCC.n628 VCC 0.300964
R1862 VCC.n387 VCC 0.294921
R1863 VCC VCC.n919 0.294921
R1864 VCC VCC.n732 0.287536
R1865 VCC.n793 VCC.n792 0.274786
R1866 VCC.n853 VCC.n852 0.274786
R1867 VCC.n411 VCC.n377 0.274786
R1868 VCC.n437 VCC.n356 0.274786
R1869 VCC.n459 VCC.n354 0.274786
R1870 VCC.n487 VCC.n486 0.274786
R1871 VCC.n33 VCC.n9 0.274786
R1872 VCC.n83 VCC.n81 0.274786
R1873 VCC.n89 VCC.n80 0.274786
R1874 VCC.n682 VCC.n75 0.274786
R1875 VCC.n733 VCC 0.213679
R1876 VCC.n562 VCC.n302 0.183357
R1877 VCC.n563 VCC.n562 0.183357
R1878 VCC.n595 VCC.n283 0.183357
R1879 VCC.n595 VCC.n284 0.183357
R1880 VCC.n220 VCC.n185 0.183357
R1881 VCC.n221 VCC.n220 0.183357
R1882 VCC.n239 VCC.n229 0.183357
R1883 VCC.n239 VCC.n230 0.183357
R1884 VCC VCC.n520 0.114307
R1885 VCC VCC.n131 0.114307
R1886 VCC.n813 VCC.n812 0.0919286
R1887 VCC.n872 VCC.n871 0.0919286
R1888 VCC.n430 VCC.n365 0.0919286
R1889 VCC.n470 VCC.n350 0.0919286
R1890 VCC.n603 VCC.n602 0.0919286
R1891 VCC.n618 VCC.n268 0.0919286
R1892 VCC.n717 VCC.n39 0.0919286
R1893 VCC.n98 VCC.n97 0.0919286
R1894 VCC.n247 VCC.n246 0.0919286
R1895 VCC.n255 VCC.n171 0.0919286
R1896 VCC VCC.n627 0.0246714
R1897 VCC.n389 VCC.n373 0.024
R1898 VCC.n515 VCC.n514 0.024
R1899 VCC.n533 VCC.n532 0.024
R1900 VCC.n609 VCC.n608 0.024
R1901 VCC.n910 VCC.n909 0.024
R1902 VCC.n741 VCC.n740 0.024
R1903 VCC.n728 VCC.n727 0.024
R1904 VCC.n126 VCC.n125 0.024
R1905 VCC.n664 VCC.n663 0.024
R1906 VCC.n634 VCC.n633 0.024
R1907 VCC.n306 VCC.n297 0.0228214
R1908 VCC.n581 VCC.n580 0.0228214
R1909 VCC.n589 VCC.n275 0.0228214
R1910 VCC.n653 VCC.n652 0.0228214
R1911 VCC.n645 VCC.n644 0.0228214
R1912 VCC.n637 VCC.n160 0.0228214
R1913 VCC.n627 VCC 0.0199714
R1914 VCC.n890 VCC.n889 0.0174643
R1915 VCC.n448 VCC.n358 0.0174643
R1916 VCC.n449 VCC.n448 0.0174643
R1917 VCC.n453 VCC.n360 0.0174643
R1918 VCC.n450 VCC.n360 0.0174643
R1919 VCC.n573 VCC.n572 0.0174643
R1920 VCC.n572 VCC.n291 0.0174643
R1921 VCC.n574 VCC.n296 0.0174643
R1922 VCC.n296 VCC.n292 0.0174643
R1923 VCC.n707 VCC.n706 0.0174643
R1924 VCC.n706 VCC.n705 0.0174643
R1925 VCC.n708 VCC.n62 0.0174643
R1926 VCC.n704 VCC.n62 0.0174643
R1927 VCC.n151 VCC.n144 0.0174643
R1928 VCC.n646 VCC.n151 0.0174643
R1929 VCC.n650 VCC.n147 0.0174643
R1930 VCC.n647 VCC.n147 0.0174643
R1931 VCC.n807 VCC.n806 0.0165714
R1932 VCC.n831 VCC.n830 0.0165714
R1933 VCC.n913 VCC.n912 0.0165714
R1934 VCC.n905 VCC.n904 0.0165714
R1935 VCC.n893 VCC.n892 0.0165714
R1936 VCC.n745 VCC.n744 0.0165714
R1937 VCC.n473 VCC.n472 0.0165714
R1938 VCC.n401 VCC.n393 0.0165714
R1939 VCC.n426 VCC.n420 0.0165714
R1940 VCC.n481 VCC.n345 0.0165714
R1941 VCC.n508 VCC.n507 0.0165714
R1942 VCC.n526 VCC.n319 0.0165714
R1943 VCC.n586 VCC.n288 0.0165714
R1944 VCC.n615 VCC.n271 0.0165714
R1945 VCC.n95 VCC.n70 0.0165714
R1946 VCC.n29 VCC.n27 0.0165714
R1947 VCC.n57 VCC.n56 0.0165714
R1948 VCC.n693 VCC.n692 0.0165714
R1949 VCC.n678 VCC.n106 0.0165714
R1950 VCC.n202 VCC.n201 0.0165714
R1951 VCC.n639 VCC.n638 0.0165714
R1952 VCC.n252 VCC.n250 0.0165714
R1953 VCC.n865 VCC.n864 0.0156786
R1954 VCC.n906 VCC.n905 0.0156786
R1955 VCC.n428 VCC.n427 0.0156786
R1956 VCC.n482 VCC.n481 0.0156786
R1957 VCC.n552 VCC.n309 0.0156786
R1958 VCC.n55 VCC.n50 0.0156786
R1959 VCC.n692 VCC.n691 0.0156786
R1960 VCC.n659 VCC.n658 0.0156786
R1961 VCC.n419 VCC.n361 0.0152714
R1962 VCC.n480 VCC.n479 0.0152714
R1963 VCC.n557 VCC.n553 0.0152714
R1964 VCC.n585 VCC.n584 0.0152714
R1965 VCC.n899 VCC.n898 0.0152714
R1966 VCC.n752 VCC.n751 0.0152714
R1967 VCC.n59 VCC.n58 0.0152714
R1968 VCC.n699 VCC.n66 0.0152714
R1969 VCC.n657 VCC.n656 0.0152714
R1970 VCC.n641 VCC.n640 0.0152714
R1971 VCC.n743 VCC.n742 0.0147857
R1972 VCC.n420 VCC.n372 0.0147857
R1973 VCC.n534 VCC.n311 0.0147857
R1974 VCC.n57 VCC.n45 0.0147857
R1975 VCC.n660 VCC.n138 0.0147857
R1976 VCC.n452 VCC.n451 0.0132571
R1977 VCC.n576 VCC.n575 0.0132571
R1978 VCC.n765 VCC.n764 0.0132571
R1979 VCC.n709 VCC.n60 0.0132571
R1980 VCC.n649 VCC.n648 0.0132571
R1981 VCC.n787 VCC.n786 0.013
R1982 VCC.n335 VCC.n333 0.013
R1983 VCC.n616 VCC.n270 0.013
R1984 VCC.n624 VCC.n263 0.013
R1985 VCC.n615 VCC.n614 0.013
R1986 VCC.n680 VCC.n104 0.013
R1987 VCC.n253 VCC.n174 0.013
R1988 VCC.n631 VCC.n630 0.013
R1989 VCC.n252 VCC.n251 0.013
R1990 VCC.n845 VCC.n844 0.0121071
R1991 VCC.n914 VCC.n913 0.0121071
R1992 VCC.n399 VCC.n396 0.0121071
R1993 VCC.n518 VCC.n517 0.0121071
R1994 VCC.n507 VCC.n334 0.0121071
R1995 VCC.n530 VCC.n523 0.0121071
R1996 VCC.n528 VCC.n525 0.0121071
R1997 VCC.n527 VCC.n526 0.0121071
R1998 VCC.n277 VCC.n274 0.0121071
R1999 VCC.n31 VCC.n30 0.0121071
R2000 VCC.n129 VCC.n128 0.0121071
R2001 VCC.n678 VCC.n677 0.0121071
R2002 VCC.n668 VCC.n115 0.0121071
R2003 VCC.n200 VCC.n198 0.0121071
R2004 VCC.n201 VCC.n195 0.0121071
R2005 VCC.n175 VCC.n162 0.0121071
R2006 VCC.n789 VCC.n788 0.0112143
R2007 VCC.n846 VCC.n845 0.0112143
R2008 VCC.n833 VCC.n832 0.0112143
R2009 VCC.n901 VCC.n900 0.0112143
R2010 VCC.n746 VCC.n745 0.0112143
R2011 VCC.n396 VCC.n395 0.0112143
R2012 VCC.n511 VCC.n510 0.0112143
R2013 VCC.n402 VCC.n401 0.0112143
R2014 VCC.n394 VCC.n393 0.0112143
R2015 VCC.n509 VCC.n331 0.0112143
R2016 VCC.n525 VCC.n524 0.0112143
R2017 VCC.n539 VCC.n318 0.0112143
R2018 VCC.n605 VCC.n604 0.0112143
R2019 VCC.n538 VCC.n537 0.0112143
R2020 VCC.n30 VCC.n16 0.0112143
R2021 VCC.n122 VCC.n121 0.0112143
R2022 VCC.n27 VCC.n26 0.0112143
R2023 VCC.n29 VCC.n28 0.0112143
R2024 VCC.n120 VCC.n119 0.0112143
R2025 VCC.n200 VCC.n199 0.0112143
R2026 VCC.n204 VCC.n137 0.0112143
R2027 VCC.n176 VCC.n161 0.0112143
R2028 VCC.n203 VCC.n135 0.0112143
R2029 VCC.n788 VCC.n787 0.0103214
R2030 VCC.n811 VCC.n810 0.0103214
R2031 VCC.n884 VCC.n883 0.0103214
R2032 VCC.n868 VCC.n867 0.0103214
R2033 VCC.n847 VCC.n846 0.0103214
R2034 VCC.n768 VCC.n767 0.0103214
R2035 VCC.n759 VCC.n758 0.0103214
R2036 VCC.n747 VCC.n746 0.0103214
R2037 VCC.n735 VCC.n734 0.0103214
R2038 VCC.n404 VCC.n403 0.0103214
R2039 VCC.n395 VCC.n375 0.0103214
R2040 VCC.n423 VCC.n422 0.0103214
R2041 VCC.n462 VCC.n461 0.0103214
R2042 VCC.n477 VCC.n476 0.0103214
R2043 VCC.n510 VCC.n333 0.0103214
R2044 VCC.n402 VCC.n391 0.0103214
R2045 VCC.n394 VCC.n374 0.0103214
R2046 VCC.n421 VCC.n362 0.0103214
R2047 VCC.n478 VCC.n348 0.0103214
R2048 VCC.n509 VCC.n508 0.0103214
R2049 VCC.n539 VCC.n317 0.0103214
R2050 VCC.n535 VCC.n534 0.0103214
R2051 VCC.n560 VCC.n304 0.0103214
R2052 VCC.n582 VCC.n285 0.0103214
R2053 VCC.n617 VCC.n616 0.0103214
R2054 VCC.n538 VCC.n319 0.0103214
R2055 VCC.n559 VCC.n558 0.0103214
R2056 VCC.n554 VCC.n295 0.0103214
R2057 VCC.n583 VCC.n287 0.0103214
R2058 VCC.n591 VCC.n590 0.0103214
R2059 VCC.n25 VCC.n2 0.0103214
R2060 VCC.n16 VCC.n7 0.0103214
R2061 VCC.n52 VCC.n41 0.0103214
R2062 VCC.n92 VCC.n91 0.0103214
R2063 VCC.n697 VCC.n696 0.0103214
R2064 VCC.n121 VCC.n104 0.0103214
R2065 VCC.n26 VCC.n3 0.0103214
R2066 VCC.n28 VCC.n5 0.0103214
R2067 VCC.n51 VCC.n43 0.0103214
R2068 VCC.n698 VCC.n68 0.0103214
R2069 VCC.n120 VCC.n106 0.0103214
R2070 VCC.n204 VCC.n194 0.0103214
R2071 VCC.n661 VCC.n660 0.0103214
R2072 VCC.n654 VCC.n143 0.0103214
R2073 VCC.n231 VCC.n152 0.0103214
R2074 VCC.n254 VCC.n253 0.0103214
R2075 VCC.n203 VCC.n202 0.0103214
R2076 VCC.n655 VCC.n141 0.0103214
R2077 VCC.n651 VCC.n146 0.0103214
R2078 VCC.n642 VCC.n155 0.0103214
R2079 VCC.n235 VCC.n158 0.0103214
R2080 VCC.n783 VCC.n772 0.00942857
R2081 VCC.n824 VCC.n823 0.00942857
R2082 VCC.n888 VCC.n885 0.00942857
R2083 VCC.n841 VCC.n835 0.00942857
R2084 VCC.n915 VCC.n914 0.00942857
R2085 VCC.n755 VCC.n754 0.00942857
R2086 VCC.n439 VCC.n364 0.00942857
R2087 VCC.n455 VCC.n357 0.00942857
R2088 VCC.n336 VCC.n327 0.00942857
R2089 VCC.n454 VCC.n359 0.00942857
R2090 VCC.n334 VCC.n328 0.00942857
R2091 VCC.n529 VCC.n528 0.00942857
R2092 VCC.n606 VCC.n275 0.00942857
R2093 VCC.n278 VCC.n276 0.00942857
R2094 VCC.n527 VCC.n323 0.00942857
R2095 VCC.n551 VCC.n310 0.00942857
R2096 VCC.n579 VCC.n578 0.00942857
R2097 VCC.n277 VCC.n271 0.00942857
R2098 VCC.n714 VCC.n42 0.00942857
R2099 VCC.n82 VCC.n63 0.00942857
R2100 VCC.n676 VCC.n108 0.00942857
R2101 VCC.n61 VCC.n44 0.00942857
R2102 VCC.n677 VCC.n107 0.00942857
R2103 VCC.n198 VCC.n197 0.00942857
R2104 VCC.n637 VCC.n636 0.00942857
R2105 VCC.n249 VCC.n248 0.00942857
R2106 VCC.n196 VCC.n195 0.00942857
R2107 VCC.n209 VCC.n139 0.00942857
R2108 VCC.n153 VCC.n150 0.00942857
R2109 VCC.n250 VCC.n175 0.00942857
R2110 VCC.n804 VCC.n791 0.00853571
R2111 VCC.n806 VCC.n805 0.00853571
R2112 VCC.n829 VCC.n825 0.00853571
R2113 VCC.n863 VCC.n862 0.00853571
R2114 VCC.n895 VCC.n894 0.00853571
R2115 VCC.n414 VCC.n376 0.00853571
R2116 VCC.n428 VCC.n370 0.00853571
R2117 VCC.n460 VCC.n355 0.00853571
R2118 VCC.n483 VCC.n344 0.00853571
R2119 VCC.n447 VCC.n446 0.00853571
R2120 VCC.n550 VCC.n311 0.00853571
R2121 VCC.n614 VCC.n613 0.00853571
R2122 VCC.n625 VCC.n262 0.00853571
R2123 VCC.n724 VCC.n8 0.00853571
R2124 VCC.n50 VCC.n47 0.00853571
R2125 VCC.n90 VCC.n64 0.00853571
R2126 VCC.n690 VCC.n72 0.00853571
R2127 VCC.n703 VCC.n702 0.00853571
R2128 VCC.n206 VCC.n138 0.00853571
R2129 VCC.n251 VCC.n164 0.00853571
R2130 VCC.n629 VCC.n165 0.00853571
R2131 VCC.n388 VCC.n387 0.00822143
R2132 VCC.n419 VCC.n418 0.00822143
R2133 VCC.n480 VCC.n329 0.00822143
R2134 VCC.n520 VCC.n325 0.00822143
R2135 VCC.n521 VCC.n321 0.00822143
R2136 VCC.n553 VCC.n308 0.00822143
R2137 VCC.n585 VCC.n272 0.00822143
R2138 VCC.n626 VCC.n261 0.00822143
R2139 VCC.n919 VCC.n918 0.00822143
R2140 VCC.n908 VCC.n899 0.00822143
R2141 VCC.n751 VCC.n750 0.00822143
R2142 VCC.n739 VCC.n733 0.00822143
R2143 VCC.n732 VCC.n0 0.00822143
R2144 VCC.n58 VCC.n4 0.00822143
R2145 VCC.n118 VCC.n66 0.00822143
R2146 VCC.n131 VCC.n116 0.00822143
R2147 VCC.n665 VCC.n132 0.00822143
R2148 VCC.n657 VCC.n134 0.00822143
R2149 VCC.n640 VCC.n157 0.00822143
R2150 VCC.n628 VCC.n163 0.00822143
R2151 VCC.n805 VCC.n804 0.00764286
R2152 VCC.n810 VCC.n809 0.00764286
R2153 VCC.n866 VCC.n865 0.00764286
R2154 VCC.n864 VCC.n863 0.00764286
R2155 VCC.n862 VCC.n849 0.00764286
R2156 VCC.n917 VCC.n911 0.00764286
R2157 VCC.n896 VCC.n895 0.00764286
R2158 VCC.n761 VCC.n755 0.00764286
R2159 VCC.n760 VCC.n759 0.00764286
R2160 VCC.n757 VCC.n756 0.00764286
R2161 VCC.n376 VCC.n370 0.00764286
R2162 VCC.n476 VCC.n475 0.00764286
R2163 VCC.n472 VCC.n344 0.00764286
R2164 VCC.n483 VCC.n332 0.00764286
R2165 VCC.n426 VCC.n425 0.00764286
R2166 VCC.n440 VCC.n362 0.00764286
R2167 VCC.n441 VCC.n359 0.00764286
R2168 VCC.n446 VCC.n445 0.00764286
R2169 VCC.n474 VCC.n348 0.00764286
R2170 VCC.n519 VCC.n326 0.00764286
R2171 VCC.n549 VCC.n312 0.00764286
R2172 VCC.n588 VCC.n286 0.00764286
R2173 VCC.n522 VCC.n322 0.00764286
R2174 VCC.n552 VCC.n551 0.00764286
R2175 VCC.n559 VCC.n305 0.00764286
R2176 VCC.n555 VCC.n554 0.00764286
R2177 VCC.n578 VCC.n293 0.00764286
R2178 VCC.n592 VCC.n287 0.00764286
R2179 VCC.n47 VCC.n8 0.00764286
R2180 VCC.n696 VCC.n695 0.00764286
R2181 VCC.n95 VCC.n72 0.00764286
R2182 VCC.n690 VCC.n73 0.00764286
R2183 VCC.n56 VCC.n46 0.00764286
R2184 VCC.n713 VCC.n43 0.00764286
R2185 VCC.n712 VCC.n44 0.00764286
R2186 VCC.n702 VCC.n65 0.00764286
R2187 VCC.n694 VCC.n68 0.00764286
R2188 VCC.n130 VCC.n117 0.00764286
R2189 VCC.n211 VCC.n210 0.00764286
R2190 VCC.n234 VCC.n233 0.00764286
R2191 VCC.n667 VCC.n666 0.00764286
R2192 VCC.n658 VCC.n139 0.00764286
R2193 VCC.n208 VCC.n141 0.00764286
R2194 VCC.n146 VCC.n145 0.00764286
R2195 VCC.n154 VCC.n153 0.00764286
R2196 VCC.n236 VCC.n155 0.00764286
R2197 VCC.n785 VCC.n784 0.00675
R2198 VCC.n823 VCC.n811 0.00675
R2199 VCC.n867 VCC.n866 0.00675
R2200 VCC.n842 VCC.n841 0.00675
R2201 VCC.n904 VCC.n903 0.00675
R2202 VCC.n769 VCC.n768 0.00675
R2203 VCC.n758 VCC.n757 0.00675
R2204 VCC.n749 VCC.n743 0.00675
R2205 VCC.n738 VCC.n737 0.00675
R2206 VCC.n424 VCC.n423 0.00675
R2207 VCC.n439 VCC.n363 0.00675
R2208 VCC.n475 VCC.n473 0.00675
R2209 VCC.n505 VCC.n336 0.00675
R2210 VCC.n386 VCC.n385 0.00675
R2211 VCC.n417 VCC.n372 0.00675
R2212 VCC.n425 VCC.n421 0.00675
R2213 VCC.n478 VCC.n347 0.00675
R2214 VCC.n474 VCC.n345 0.00675
R2215 VCC.n312 VCC.n303 0.00675
R2216 VCC.n306 VCC.n304 0.00675
R2217 VCC.n593 VCC.n286 0.00675
R2218 VCC.n310 VCC.n305 0.00675
R2219 VCC.n558 VCC.n307 0.00675
R2220 VCC.n293 VCC.n290 0.00675
R2221 VCC.n592 VCC.n591 0.00675
R2222 VCC.n590 VCC.n586 0.00675
R2223 VCC.n53 VCC.n52 0.00675
R2224 VCC.n715 VCC.n714 0.00675
R2225 VCC.n695 VCC.n70 0.00675
R2226 VCC.n676 VCC.n105 0.00675
R2227 VCC.n731 VCC.n1 0.00675
R2228 VCC.n45 VCC.n6 0.00675
R2229 VCC.n51 VCC.n46 0.00675
R2230 VCC.n698 VCC.n67 0.00675
R2231 VCC.n694 VCC.n693 0.00675
R2232 VCC.n210 VCC.n207 0.00675
R2233 VCC.n654 VCC.n653 0.00675
R2234 VCC.n237 VCC.n234 0.00675
R2235 VCC.n209 VCC.n208 0.00675
R2236 VCC.n655 VCC.n142 0.00675
R2237 VCC.n643 VCC.n154 0.00675
R2238 VCC.n236 VCC.n235 0.00675
R2239 VCC.n639 VCC.n158 0.00675
R2240 VCC.n784 VCC.n783 0.00585714
R2241 VCC.n808 VCC.n807 0.00585714
R2242 VCC.n883 VCC.n869 0.00585714
R2243 VCC.n907 VCC.n906 0.00585714
R2244 VCC.n896 VCC.n769 0.00585714
R2245 VCC.n403 VCC.n392 0.00585714
R2246 VCC.n400 VCC.n392 0.00585714
R2247 VCC.n427 VCC.n371 0.00585714
R2248 VCC.n462 VCC.n349 0.00585714
R2249 VCC.n506 VCC.n505 0.00585714
R2250 VCC.n445 VCC.n347 0.00585714
R2251 VCC.n482 VCC.n330 0.00585714
R2252 VCC.n524 VCC.n317 0.00585714
R2253 VCC.n561 VCC.n560 0.00585714
R2254 VCC.n582 VCC.n581 0.00585714
R2255 VCC.n594 VCC.n285 0.00585714
R2256 VCC.n276 VCC.n269 0.00585714
R2257 VCC.n611 VCC.n270 0.00585714
R2258 VCC.n320 VCC.n309 0.00585714
R2259 VCC.n555 VCC.n307 0.00585714
R2260 VCC.n583 VCC.n290 0.00585714
R2261 VCC.n25 VCC.n17 0.00585714
R2262 VCC.n17 VCC.n15 0.00585714
R2263 VCC.n55 VCC.n54 0.00585714
R2264 VCC.n92 VCC.n69 0.00585714
R2265 VCC.n679 VCC.n105 0.00585714
R2266 VCC.n67 VCC.n65 0.00585714
R2267 VCC.n691 VCC.n71 0.00585714
R2268 VCC.n199 VCC.n194 0.00585714
R2269 VCC.n186 VCC.n143 0.00585714
R2270 VCC.n644 VCC.n152 0.00585714
R2271 VCC.n238 VCC.n231 0.00585714
R2272 VCC.n249 VCC.n172 0.00585714
R2273 VCC.n174 VCC.n173 0.00585714
R2274 VCC.n659 VCC.n136 0.00585714
R2275 VCC.n145 VCC.n142 0.00585714
R2276 VCC.n643 VCC.n642 0.00585714
R2277 VCC.n844 VCC.n843 0.00496429
R2278 VCC.n843 VCC.n842 0.00496429
R2279 VCC.n917 VCC.n916 0.00496429
R2280 VCC.n907 VCC.n902 0.00496429
R2281 VCC.n761 VCC.n760 0.00496429
R2282 VCC.n749 VCC.n748 0.00496429
R2283 VCC.n738 VCC.n736 0.00496429
R2284 VCC.n400 VCC.n399 0.00496429
R2285 VCC.n390 VCC.n385 0.00496429
R2286 VCC.n417 VCC.n416 0.00496429
R2287 VCC.n441 VCC.n440 0.00496429
R2288 VCC.n513 VCC.n330 0.00496429
R2289 VCC.n516 VCC.n326 0.00496429
R2290 VCC.n531 VCC.n322 0.00496429
R2291 VCC.n536 VCC.n320 0.00496429
R2292 VCC.n288 VCC.n273 0.00496429
R2293 VCC.n607 VCC.n273 0.00496429
R2294 VCC.n610 VCC.n262 0.00496429
R2295 VCC.n31 VCC.n15 0.00496429
R2296 VCC.n729 VCC.n1 0.00496429
R2297 VCC.n726 VCC.n6 0.00496429
R2298 VCC.n713 VCC.n712 0.00496429
R2299 VCC.n124 VCC.n71 0.00496429
R2300 VCC.n127 VCC.n117 0.00496429
R2301 VCC.n666 VCC.n133 0.00496429
R2302 VCC.n662 VCC.n136 0.00496429
R2303 VCC.n638 VCC.n159 0.00496429
R2304 VCC.n635 VCC.n159 0.00496429
R2305 VCC.n632 VCC.n165 0.00496429
R2306 VCC.n442 VCC.n361 0.00486429
R2307 VCC.n452 VCC.n443 0.00486429
R2308 VCC.n451 VCC.n444 0.00486429
R2309 VCC.n479 VCC.n346 0.00486429
R2310 VCC.n557 VCC.n556 0.00486429
R2311 VCC.n575 VCC.n294 0.00486429
R2312 VCC.n577 VCC.n576 0.00486429
R2313 VCC.n584 VCC.n289 0.00486429
R2314 VCC.n898 VCC.n897 0.00486429
R2315 VCC.n766 VCC.n765 0.00486429
R2316 VCC.n764 VCC.n763 0.00486429
R2317 VCC.n762 VCC.n752 0.00486429
R2318 VCC.n711 VCC.n59 0.00486429
R2319 VCC.n710 VCC.n709 0.00486429
R2320 VCC.n701 VCC.n60 0.00486429
R2321 VCC.n700 VCC.n699 0.00486429
R2322 VCC.n656 VCC.n140 0.00486429
R2323 VCC.n649 VCC.n148 0.00486429
R2324 VCC.n648 VCC.n149 0.00486429
R2325 VCC.n641 VCC.n156 0.00486429
R2326 VCC.n786 VCC.n785 0.00407143
R2327 VCC.n825 VCC.n824 0.00407143
R2328 VCC.n830 VCC.n829 0.00407143
R2329 VCC.n849 VCC.n848 0.00407143
R2330 VCC.n894 VCC.n893 0.00407143
R2331 VCC.n449 VCC.n355 0.00407143
R2332 VCC.n506 VCC.n335 0.00407143
R2333 VCC.n450 VCC.n447 0.00407143
R2334 VCC.n705 VCC.n64 0.00407143
R2335 VCC.n680 VCC.n679 0.00407143
R2336 VCC.n704 VCC.n703 0.00407143
R2337 VCC.n443 VCC.n442 0.00318571
R2338 VCC.n444 VCC.n346 0.00318571
R2339 VCC.n556 VCC.n294 0.00318571
R2340 VCC.n577 VCC.n289 0.00318571
R2341 VCC.n897 VCC.n766 0.00318571
R2342 VCC.n763 VCC.n762 0.00318571
R2343 VCC.n711 VCC.n710 0.00318571
R2344 VCC.n701 VCC.n700 0.00318571
R2345 VCC.n148 VCC.n140 0.00318571
R2346 VCC.n156 VCC.n149 0.00318571
R2347 VCC.n790 VCC.n789 0.00317857
R2348 VCC.n889 VCC.n888 0.00317857
R2349 VCC.n848 VCC.n847 0.00317857
R2350 VCC.n834 VCC.n833 0.00317857
R2351 VCC.n916 VCC.n915 0.00317857
R2352 VCC.n902 VCC.n901 0.00317857
R2353 VCC.n754 VCC.n753 0.00317857
R2354 VCC.n748 VCC.n747 0.00317857
R2355 VCC.n736 VCC.n735 0.00317857
R2356 VCC.n404 VCC.n384 0.00317857
R2357 VCC.n415 VCC.n375 0.00317857
R2358 VCC.n415 VCC.n414 0.00317857
R2359 VCC.n364 VCC.n357 0.00317857
R2360 VCC.n455 VCC.n358 0.00317857
R2361 VCC.n461 VCC.n460 0.00317857
R2362 VCC.n512 VCC.n332 0.00317857
R2363 VCC.n512 VCC.n511 0.00317857
R2364 VCC.n517 VCC.n327 0.00317857
R2365 VCC.n391 VCC.n390 0.00317857
R2366 VCC.n416 VCC.n374 0.00317857
R2367 VCC.n454 VCC.n453 0.00317857
R2368 VCC.n513 VCC.n331 0.00317857
R2369 VCC.n516 VCC.n328 0.00317857
R2370 VCC.n530 VCC.n529 0.00317857
R2371 VCC.n535 VCC.n318 0.00317857
R2372 VCC.n580 VCC.n291 0.00317857
R2373 VCC.n589 VCC.n588 0.00317857
R2374 VCC.n606 VCC.n605 0.00317857
R2375 VCC.n612 VCC.n611 0.00317857
R2376 VCC.n612 VCC.n263 0.00317857
R2377 VCC.n531 VCC.n323 0.00317857
R2378 VCC.n537 VCC.n536 0.00317857
R2379 VCC.n579 VCC.n292 0.00317857
R2380 VCC.n607 VCC.n274 0.00317857
R2381 VCC.n613 VCC.n610 0.00317857
R2382 VCC.n730 VCC.n2 0.00317857
R2383 VCC.n725 VCC.n7 0.00317857
R2384 VCC.n725 VCC.n724 0.00317857
R2385 VCC.n82 VCC.n42 0.00317857
R2386 VCC.n707 VCC.n63 0.00317857
R2387 VCC.n91 VCC.n90 0.00317857
R2388 VCC.n123 VCC.n73 0.00317857
R2389 VCC.n123 VCC.n122 0.00317857
R2390 VCC.n128 VCC.n108 0.00317857
R2391 VCC.n729 VCC.n3 0.00317857
R2392 VCC.n726 VCC.n5 0.00317857
R2393 VCC.n708 VCC.n61 0.00317857
R2394 VCC.n124 VCC.n119 0.00317857
R2395 VCC.n127 VCC.n107 0.00317857
R2396 VCC.n197 VCC.n115 0.00317857
R2397 VCC.n661 VCC.n137 0.00317857
R2398 VCC.n646 VCC.n645 0.00317857
R2399 VCC.n233 VCC.n160 0.00317857
R2400 VCC.n636 VCC.n161 0.00317857
R2401 VCC.n173 VCC.n166 0.00317857
R2402 VCC.n631 VCC.n166 0.00317857
R2403 VCC.n196 VCC.n133 0.00317857
R2404 VCC.n662 VCC.n135 0.00317857
R2405 VCC.n647 VCC.n150 0.00317857
R2406 VCC.n635 VCC.n162 0.00317857
R2407 VCC.n632 VCC.n164 0.00317857
R2408 VCC.n771 VCC.n770 0.00228571
R2409 VCC.n791 VCC.n790 0.00228571
R2410 VCC.n885 VCC.n884 0.00228571
R2411 VCC.n869 VCC.n868 0.00228571
R2412 VCC.n424 VCC.n371 0.00228571
R2413 VCC.n550 VCC.n549 0.00228571
R2414 VCC.n561 VCC.n303 0.00228571
R2415 VCC.n573 VCC.n297 0.00228571
R2416 VCC.n594 VCC.n593 0.00228571
R2417 VCC.n574 VCC.n295 0.00228571
R2418 VCC.n54 VCC.n53 0.00228571
R2419 VCC.n211 VCC.n206 0.00228571
R2420 VCC.n207 VCC.n186 0.00228571
R2421 VCC.n652 VCC.n144 0.00228571
R2422 VCC.n238 VCC.n237 0.00228571
R2423 VCC.n651 VCC.n650 0.00228571
R2424 VCC.n389 VCC.n388 0.00217857
R2425 VCC.n418 VCC.n373 0.00217857
R2426 VCC.n514 VCC.n329 0.00217857
R2427 VCC.n515 VCC.n325 0.00217857
R2428 VCC.n532 VCC.n321 0.00217857
R2429 VCC.n533 VCC.n308 0.00217857
R2430 VCC.n608 VCC.n272 0.00217857
R2431 VCC.n609 VCC.n261 0.00217857
R2432 VCC.n918 VCC.n910 0.00217857
R2433 VCC.n909 VCC.n908 0.00217857
R2434 VCC.n750 VCC.n741 0.00217857
R2435 VCC.n740 VCC.n739 0.00217857
R2436 VCC.n728 VCC.n0 0.00217857
R2437 VCC.n727 VCC.n4 0.00217857
R2438 VCC.n125 VCC.n118 0.00217857
R2439 VCC.n126 VCC.n116 0.00217857
R2440 VCC.n665 VCC.n664 0.00217857
R2441 VCC.n663 VCC.n134 0.00217857
R2442 VCC.n634 VCC.n157 0.00217857
R2443 VCC.n633 VCC.n163 0.00217857
R2444 VCC.n772 VCC.n771 0.00139286
R2445 VCC.n809 VCC.n808 0.00139286
R2446 VCC.n890 VCC.n831 0.00139286
R2447 VCC.n835 VCC.n834 0.00139286
R2448 VCC.n892 VCC.n891 0.00139286
R2449 VCC.n422 VCC.n363 0.00139286
R2450 VCC.n477 VCC.n349 0.00139286
R2451 VCC.n604 VCC.n278 0.00139286
R2452 VCC.n617 VCC.n269 0.00139286
R2453 VCC.n715 VCC.n41 0.00139286
R2454 VCC.n697 VCC.n69 0.00139286
R2455 VCC.n248 VCC.n176 0.00139286
R2456 VCC.n254 VCC.n172 0.00139286
R2457 D0_BUF.n15 D0_BUF.n0 400.238
R2458 D0_BUF.n3 D0_BUF.n2 292.5
R2459 D0_BUF.n17 D0_BUF.n16 153.333
R2460 D0_BUF D0_BUF.n17 105.805
R2461 D0_BUF.n0 D0_BUF.t3 83.8685
R2462 D0_BUF.n16 D0_BUF.t2 80.9765
R2463 D0_BUF.n16 D0_BUF.t4 57.8405
R2464 D0_BUF.n0 D0_BUF.t5 54.9485
R2465 D0_BUF.n5 D0_BUF.t1 47.274
R2466 D0_BUF.n2 D0_BUF.t0 27.6955
R2467 D0_BUF.n17 D0_BUF.n15 23.9595
R2468 D0_BUF.n11 D0_BUF.n3 13.177
R2469 D0_BUF.n8 D0_BUF.n3 13.177
R2470 D0_BUF.n11 D0_BUF.n10 9.3005
R2471 D0_BUF.n9 D0_BUF.n8 9.3005
R2472 D0_BUF.n6 D0_BUF.n5 9.3005
R2473 D0_BUF.n7 D0_BUF.n4 9.3005
R2474 D0_BUF.n12 D0_BUF.n1 9.3005
R2475 D0_BUF.n14 D0_BUF.n13 9.3005
R2476 D0_BUF.n13 D0_BUF.n2 9.02061
R2477 D0_BUF.n6 D0_BUF.n2 9.0206
R2478 D0_BUF.n13 D0_BUF.n12 6.02403
R2479 D0_BUF.n7 D0_BUF.n6 6.02403
R2480 D0_BUF.n15 D0_BUF 5.08342
R2481 D0_BUF D0_BUF.n14 2.37139
R2482 D0_BUF.n12 D0_BUF.n11 0.376971
R2483 D0_BUF.n8 D0_BUF.n7 0.376971
R2484 D0_BUF.n10 D0_BUF.n9 0.190717
R2485 D0_BUF.n14 D0_BUF.n1 0.0439783
R2486 D0_BUF.n5 D0_BUF.n4 0.0439783
R2487 D0_BUF.n10 D0_BUF.n1 0.00321739
R2488 D0_BUF.n9 D0_BUF.n4 0.00321739
R2489 VREFL.n1 VREFL.t1 99.7169
R2490 VREFL.n0 VREFL.t0 44.9543
R2491 VREFL.n0 VREFL.t2 37.5373
R2492 VREFL.n1 VREFL.n0 2.88557
R2493 VREFL VREFL.n1 1.84958
R2494 D1.n1 D1.n0 127.099
R2495 D1.n0 D1.t0 77.6025
R2496 D1.n0 D1.t1 61.2145
R2497 D1.n1 D1 0.0485769
R2498 D1 D1.n1 0.0365577
R2499 VOUT.n0 VOUT.t1 46.8495
R2500 VOUT.n0 VOUT.t3 46.5654
R2501 VOUT.n5 VOUT.t0 34.887
R2502 VOUT.n10 VOUT.t2 27.6955
R2503 VOUT.n4 VOUT.n3 13.362
R2504 VOUT.n2 VOUT.n1 9.3005
R2505 VOUT.n7 VOUT.n6 9.3005
R2506 VOUT.n9 VOUT.n8 9.3005
R2507 VOUT.n12 VOUT.n11 9.3005
R2508 VOUT.n11 VOUT.n10 9.02061
R2509 VOUT.n5 VOUT.n4 4.55875
R2510 VOUT.n0 VOUT 3.09322
R2511 VOUT VOUT.n12 0.815717
R2512 VOUT.n2 VOUT.n0 0.613
R2513 VOUT.n12 VOUT.n9 0.0439783
R2514 VOUT.n7 VOUT.n5 0.0439783
R2515 VOUT.n5 VOUT.n2 0.014087
R2516 VOUT.n9 VOUT.n7 0.00321739
R2517 D2_BUF.n2 D2_BUF.n1 173.293
R2518 D2_BUF.n1 D2_BUF.t2 84.3505
R2519 D2_BUF.n1 D2_BUF.t3 53.5025
R2520 D2_BUF.n0 D2_BUF.t1 46.9077
R2521 D2_BUF.n0 D2_BUF.t0 35.0239
R2522 D2_BUF D2_BUF.n2 3.75226
R2523 D2_BUF.n2 D2_BUF.n0 0.204238
R2524 D1_BUF.n2 D1_BUF.n1 169.566
R2525 D1_BUF.n1 D1_BUF.t2 84.8325
R2526 D1_BUF.n1 D1_BUF.t3 53.0205
R2527 D1_BUF.n0 D1_BUF.t1 46.9158
R2528 D1_BUF.n0 D1_BUF.t0 35.0302
R2529 D1_BUF.n3 D1_BUF.n2 3.65455
R2530 D1_BUF D1_BUF.n3 2.60341
R2531 D1_BUF.n2 D1_BUF.n0 0.199588
R2532 D1_BUF.n3 D1_BUF 0.0389615
R2533 D2 D2.n0 125.046
R2534 D2.n0 D2.t0 77.1205
R2535 D2.n0 D2.t1 61.6965
R2536 VREFH VREFH.t0 98.071
C330 switch_n_3v3_1.D3 VSS 0.107f
C331 switch_n_3v3_1.D7 VSS 0.259f
C332 switch_n_3v3_1.D6 VSS 0.11f
C333 switch_n_3v3_1.D5 VSS 0.108f
C334 switch_n_3v3_1.D4 VSS 0.108f
C335 2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS 0.667f 
C336 2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS 1.53f 
C337 D1_BUF VSS 1.17f
C338 2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS 1.13f 
C339 D0_BUF VSS 2.53f
C340 a_1438_406# VSS 1.22f 
C341 2_bit_dac_0[0].switch2n_3v3_0.R_L VSS 0.676f 
C342 2_bit_dac_0[0].switch2n_3v3_0.R_H VSS 0.519f 
C343 VREFH VSS 0.29f
C344 2_bit_dac_0[0].switch2n_3v3_0.VREFH VSS 0.544f 
C345 2_bit_dac_0[0].VOUT VSS 1.32f 
C346 VOUT VSS 0.406f
C347 2_bit_dac_0[1].VOUT VSS 1.4f 
C348 2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS 0.905f 
C349 VREFL VSS 1.15f
C350 2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS 1.11f 
C351 D2_BUF VSS 1.15f
C352 switch_n_3v3_1.DX_ VSS 1.15f 
C353 D2 VSS 0.6f
C354 2_bit_dac_0[0].D1 VSS 1.63f 
C355 2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS 1.08f 
C356 D1 VSS 0.48f
C357 2_bit_dac_0[0].D0 VSS 3.37f 
C358 a_1438_1634# VSS 1.18f 
C359 D0 VSS 0.729f
C360 2_bit_dac_0[1].switch2n_3v3_0.R_L VSS 0.68f 
C361 2_bit_dac_0[1].switch2n_3v3_0.R_H VSS 0.521f 
C362 2_bit_dac_0[1].VREFH VSS 1.5f 
C363 2_bit_dac_0[1].switch2n_3v3_0.VREFH VSS 0.714f 
C364 VCC VSS 20.2f
.ends

X1 D0 VREFL D0_BUF VREFH D1 D1_BUF D2 D2_BUF VOUT VSS VCC x3_bit_dac


.param mc_mm_switch=0
.param mc_pr_switch=0
.lib "/foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice.tt.red" tt

*.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt.spice
*.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
*.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
*.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

V1 VSS 0 dc 0
V2 VCC 0 dc 3.3

V3 VREFL 0 dc 0
V4 VREFH 0 dc 3.3

V5  D0 0 PULSE(0 1.8 4n 1p 1p 4n 8n)
V6  D1 0 PULSE(0 1.8 8n 1p 1p 8n 16n)
V7  D2 0 PULSE(0 1.8 16n 1p 1p 16n 32n)



.tran 0.1n 128n uic


.control
run

set xbrushwidth=3
set hcopydevtype = svg

plot D0 D1 D2 VOUT

hardcopy 3_bit_dac_RCX.svg D0 D1 D2 VOUT

.endc
.end
