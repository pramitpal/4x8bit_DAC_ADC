* NGSPICE file created from Mux.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_g5v0d10v5_AWMFT3 a_n108_n84# w_n144_n146# a_50_n84# a_n50_n110#
X0 a_50_n84# a_n50_n110# a_n108_n84# w_n144_n146# sky130_fd_pr__pfet_g5v0d10v5 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.5
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_NQZZCX a_50_n42# a_n50_n68# a_n108_n42# VSUBS
X0 a_50_n42# a_n50_n68# a_n108_n42# VSUBS sky130_fd_pr__nfet_g5v0d10v5 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.5
.ends

.subckt Mux VCC VSS OUT SEL A B
Xsky130_fd_pr__pfet_g5v0d10v5_AWMFT3_0 VCC VCC a_8221_5082# SEL sky130_fd_pr__pfet_g5v0d10v5_AWMFT3
Xsky130_fd_pr__pfet_g5v0d10v5_AWMFT3_2 B VCC OUT SEL sky130_fd_pr__pfet_g5v0d10v5_AWMFT3
Xsky130_fd_pr__pfet_g5v0d10v5_AWMFT3_3 A VCC OUT a_8221_5082# sky130_fd_pr__pfet_g5v0d10v5_AWMFT3
Xsky130_fd_pr__nfet_g5v0d10v5_NQZZCX_0 OUT a_8221_5082# B VSS sky130_fd_pr__nfet_g5v0d10v5_NQZZCX
Xsky130_fd_pr__nfet_g5v0d10v5_NQZZCX_1 a_8221_5082# SEL VSS VSS sky130_fd_pr__nfet_g5v0d10v5_NQZZCX
Xsky130_fd_pr__nfet_g5v0d10v5_NQZZCX_2 OUT SEL A VSS sky130_fd_pr__nfet_g5v0d10v5_NQZZCX
.ends

