* NGSPICE file created from 4x8bit_tx_buffer.ext - technology: sky130A

.subckt switch_n_3v3 VREFH DX_BUF m2_n6802_n991# m2_n6562_n991# D7 D6 D5 D4 DX D3
+ D2 m2_n6722_n991# m2_n6482_n991# m2_n6882_n991# VCC VSS VOUT m2_n6642_n991# VREFL
X0 VOUT DX_BUF VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1 DX_ DX VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2 DX_BUF DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X3 VOUT DX_BUF VREFL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X4 DX_ DX VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5 VREFL DX_ VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6 DX_BUF DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7 VREFH DX_ VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt switch_n_3v3_v2 VREFH DX_BUF DX VCC VSS VOUT VREFL
X0 VOUT DX_BUF VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1 DX_ DX VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2 DX_BUF DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X3 VOUT DX_BUF VREFL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X4 DX_ DX VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5 VREFL DX_ VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6 DX_BUF DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7 VREFH DX_ VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt switch2n_3v3 VOUTL DX_BUF VOUTH DX VCC VSS a_n7536_n590# VREFL
X0 VOUTH a_n6524_n498# VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1 VREFH DX_BUF VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X2 VREFH R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X3 DX_BUF a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4 VREFL DX_BUF VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X5 VREFH a_n7536_n590# VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X6 a_n6524_n498# DX VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7 VOUTL a_n6524_n498# VREFL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X8 VOUTH a_n6524_n498# R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9 R_H DX_BUF VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X10 R_H R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X11 R_L VREFL VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X12 R_L DX_BUF VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X13 DX_BUF a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X14 a_n6524_n498# DX VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X15 VOUTL a_n6524_n498# R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
.ends

.subckt x2_bit_dac VREFH D1_BUF D1 D0 VCC D0_BUF VOUT VREFL VSS
Xswitch_n_3v3_v2_0 switch2n_3v3_0/VOUTH D1_BUF D1 VCC VSS VOUT switch2n_3v3_0/VOUTL
+ switch_n_3v3_v2
Xswitch2n_3v3_0 switch2n_3v3_0/VOUTL D0_BUF switch2n_3v3_0/VOUTH D0 VCC VSS VREFH
+ VREFL switch2n_3v3
.ends

.subckt x3_bit_dac VREFH D1_BUF switch_n_3v3_1/D6 switch_n_3v3_1/D7 switch_n_3v3_1/D5
+ switch_n_3v3_1/D4 switch_n_3v3_1/D3 D2_BUF D2 D1 D0 D0_BUF VCC VOUT VREFL VSS
X2_bit_dac_0[0] VREFH D1_BUF 2_bit_dac_0[0]/D1 2_bit_dac_0[0]/D0 VCC D0_BUF 2_bit_dac_0[0]/VOUT
+ 2_bit_dac_0[1]/VREFH VSS x2_bit_dac
X2_bit_dac_0[1] 2_bit_dac_0[1]/VREFH 2_bit_dac_0[0]/D1 D1 D0 VCC 2_bit_dac_0[0]/D0
+ 2_bit_dac_0[1]/VOUT VREFL VSS x2_bit_dac
Xswitch_n_3v3_1 2_bit_dac_0[0]/VOUT D2_BUF switch_n_3v3_1/D3 switch_n_3v3_1/D6 switch_n_3v3_1/D7
+ switch_n_3v3_1/D6 switch_n_3v3_1/D5 switch_n_3v3_1/D4 D2 switch_n_3v3_1/D3 D2 switch_n_3v3_1/D4
+ switch_n_3v3_1/D7 D2_BUF VCC VSS VOUT switch_n_3v3_1/D5 2_bit_dac_0[1]/VOUT switch_n_3v3
.ends

.subckt x4_bit_dac VREFH D1_BUF D2_BUF D3 D2 switch_n_3v3_0/D7 D1 switch_n_3v3_0/D6
+ D0 switch_n_3v3_0/D5 switch_n_3v3_0/D4 D3_BUF D0_BUF VCC VOUT VREFL VSS
X3_bit_dac_0[0] VREFH D1_BUF switch_n_3v3_0/D6 switch_n_3v3_0/D7 switch_n_3v3_0/D5
+ switch_n_3v3_0/D4 D3_BUF D2_BUF switch_n_3v3_0/D2 3_bit_dac_0[0]/D1 3_bit_dac_0[0]/D0
+ D0_BUF VCC 3_bit_dac_0[0]/VOUT 3_bit_dac_0[1]/VREFH VSS x3_bit_dac
X3_bit_dac_0[1] 3_bit_dac_0[1]/VREFH 3_bit_dac_0[0]/D1 switch_n_3v3_0/D6 switch_n_3v3_0/D7
+ switch_n_3v3_0/D5 switch_n_3v3_0/D4 D3 switch_n_3v3_0/D2 D2 D1 D0 3_bit_dac_0[0]/D0
+ VCC 3_bit_dac_0[1]/VOUT VREFL VSS x3_bit_dac
Xswitch_n_3v3_0 3_bit_dac_0[0]/VOUT D3_BUF D3_BUF switch_n_3v3_0/D6 switch_n_3v3_0/D7
+ switch_n_3v3_0/D6 switch_n_3v3_0/D5 switch_n_3v3_0/D4 D3 D3 switch_n_3v3_0/D2 switch_n_3v3_0/D4
+ switch_n_3v3_0/D7 switch_n_3v3_0/D2 VCC VSS VOUT switch_n_3v3_0/D5 3_bit_dac_0[1]/VOUT
+ switch_n_3v3
.ends

.subckt x5_bit_dac D4_BUF VREFH D1_BUF D2_BUF D4 D3 D2 switch_n_3v3_0/D7 D1 switch_n_3v3_0/D6
+ D0 switch_n_3v3_0/D5 D3_BUF D0_BUF VOUT VREFL VSS
X4_bit_dac_0[0] VREFH D1_BUF D2_BUF switch_n_3v3_0/D3 switch_n_3v3_0/D2 switch_n_3v3_0/D7
+ 4_bit_dac_0[0]/D1 switch_n_3v3_0/D6 4_bit_dac_0[0]/D0 switch_n_3v3_0/D5 D4_BUF D3_BUF
+ D0_BUF VCC 4_bit_dac_0[0]/VOUT 4_bit_dac_0[1]/VREFH VSS x4_bit_dac
X4_bit_dac_0[1] 4_bit_dac_0[1]/VREFH 4_bit_dac_0[0]/D1 switch_n_3v3_0/D2 D3 D2 switch_n_3v3_0/D7
+ D1 switch_n_3v3_0/D6 D0 switch_n_3v3_0/D5 D4 switch_n_3v3_0/D3 4_bit_dac_0[0]/D0
+ VCC 4_bit_dac_0[1]/VOUT VREFL VSS x4_bit_dac
Xswitch_n_3v3_0 4_bit_dac_0[0]/VOUT D4_BUF switch_n_3v3_0/D3 switch_n_3v3_0/D6 switch_n_3v3_0/D7
+ switch_n_3v3_0/D6 switch_n_3v3_0/D5 D4 D4 switch_n_3v3_0/D3 switch_n_3v3_0/D2 D4_BUF
+ switch_n_3v3_0/D7 switch_n_3v3_0/D2 VCC VSS VOUT switch_n_3v3_0/D5 4_bit_dac_0[1]/VOUT
+ switch_n_3v3
.ends

.subckt x6_bit_dac D4_BUF VREFH D1_BUF D5_BUF D2_BUF D5 D4 D3 D2 D1 D0 D3_BUF D0_BUF
+ VOUT VREFL VSS
Xswitch_n_3v3_0 5_bit_dac_0[0]/VOUT D5_BUF switch_n_3v3_0/D3 switch_n_3v3_0/D6 switch_n_3v3_0/D7
+ switch_n_3v3_0/D6 D5 switch_n_3v3_0/D4 D5 switch_n_3v3_0/D3 switch_n_3v3_0/D2 switch_n_3v3_0/D4
+ switch_n_3v3_0/D7 switch_n_3v3_0/D2 VCC VSS VOUT D5_BUF 5_bit_dac_0[1]/VOUT switch_n_3v3
X5_bit_dac_0[0] D4_BUF VREFH D1_BUF D2_BUF switch_n_3v3_0/D4 switch_n_3v3_0/D3 switch_n_3v3_0/D2
+ switch_n_3v3_0/D7 5_bit_dac_0[0]/D1 switch_n_3v3_0/D6 5_bit_dac_0[0]/D0 D5_BUF D3_BUF
+ D0_BUF 5_bit_dac_0[0]/VOUT 5_bit_dac_0[1]/VREFH VSS x5_bit_dac
X5_bit_dac_0[1] switch_n_3v3_0/D4 5_bit_dac_0[1]/VREFH 5_bit_dac_0[0]/D1 switch_n_3v3_0/D2
+ D4 D3 D2 switch_n_3v3_0/D7 D1 switch_n_3v3_0/D6 D0 D5 switch_n_3v3_0/D3 5_bit_dac_0[0]/D0
+ 5_bit_dac_0[1]/VOUT VREFL VSS x5_bit_dac
.ends

.subckt x7_bit_dac D4_BUF VREFH D1_BUF D5_BUF D2_BUF D6 D5 D4 D3 D2 D1 D0 D6_BUF D3_BUF
+ D0_BUF VCC VOUT VREFL VSS
X6_bit_dac_0[0] D4_BUF VREFH D1_BUF D5_BUF D2_BUF switch_n_3v3_1/D5 switch_n_3v3_1/D4
+ switch_n_3v3_1/D3 switch_n_3v3_1/D2 6_bit_dac_0[0]/D1 6_bit_dac_0[0]/D0 D3_BUF D0_BUF
+ 6_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/VREFH VSS x6_bit_dac
X6_bit_dac_0[1] switch_n_3v3_1/D4 6_bit_dac_0[1]/VREFH 6_bit_dac_0[0]/D1 switch_n_3v3_1/D5
+ switch_n_3v3_1/D2 D5 D4 D3 D2 D1 D0 switch_n_3v3_1/D3 6_bit_dac_0[0]/D0 6_bit_dac_0[1]/VOUT
+ VREFL VSS x6_bit_dac
Xswitch_n_3v3_1 6_bit_dac_0[0]/VOUT D6_BUF switch_n_3v3_1/D3 D6_BUF switch_n_3v3_1/D7
+ D6 switch_n_3v3_1/D5 switch_n_3v3_1/D4 D6 switch_n_3v3_1/D3 switch_n_3v3_1/D2 switch_n_3v3_1/D4
+ switch_n_3v3_1/D7 switch_n_3v3_1/D2 VCC VSS VOUT switch_n_3v3_1/D5 6_bit_dac_0[1]/VOUT
+ switch_n_3v3
.ends

.subckt x8_bit_dac VREFH D7 D6 D5 D4 D3 D2 D1 D0 VOUT VREFL VSS VCC
X7_bit_dac_0[0] D4_BUF VREFH D1_BUF D5_BUF D2_BUF switch_n_3v3_1/D6 switch_n_3v3_1/D5
+ switch_n_3v3_1/D4 switch_n_3v3_1/D3 switch_n_3v3_1/D2 7_bit_dac_0[0]/D1 7_bit_dac_0[0]/D0
+ D6_BUF D3_BUF D0_BUF VCC 7_bit_dac_0[0]/VOUT 7_bit_dac_0[1]/VREFH VSS x7_bit_dac
X7_bit_dac_0[1] switch_n_3v3_1/D4 7_bit_dac_0[1]/VREFH 7_bit_dac_0[0]/D1 switch_n_3v3_1/D5
+ switch_n_3v3_1/D2 D6 D5 D4 D3 D2 D1 D0 switch_n_3v3_1/D6 switch_n_3v3_1/D3 7_bit_dac_0[0]/D0
+ VCC 7_bit_dac_0[1]/VOUT VREFL VSS x7_bit_dac
Xswitch_n_3v3_1 7_bit_dac_0[0]/VOUT D7_BUF switch_n_3v3_1/D3 switch_n_3v3_1/D6 D7
+ switch_n_3v3_1/D6 switch_n_3v3_1/D5 switch_n_3v3_1/D4 D7 switch_n_3v3_1/D3 switch_n_3v3_1/D2
+ switch_n_3v3_1/D4 D7_BUF switch_n_3v3_1/D2 VCC VSS VOUT switch_n_3v3_1/D5 7_bit_dac_0[1]/VOUT
+ switch_n_3v3
.ends

.subckt level_tx_1bit VCCL VIN DVSS VCC VOUT
X0 DVSS a_n1600_540# a_n1428_490# DVSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X1 VOUT a_n1810_540# DVSS DVSS sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X2 a_n1600_540# a_n1810_540# VCCL VCCL sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X3 VCC a_n1428_490# VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X4 a_n1428_490# VOUT VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X5 a_n1810_540# VIN VCCL VCCL sky130_fd_pr__pfet_01v8 ad=0.244 pd=2.26 as=0.244 ps=2.26 w=0.84 l=0.15
X6 a_n1600_540# a_n1810_540# DVSS DVSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X7 a_n1810_540# VIN DVSS DVSS sky130_fd_pr__nfet_01v8 ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
.ends

.subckt level_tx_8bit VIN7 VIN6 VIN5 VIN4 VCCL VIN3 VIN2 VIN1 VIN0 VOUT7 VOUT6 VOUT5
+ VOUT4 VOUT3 VOUT2 VCC VOUT1 VOUT0 DVSS
Xlevel_tx_1bit_0[0] VCCL VIN0 DVSS VCC VOUT0 level_tx_1bit
Xlevel_tx_1bit_0[1] VCCL VIN1 DVSS VCC VOUT1 level_tx_1bit
Xlevel_tx_1bit_0[2] VCCL VIN2 DVSS VCC VOUT2 level_tx_1bit
Xlevel_tx_1bit_0[3] VCCL VIN3 DVSS VCC VOUT3 level_tx_1bit
Xlevel_tx_1bit_0[4] VCCL VIN4 DVSS VCC VOUT4 level_tx_1bit
Xlevel_tx_1bit_0[5] VCCL VIN5 DVSS VCC VOUT5 level_tx_1bit
Xlevel_tx_1bit_0[6] VCCL VIN6 DVSS VCC VOUT6 level_tx_1bit
Xlevel_tx_1bit_0[7] VCCL VIN7 DVSS VCC VOUT7 level_tx_1bit
.ends

.subckt opamp OUT VIN VDD GND
X0 a_1549_3140# a_550_1291# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X1 OUT a_2027_304# GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.5
X2 GND a_2027_304# OUT GND sky130_fd_pr__nfet_g5v0d10v5 ad=1.74 pd=12.6 as=0.87 ps=6.29 w=6 l=0.5
X3 a_925_2276# a_925_2276# GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X4 a_1095_1321# OUT a_937_1321# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X5 GND a_2027_304# OUT GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=0.87 ps=6.29 w=6 l=0.5
X6 a_925_2276# a_550_1291# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X7 GND a_925_2276# a_1392_2207# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
R0 a_550_1291# GND sky130_fd_pr__res_generic_po w=0.33 l=65.2
X8 a_937_1321# a_n804_1718# a_1473_304# w_1403_231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X9 a_1708_2207# VIN a_1549_3140# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
X10 VDD a_2388_2094# OUT VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X11 a_1549_3140# OUT a_1392_2207# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X12 a_1253_1321# VIN a_1095_1321# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X13 a_1095_1321# a_925_2276# GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.5
X14 OUT a_2027_304# GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.29 as=1.74 ps=12.6 w=6 l=0.5
X15 a_2027_304# a_n804_1718# a_1253_1321# w_1403_231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X16 VDD a_2168_2788# a_2168_2788# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X17 OUT a_2388_2094# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.3 as=1.45 ps=10.3 w=10 l=0.5
X18 a_1253_1321# a_550_1291# VDD w_1403_231# sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
R1 VDD a_n804_1718# sky130_fd_pr__res_generic_po w=0.33 l=38.5
X19 VDD a_550_1291# a_937_1321# w_1403_231# sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X20 VDD a_550_1291# a_550_1291# VDD sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=4.29 as=1.16 ps=8.58 w=4 l=0.5
X21 OUT a_2388_2094# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.3 as=2.9 ps=20.6 w=10 l=0.5
X22 VDD a_2388_2094# OUT VDD sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.6 as=1.45 ps=10.3 w=10 l=0.5
X23 a_1708_2207# a_925_2276# GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X24 GND a_1473_304# a_1473_304# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X25 a_2168_2788# a_n804_1718# a_1392_2207# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X26 a_1708_2207# a_n804_1718# a_2388_2094# GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
R2 a_n804_1718# GND sky130_fd_pr__res_generic_po w=0.33 l=23.6
X27 a_2027_304# a_1473_304# GND GND sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X28 a_2388_2094# a_2168_2788# VDD VDD sky130_fd_pr__pfet_g5v0d10v5 ad=1.16 pd=8.58 as=0.58 ps=4.29 w=4 l=0.5
.ends

.subckt x8_bit_dac_tx_buffer_v2 VREFH VCCD D7 VSSD D6 D5 D4 D3 D2 D1 D0 VDDA VREFL
+ VOUT 8_bit_dac_0/VCC VSSA
X8_bit_dac_0 VREFH 8_bit_dac_0/D7 8_bit_dac_0/D6 8_bit_dac_0/D5 8_bit_dac_0/D4 8_bit_dac_0/D3
+ 8_bit_dac_0/D2 8_bit_dac_0/D1 8_bit_dac_0/D0 opamp_0/VIN VREFL VSSA 8_bit_dac_0/VCC
+ x8_bit_dac
Xlevel_tx_8bit_0 D7 D6 D5 D4 VCCD D3 D2 D1 D0 8_bit_dac_0/D7 8_bit_dac_0/D6 8_bit_dac_0/D5
+ 8_bit_dac_0/D4 8_bit_dac_0/D3 8_bit_dac_0/D2 8_bit_dac_0/VCC 8_bit_dac_0/D1 8_bit_dac_0/D0
+ VSSD level_tx_8bit
Xopamp_0 VOUT opamp_0/VIN VDDA VSSA opamp
.ends

.subckt x2x8bit_tx_buffer D11 D10 D00 VREFH VCCD VSSD VOUT1 D07 D17 VOUT0 D06 D16
+ D05 VDDA D15 D04 D14 D03 VREFL D13 D02 D12 D01 VSSA
X8_bit_dac_tx_buffer_v2_0[0] VREFH VCCD D07 VSSD D06 D05 D04 D03 D02 D01 D00 VDDA
+ VREFL VOUT0 VDDA VSSA x8_bit_dac_tx_buffer_v2
X8_bit_dac_tx_buffer_v2_0[1] VREFH VCCD D17 VSSD D16 D15 D14 D13 D12 D11 D10 VDDA
+ VREFL VOUT1 VDDA VSSA x8_bit_dac_tx_buffer_v2
.ends

.subckt x4x8bit_tx_buffer D00 D01 D02 D03 D04 D05 D06 D07 D10 D11 D12 D13 D14 D15
+ D16 D17 D20 D21 D22 D23 D24 D25 D26 D27 D30 D31 D32 D33 D34 D35 D36 D37 VCCD VDDA
+ VOUT0 VOUT1 VOUT2 VOUT3 VREFH VREFL VSSA VSSD
X2x8bit_tx_buffer_0[0] D11 D10 D00 VREFH VCCD VSSD VOUT1 D07 D17 VOUT0 D06 D16 D05
+ VDDA D15 D04 D14 D03 VREFL D13 D02 D12 D01 VSSA x2x8bit_tx_buffer
X2x8bit_tx_buffer_0[1] D31 D30 D20 VREFH VCCD VSSD VOUT3 D27 D37 VOUT2 D26 D36 D25
+ VDDA D35 D24 D34 D23 VREFL D33 D22 D32 D21 VSSA x2x8bit_tx_buffer
.ends

