magic
tech sky130A
magscale 1 2
timestamp 1687028152
<< isosubstrate >>
rect 946 78804 6730 80552
<< metal2 >>
rect 35 84716 44 84784
rect 112 84716 121 84784
rect 44 80346 112 84716
rect 277 81506 286 81574
rect 354 81506 363 81574
rect 35 80278 44 80346
rect 112 80278 121 80346
rect 44 78198 112 80278
rect 286 79940 354 81506
rect 642 80648 682 85090
rect 780 80738 820 85090
rect 916 80828 956 85090
rect 1050 80918 1090 85090
rect 1182 81010 1222 85090
rect 1314 81110 1354 85090
rect 1446 81208 1486 85090
rect 1580 81316 1620 85090
rect 6408 82750 6456 85090
rect 6262 82702 6456 82750
rect 6278 81952 6388 81992
rect 1580 81276 5948 81316
rect 1446 81168 5272 81208
rect 1314 81070 4588 81110
rect 1182 80970 3920 81010
rect 1050 80878 3224 80918
rect 916 80788 2544 80828
rect 780 80698 1860 80738
rect 642 80608 1200 80648
rect 146 79872 354 79940
rect 146 77496 214 79872
rect 1160 79850 1200 80608
rect 1160 79810 1300 79850
rect 1260 79612 1300 79810
rect 1820 79848 1860 80698
rect 2504 79848 2544 80788
rect 1820 79808 1980 79848
rect 2504 79808 2660 79848
rect 1807 79667 1877 79702
rect 1842 78722 1877 79667
rect 1940 79612 1980 79808
rect 2487 79667 2561 79702
rect 2526 78770 2561 79667
rect 2620 79612 2660 79808
rect 3184 79838 3224 80878
rect 3880 79862 3920 80970
rect 3184 79798 3340 79838
rect 3880 79822 4020 79862
rect 3167 79667 3237 79702
rect 3202 78858 3237 79667
rect 3300 79612 3340 79798
rect 3847 79667 3919 79702
rect 3202 78823 3819 78858
rect 2526 78735 3605 78770
rect 276 78687 1877 78722
rect 276 78500 331 78687
rect 3570 78433 3605 78735
rect 3784 78630 3819 78823
rect 3884 78714 3919 79667
rect 3980 79612 4020 79822
rect 4548 79856 4588 81070
rect 5232 79880 5272 81168
rect 5908 79884 5948 81276
rect 6336 80746 6388 81952
rect 6336 80694 7658 80746
rect 4548 79816 4700 79856
rect 5232 79840 5380 79880
rect 5908 79844 6060 79884
rect 4516 79667 4597 79702
rect 4562 78786 4597 79667
rect 4660 79612 4700 79816
rect 5207 79667 5275 79702
rect 5240 78866 5275 79667
rect 5340 79612 5380 79840
rect 5887 79667 5955 79702
rect 5240 78831 5401 78866
rect 4562 78751 5321 78786
rect 3884 78679 5243 78714
rect 3784 78595 5165 78630
rect 5124 78536 5165 78595
rect 5208 78561 5243 78679
rect 5286 78517 5321 78751
rect 5366 78537 5401 78831
rect 5920 78716 5955 79667
rect 6020 79612 6060 79844
rect 6567 79667 6655 79702
rect 5445 78681 5955 78716
rect 5445 78567 5480 78681
rect 6620 78632 6655 79667
rect 5524 78597 6655 78632
rect 5524 78528 5565 78597
rect 7606 78418 7658 80694
rect 380 0 435 301
<< via2 >>
rect 44 84716 112 84784
rect 286 81506 354 81574
rect 44 80278 112 80346
<< metal3 >>
rect 0 84784 7726 84902
rect 0 84716 44 84784
rect 112 84716 7726 84784
rect 0 84602 7726 84716
rect 0 81574 7726 81692
rect 0 81506 286 81574
rect 354 81506 7726 81574
rect 0 81392 7726 81506
rect 0 80346 7726 80362
rect 0 80278 44 80346
rect 112 80278 7726 80346
rect 0 80262 7726 80278
rect 0 79392 7726 79492
rect 0 78932 7726 79032
rect 80 77584 670 77724
use 8_bit_dac  8_bit_dac_0
timestamp 1687027365
transform 1 0 2 0 1 0
box -2 0 7724 78592
use level_tx_8bit  level_tx_8bit_0
timestamp 1687027365
transform 1 0 1160 0 1 78842
box 20 40 5460 1590
use opamp  opamp_0
timestamp 1687027365
transform 1 0 1622 0 1 82702
box 272 -1310 4740 2280
<< labels >>
rlabel metal3 476 80300 476 80300 1 VDDA
rlabel metal3 450 79430 450 79430 1 VSSD
rlabel metal3 440 78980 440 78980 1 VCCD
rlabel metal3 250 77660 250 77660 1 VSSA
rlabel metal2 1180 80450 1180 80450 1 D0
rlabel metal2 1840 80470 1840 80470 1 D1
rlabel metal2 2520 80480 2520 80480 1 D2
rlabel metal2 3200 80470 3200 80470 1 D3
rlabel metal2 3900 80470 3900 80470 1 D4
rlabel metal2 4570 80470 4570 80470 1 D5
rlabel metal2 5250 80470 5250 80470 1 D6
rlabel metal2 5930 80470 5930 80470 1 D7
rlabel metal2 7630 78540 7630 78540 1 VOUT
rlabel metal2 416 68 416 68 1 VREFH
rlabel metal2 6430 85040 6430 85040 1 VOUT_BUF
<< end >>
