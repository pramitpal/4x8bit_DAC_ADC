magic
tech sky130A
magscale 1 2
timestamp 1686247030
<< nwell >>
rect 677 3755 3685 3957
rect 697 2969 3685 3755
rect 1323 2691 3685 2969
rect 1323 2141 1832 2691
rect 1478 784 2021 1813
rect 2837 1707 3683 2691
rect 1403 231 2159 784
<< pwell >>
rect 841 2276 1109 2728
rect 2362 2516 2630 2520
rect 2085 2068 2630 2516
rect 2085 2064 2353 2068
rect 911 1295 1337 1747
rect 915 350 1183 1295
rect 2155 1263 2581 1715
rect 2893 617 3635 1504
rect 2312 252 3635 617
rect 2312 165 2738 252
rect -490 -4 1239 157
<< mvnmos >>
rect 925 2302 1025 2702
rect 2169 2090 2269 2490
rect 2446 2094 2546 2494
rect 995 1321 1095 1721
rect 1153 1321 1253 1721
rect 999 376 1099 1176
rect 2239 1289 2339 1689
rect 2397 1289 2497 1689
rect 2396 191 2496 591
rect 2554 191 2654 591
rect 2977 278 3077 1478
rect 3135 278 3235 1478
rect 3293 278 3393 1478
rect 3451 278 3551 1478
<< mvpmos >>
rect 825 3036 925 3836
rect 983 3036 1083 3836
rect 1449 3140 1549 3540
rect 1450 2207 1550 3007
rect 1608 2207 1708 3007
rect 2226 2788 2326 3588
rect 2384 2788 2484 3588
rect 2972 1811 3072 3811
rect 3130 1811 3230 3811
rect 3288 1811 3388 3811
rect 3446 1811 3546 3811
rect 1630 941 1730 1741
rect 1788 941 1888 1741
rect 1531 304 1631 704
rect 1927 304 2027 704
<< mvndiff >>
rect 867 2689 925 2702
rect 867 2655 879 2689
rect 913 2655 925 2689
rect 867 2621 925 2655
rect 867 2587 879 2621
rect 913 2587 925 2621
rect 867 2553 925 2587
rect 867 2519 879 2553
rect 913 2519 925 2553
rect 867 2485 925 2519
rect 867 2451 879 2485
rect 913 2451 925 2485
rect 867 2417 925 2451
rect 867 2383 879 2417
rect 913 2383 925 2417
rect 867 2349 925 2383
rect 867 2315 879 2349
rect 913 2315 925 2349
rect 867 2302 925 2315
rect 1025 2689 1083 2702
rect 1025 2655 1037 2689
rect 1071 2655 1083 2689
rect 1025 2621 1083 2655
rect 1025 2587 1037 2621
rect 1071 2587 1083 2621
rect 1025 2553 1083 2587
rect 1025 2519 1037 2553
rect 1071 2519 1083 2553
rect 1025 2485 1083 2519
rect 1025 2451 1037 2485
rect 1071 2451 1083 2485
rect 1025 2417 1083 2451
rect 1025 2383 1037 2417
rect 1071 2383 1083 2417
rect 1025 2349 1083 2383
rect 1025 2315 1037 2349
rect 1071 2315 1083 2349
rect 1025 2302 1083 2315
rect 2111 2477 2169 2490
rect 2111 2443 2123 2477
rect 2157 2443 2169 2477
rect 2111 2409 2169 2443
rect 2111 2375 2123 2409
rect 2157 2375 2169 2409
rect 2111 2341 2169 2375
rect 2111 2307 2123 2341
rect 2157 2307 2169 2341
rect 2111 2273 2169 2307
rect 2111 2239 2123 2273
rect 2157 2239 2169 2273
rect 2111 2205 2169 2239
rect 2111 2171 2123 2205
rect 2157 2171 2169 2205
rect 2111 2137 2169 2171
rect 2111 2103 2123 2137
rect 2157 2103 2169 2137
rect 2111 2090 2169 2103
rect 2269 2477 2327 2490
rect 2269 2443 2281 2477
rect 2315 2443 2327 2477
rect 2269 2409 2327 2443
rect 2269 2375 2281 2409
rect 2315 2375 2327 2409
rect 2269 2341 2327 2375
rect 2269 2307 2281 2341
rect 2315 2307 2327 2341
rect 2269 2273 2327 2307
rect 2269 2239 2281 2273
rect 2315 2239 2327 2273
rect 2269 2205 2327 2239
rect 2269 2171 2281 2205
rect 2315 2171 2327 2205
rect 2269 2137 2327 2171
rect 2269 2103 2281 2137
rect 2315 2103 2327 2137
rect 2269 2090 2327 2103
rect 2388 2481 2446 2494
rect 2388 2447 2400 2481
rect 2434 2447 2446 2481
rect 2388 2413 2446 2447
rect 2388 2379 2400 2413
rect 2434 2379 2446 2413
rect 2388 2345 2446 2379
rect 2388 2311 2400 2345
rect 2434 2311 2446 2345
rect 2388 2277 2446 2311
rect 2388 2243 2400 2277
rect 2434 2243 2446 2277
rect 2388 2209 2446 2243
rect 2388 2175 2400 2209
rect 2434 2175 2446 2209
rect 2388 2141 2446 2175
rect 2388 2107 2400 2141
rect 2434 2107 2446 2141
rect 2388 2094 2446 2107
rect 2546 2481 2604 2494
rect 2546 2447 2558 2481
rect 2592 2447 2604 2481
rect 2546 2413 2604 2447
rect 2546 2379 2558 2413
rect 2592 2379 2604 2413
rect 2546 2345 2604 2379
rect 2546 2311 2558 2345
rect 2592 2311 2604 2345
rect 2546 2277 2604 2311
rect 2546 2243 2558 2277
rect 2592 2243 2604 2277
rect 2546 2209 2604 2243
rect 2546 2175 2558 2209
rect 2592 2175 2604 2209
rect 2546 2141 2604 2175
rect 2546 2107 2558 2141
rect 2592 2107 2604 2141
rect 2546 2094 2604 2107
rect 937 1708 995 1721
rect 937 1674 949 1708
rect 983 1674 995 1708
rect 937 1640 995 1674
rect 937 1606 949 1640
rect 983 1606 995 1640
rect 937 1572 995 1606
rect 937 1538 949 1572
rect 983 1538 995 1572
rect 937 1504 995 1538
rect 937 1470 949 1504
rect 983 1470 995 1504
rect 937 1436 995 1470
rect 937 1402 949 1436
rect 983 1402 995 1436
rect 937 1368 995 1402
rect 937 1334 949 1368
rect 983 1334 995 1368
rect 937 1321 995 1334
rect 1095 1708 1153 1721
rect 1095 1674 1107 1708
rect 1141 1674 1153 1708
rect 1095 1640 1153 1674
rect 1095 1606 1107 1640
rect 1141 1606 1153 1640
rect 1095 1572 1153 1606
rect 1095 1538 1107 1572
rect 1141 1538 1153 1572
rect 1095 1504 1153 1538
rect 1095 1470 1107 1504
rect 1141 1470 1153 1504
rect 1095 1436 1153 1470
rect 1095 1402 1107 1436
rect 1141 1402 1153 1436
rect 1095 1368 1153 1402
rect 1095 1334 1107 1368
rect 1141 1334 1153 1368
rect 1095 1321 1153 1334
rect 1253 1708 1311 1721
rect 1253 1674 1265 1708
rect 1299 1674 1311 1708
rect 1253 1640 1311 1674
rect 1253 1606 1265 1640
rect 1299 1606 1311 1640
rect 1253 1572 1311 1606
rect 1253 1538 1265 1572
rect 1299 1538 1311 1572
rect 1253 1504 1311 1538
rect 1253 1470 1265 1504
rect 1299 1470 1311 1504
rect 1253 1436 1311 1470
rect 1253 1402 1265 1436
rect 1299 1402 1311 1436
rect 1253 1368 1311 1402
rect 1253 1334 1265 1368
rect 1299 1334 1311 1368
rect 1253 1321 1311 1334
rect 941 1133 999 1176
rect 941 1099 953 1133
rect 987 1099 999 1133
rect 941 1065 999 1099
rect 941 1031 953 1065
rect 987 1031 999 1065
rect 941 997 999 1031
rect 941 963 953 997
rect 987 963 999 997
rect 941 929 999 963
rect 941 895 953 929
rect 987 895 999 929
rect 941 861 999 895
rect 941 827 953 861
rect 987 827 999 861
rect 941 793 999 827
rect 941 759 953 793
rect 987 759 999 793
rect 941 725 999 759
rect 941 691 953 725
rect 987 691 999 725
rect 941 657 999 691
rect 941 623 953 657
rect 987 623 999 657
rect 941 589 999 623
rect 941 555 953 589
rect 987 555 999 589
rect 941 521 999 555
rect 941 487 953 521
rect 987 487 999 521
rect 941 453 999 487
rect 941 419 953 453
rect 987 419 999 453
rect 941 376 999 419
rect 1099 1133 1157 1176
rect 1099 1099 1111 1133
rect 1145 1099 1157 1133
rect 1099 1065 1157 1099
rect 1099 1031 1111 1065
rect 1145 1031 1157 1065
rect 1099 997 1157 1031
rect 1099 963 1111 997
rect 1145 963 1157 997
rect 1099 929 1157 963
rect 2181 1676 2239 1689
rect 2181 1642 2193 1676
rect 2227 1642 2239 1676
rect 2181 1608 2239 1642
rect 2181 1574 2193 1608
rect 2227 1574 2239 1608
rect 2181 1540 2239 1574
rect 2181 1506 2193 1540
rect 2227 1506 2239 1540
rect 2181 1472 2239 1506
rect 2181 1438 2193 1472
rect 2227 1438 2239 1472
rect 2181 1404 2239 1438
rect 2181 1370 2193 1404
rect 2227 1370 2239 1404
rect 2181 1336 2239 1370
rect 2181 1302 2193 1336
rect 2227 1302 2239 1336
rect 2181 1289 2239 1302
rect 2339 1676 2397 1689
rect 2339 1642 2351 1676
rect 2385 1642 2397 1676
rect 2339 1608 2397 1642
rect 2339 1574 2351 1608
rect 2385 1574 2397 1608
rect 2339 1540 2397 1574
rect 2339 1506 2351 1540
rect 2385 1506 2397 1540
rect 2339 1472 2397 1506
rect 2339 1438 2351 1472
rect 2385 1438 2397 1472
rect 2339 1404 2397 1438
rect 2339 1370 2351 1404
rect 2385 1370 2397 1404
rect 2339 1336 2397 1370
rect 2339 1302 2351 1336
rect 2385 1302 2397 1336
rect 2339 1289 2397 1302
rect 2497 1676 2555 1689
rect 2497 1642 2509 1676
rect 2543 1642 2555 1676
rect 2497 1608 2555 1642
rect 2497 1574 2509 1608
rect 2543 1574 2555 1608
rect 2497 1540 2555 1574
rect 2497 1506 2509 1540
rect 2543 1506 2555 1540
rect 2497 1472 2555 1506
rect 2497 1438 2509 1472
rect 2543 1438 2555 1472
rect 2497 1404 2555 1438
rect 2497 1370 2509 1404
rect 2543 1370 2555 1404
rect 2497 1336 2555 1370
rect 2497 1302 2509 1336
rect 2543 1302 2555 1336
rect 2497 1289 2555 1302
rect 2919 1439 2977 1478
rect 2919 1405 2931 1439
rect 2965 1405 2977 1439
rect 2919 1371 2977 1405
rect 2919 1337 2931 1371
rect 2965 1337 2977 1371
rect 2919 1303 2977 1337
rect 2919 1269 2931 1303
rect 2965 1269 2977 1303
rect 2919 1235 2977 1269
rect 2919 1201 2931 1235
rect 2965 1201 2977 1235
rect 2919 1167 2977 1201
rect 2919 1133 2931 1167
rect 2965 1133 2977 1167
rect 2919 1099 2977 1133
rect 2919 1065 2931 1099
rect 2965 1065 2977 1099
rect 2919 1031 2977 1065
rect 2919 997 2931 1031
rect 2965 997 2977 1031
rect 2919 963 2977 997
rect 1099 895 1111 929
rect 1145 895 1157 929
rect 2919 929 2931 963
rect 2965 929 2977 963
rect 1099 861 1157 895
rect 1099 827 1111 861
rect 1145 827 1157 861
rect 1099 793 1157 827
rect 1099 759 1111 793
rect 1145 759 1157 793
rect 1099 725 1157 759
rect 1099 691 1111 725
rect 1145 691 1157 725
rect 2919 895 2977 929
rect 2919 861 2931 895
rect 2965 861 2977 895
rect 2919 827 2977 861
rect 2919 793 2931 827
rect 2965 793 2977 827
rect 1099 657 1157 691
rect 1099 623 1111 657
rect 1145 623 1157 657
rect 1099 589 1157 623
rect 1099 555 1111 589
rect 1145 555 1157 589
rect 1099 521 1157 555
rect 1099 487 1111 521
rect 1145 487 1157 521
rect 1099 453 1157 487
rect 1099 419 1111 453
rect 1145 419 1157 453
rect 1099 376 1157 419
rect 2919 759 2977 793
rect 2919 725 2931 759
rect 2965 725 2977 759
rect 2919 691 2977 725
rect 2919 657 2931 691
rect 2965 657 2977 691
rect 2919 623 2977 657
rect 2338 578 2396 591
rect 2338 544 2350 578
rect 2384 544 2396 578
rect 2338 510 2396 544
rect 2338 476 2350 510
rect 2384 476 2396 510
rect 2338 442 2396 476
rect 2338 408 2350 442
rect 2384 408 2396 442
rect 2338 374 2396 408
rect 2338 340 2350 374
rect 2384 340 2396 374
rect 2338 306 2396 340
rect 2338 272 2350 306
rect 2384 272 2396 306
rect 2338 238 2396 272
rect 2338 204 2350 238
rect 2384 204 2396 238
rect 2338 191 2396 204
rect 2496 578 2554 591
rect 2496 544 2508 578
rect 2542 544 2554 578
rect 2496 510 2554 544
rect 2496 476 2508 510
rect 2542 476 2554 510
rect 2496 442 2554 476
rect 2496 408 2508 442
rect 2542 408 2554 442
rect 2496 374 2554 408
rect 2496 340 2508 374
rect 2542 340 2554 374
rect 2496 306 2554 340
rect 2496 272 2508 306
rect 2542 272 2554 306
rect 2496 238 2554 272
rect 2496 204 2508 238
rect 2542 204 2554 238
rect 2496 191 2554 204
rect 2654 578 2712 591
rect 2654 544 2666 578
rect 2700 544 2712 578
rect 2654 510 2712 544
rect 2654 476 2666 510
rect 2700 476 2712 510
rect 2654 442 2712 476
rect 2654 408 2666 442
rect 2700 408 2712 442
rect 2654 374 2712 408
rect 2654 340 2666 374
rect 2700 340 2712 374
rect 2654 306 2712 340
rect 2654 272 2666 306
rect 2700 272 2712 306
rect 2919 589 2931 623
rect 2965 589 2977 623
rect 2919 555 2977 589
rect 2919 521 2931 555
rect 2965 521 2977 555
rect 2919 487 2977 521
rect 2919 453 2931 487
rect 2965 453 2977 487
rect 2919 419 2977 453
rect 2919 385 2931 419
rect 2965 385 2977 419
rect 2919 351 2977 385
rect 2919 317 2931 351
rect 2965 317 2977 351
rect 2919 278 2977 317
rect 3077 1439 3135 1478
rect 3077 1405 3089 1439
rect 3123 1405 3135 1439
rect 3077 1371 3135 1405
rect 3077 1337 3089 1371
rect 3123 1337 3135 1371
rect 3077 1303 3135 1337
rect 3077 1269 3089 1303
rect 3123 1269 3135 1303
rect 3077 1235 3135 1269
rect 3077 1201 3089 1235
rect 3123 1201 3135 1235
rect 3077 1167 3135 1201
rect 3077 1133 3089 1167
rect 3123 1133 3135 1167
rect 3077 1099 3135 1133
rect 3077 1065 3089 1099
rect 3123 1065 3135 1099
rect 3077 1031 3135 1065
rect 3077 997 3089 1031
rect 3123 997 3135 1031
rect 3077 963 3135 997
rect 3077 929 3089 963
rect 3123 929 3135 963
rect 3077 895 3135 929
rect 3077 861 3089 895
rect 3123 861 3135 895
rect 3077 827 3135 861
rect 3077 793 3089 827
rect 3123 793 3135 827
rect 3077 759 3135 793
rect 3077 725 3089 759
rect 3123 725 3135 759
rect 3077 691 3135 725
rect 3077 657 3089 691
rect 3123 657 3135 691
rect 3077 623 3135 657
rect 3077 589 3089 623
rect 3123 589 3135 623
rect 3077 555 3135 589
rect 3077 521 3089 555
rect 3123 521 3135 555
rect 3077 487 3135 521
rect 3077 453 3089 487
rect 3123 453 3135 487
rect 3077 419 3135 453
rect 3077 385 3089 419
rect 3123 385 3135 419
rect 3077 351 3135 385
rect 3077 317 3089 351
rect 3123 317 3135 351
rect 3077 278 3135 317
rect 3235 1439 3293 1478
rect 3235 1405 3247 1439
rect 3281 1405 3293 1439
rect 3235 1371 3293 1405
rect 3235 1337 3247 1371
rect 3281 1337 3293 1371
rect 3235 1303 3293 1337
rect 3235 1269 3247 1303
rect 3281 1269 3293 1303
rect 3235 1235 3293 1269
rect 3235 1201 3247 1235
rect 3281 1201 3293 1235
rect 3235 1167 3293 1201
rect 3235 1133 3247 1167
rect 3281 1133 3293 1167
rect 3235 1099 3293 1133
rect 3235 1065 3247 1099
rect 3281 1065 3293 1099
rect 3235 1031 3293 1065
rect 3235 997 3247 1031
rect 3281 997 3293 1031
rect 3235 963 3293 997
rect 3235 929 3247 963
rect 3281 929 3293 963
rect 3235 895 3293 929
rect 3235 861 3247 895
rect 3281 861 3293 895
rect 3235 827 3293 861
rect 3235 793 3247 827
rect 3281 793 3293 827
rect 3235 759 3293 793
rect 3235 725 3247 759
rect 3281 725 3293 759
rect 3235 691 3293 725
rect 3235 657 3247 691
rect 3281 657 3293 691
rect 3235 623 3293 657
rect 3235 589 3247 623
rect 3281 589 3293 623
rect 3235 555 3293 589
rect 3235 521 3247 555
rect 3281 521 3293 555
rect 3235 487 3293 521
rect 3235 453 3247 487
rect 3281 453 3293 487
rect 3235 419 3293 453
rect 3235 385 3247 419
rect 3281 385 3293 419
rect 3235 351 3293 385
rect 3235 317 3247 351
rect 3281 317 3293 351
rect 3235 278 3293 317
rect 3393 1439 3451 1478
rect 3393 1405 3405 1439
rect 3439 1405 3451 1439
rect 3393 1371 3451 1405
rect 3393 1337 3405 1371
rect 3439 1337 3451 1371
rect 3393 1303 3451 1337
rect 3393 1269 3405 1303
rect 3439 1269 3451 1303
rect 3393 1235 3451 1269
rect 3393 1201 3405 1235
rect 3439 1201 3451 1235
rect 3393 1167 3451 1201
rect 3393 1133 3405 1167
rect 3439 1133 3451 1167
rect 3393 1099 3451 1133
rect 3393 1065 3405 1099
rect 3439 1065 3451 1099
rect 3393 1031 3451 1065
rect 3393 997 3405 1031
rect 3439 997 3451 1031
rect 3393 963 3451 997
rect 3393 929 3405 963
rect 3439 929 3451 963
rect 3393 895 3451 929
rect 3393 861 3405 895
rect 3439 861 3451 895
rect 3393 827 3451 861
rect 3393 793 3405 827
rect 3439 793 3451 827
rect 3393 759 3451 793
rect 3393 725 3405 759
rect 3439 725 3451 759
rect 3393 691 3451 725
rect 3393 657 3405 691
rect 3439 657 3451 691
rect 3393 623 3451 657
rect 3393 589 3405 623
rect 3439 589 3451 623
rect 3393 555 3451 589
rect 3393 521 3405 555
rect 3439 521 3451 555
rect 3393 487 3451 521
rect 3393 453 3405 487
rect 3439 453 3451 487
rect 3393 419 3451 453
rect 3393 385 3405 419
rect 3439 385 3451 419
rect 3393 351 3451 385
rect 3393 317 3405 351
rect 3439 317 3451 351
rect 3393 278 3451 317
rect 3551 1439 3609 1478
rect 3551 1405 3563 1439
rect 3597 1405 3609 1439
rect 3551 1371 3609 1405
rect 3551 1337 3563 1371
rect 3597 1337 3609 1371
rect 3551 1303 3609 1337
rect 3551 1269 3563 1303
rect 3597 1269 3609 1303
rect 3551 1235 3609 1269
rect 3551 1201 3563 1235
rect 3597 1201 3609 1235
rect 3551 1167 3609 1201
rect 3551 1133 3563 1167
rect 3597 1133 3609 1167
rect 3551 1099 3609 1133
rect 3551 1065 3563 1099
rect 3597 1065 3609 1099
rect 3551 1031 3609 1065
rect 3551 997 3563 1031
rect 3597 997 3609 1031
rect 3551 963 3609 997
rect 3551 929 3563 963
rect 3597 929 3609 963
rect 3551 895 3609 929
rect 3551 861 3563 895
rect 3597 861 3609 895
rect 3551 827 3609 861
rect 3551 793 3563 827
rect 3597 793 3609 827
rect 3551 759 3609 793
rect 3551 725 3563 759
rect 3597 725 3609 759
rect 3551 691 3609 725
rect 3551 657 3563 691
rect 3597 657 3609 691
rect 3551 623 3609 657
rect 3551 589 3563 623
rect 3597 589 3609 623
rect 3551 555 3609 589
rect 3551 521 3563 555
rect 3597 521 3609 555
rect 3551 487 3609 521
rect 3551 453 3563 487
rect 3597 453 3609 487
rect 3551 419 3609 453
rect 3551 385 3563 419
rect 3597 385 3609 419
rect 3551 351 3609 385
rect 3551 317 3563 351
rect 3597 317 3609 351
rect 3551 278 3609 317
rect 2654 238 2712 272
rect 2654 204 2666 238
rect 2700 204 2712 238
rect 2654 191 2712 204
<< mvpdiff >>
rect 767 3793 825 3836
rect 767 3759 779 3793
rect 813 3759 825 3793
rect 767 3725 825 3759
rect 767 3691 779 3725
rect 813 3691 825 3725
rect 767 3657 825 3691
rect 767 3623 779 3657
rect 813 3623 825 3657
rect 767 3589 825 3623
rect 767 3555 779 3589
rect 813 3555 825 3589
rect 767 3521 825 3555
rect 767 3487 779 3521
rect 813 3487 825 3521
rect 767 3453 825 3487
rect 767 3419 779 3453
rect 813 3419 825 3453
rect 767 3385 825 3419
rect 767 3351 779 3385
rect 813 3351 825 3385
rect 767 3317 825 3351
rect 767 3283 779 3317
rect 813 3283 825 3317
rect 767 3249 825 3283
rect 767 3215 779 3249
rect 813 3215 825 3249
rect 767 3181 825 3215
rect 767 3147 779 3181
rect 813 3147 825 3181
rect 767 3113 825 3147
rect 767 3079 779 3113
rect 813 3079 825 3113
rect 767 3036 825 3079
rect 925 3793 983 3836
rect 925 3759 937 3793
rect 971 3759 983 3793
rect 925 3725 983 3759
rect 925 3691 937 3725
rect 971 3691 983 3725
rect 925 3657 983 3691
rect 925 3623 937 3657
rect 971 3623 983 3657
rect 925 3589 983 3623
rect 925 3555 937 3589
rect 971 3555 983 3589
rect 925 3521 983 3555
rect 925 3487 937 3521
rect 971 3487 983 3521
rect 925 3453 983 3487
rect 925 3419 937 3453
rect 971 3419 983 3453
rect 925 3385 983 3419
rect 925 3351 937 3385
rect 971 3351 983 3385
rect 925 3317 983 3351
rect 925 3283 937 3317
rect 971 3283 983 3317
rect 925 3249 983 3283
rect 925 3215 937 3249
rect 971 3215 983 3249
rect 925 3181 983 3215
rect 925 3147 937 3181
rect 971 3147 983 3181
rect 925 3113 983 3147
rect 925 3079 937 3113
rect 971 3079 983 3113
rect 925 3036 983 3079
rect 1083 3793 1141 3836
rect 1083 3759 1095 3793
rect 1129 3759 1141 3793
rect 1083 3725 1141 3759
rect 2914 3780 2972 3811
rect 1083 3691 1095 3725
rect 1129 3691 1141 3725
rect 1083 3657 1141 3691
rect 1083 3623 1095 3657
rect 1129 3623 1141 3657
rect 1083 3589 1141 3623
rect 2914 3746 2926 3780
rect 2960 3746 2972 3780
rect 2914 3712 2972 3746
rect 2914 3678 2926 3712
rect 2960 3678 2972 3712
rect 2914 3644 2972 3678
rect 1083 3555 1095 3589
rect 1129 3555 1141 3589
rect 2914 3610 2926 3644
rect 2960 3610 2972 3644
rect 1083 3521 1141 3555
rect 2168 3545 2226 3588
rect 1083 3487 1095 3521
rect 1129 3487 1141 3521
rect 1083 3453 1141 3487
rect 1083 3419 1095 3453
rect 1129 3419 1141 3453
rect 1083 3385 1141 3419
rect 1083 3351 1095 3385
rect 1129 3351 1141 3385
rect 1083 3317 1141 3351
rect 1083 3283 1095 3317
rect 1129 3283 1141 3317
rect 1083 3249 1141 3283
rect 1083 3215 1095 3249
rect 1129 3215 1141 3249
rect 1083 3181 1141 3215
rect 1083 3147 1095 3181
rect 1129 3147 1141 3181
rect 1083 3113 1141 3147
rect 1391 3527 1449 3540
rect 1391 3493 1403 3527
rect 1437 3493 1449 3527
rect 1391 3459 1449 3493
rect 1391 3425 1403 3459
rect 1437 3425 1449 3459
rect 1391 3391 1449 3425
rect 1391 3357 1403 3391
rect 1437 3357 1449 3391
rect 1391 3323 1449 3357
rect 1391 3289 1403 3323
rect 1437 3289 1449 3323
rect 1391 3255 1449 3289
rect 1391 3221 1403 3255
rect 1437 3221 1449 3255
rect 1391 3187 1449 3221
rect 1391 3153 1403 3187
rect 1437 3153 1449 3187
rect 1391 3140 1449 3153
rect 1549 3527 1607 3540
rect 1549 3493 1561 3527
rect 1595 3493 1607 3527
rect 1549 3459 1607 3493
rect 1549 3425 1561 3459
rect 1595 3425 1607 3459
rect 1549 3391 1607 3425
rect 1549 3357 1561 3391
rect 1595 3357 1607 3391
rect 1549 3323 1607 3357
rect 1549 3289 1561 3323
rect 1595 3289 1607 3323
rect 1549 3255 1607 3289
rect 1549 3221 1561 3255
rect 1595 3221 1607 3255
rect 1549 3187 1607 3221
rect 1549 3153 1561 3187
rect 1595 3153 1607 3187
rect 1549 3140 1607 3153
rect 2168 3511 2180 3545
rect 2214 3511 2226 3545
rect 2168 3477 2226 3511
rect 2168 3443 2180 3477
rect 2214 3443 2226 3477
rect 2168 3409 2226 3443
rect 2168 3375 2180 3409
rect 2214 3375 2226 3409
rect 2168 3341 2226 3375
rect 2168 3307 2180 3341
rect 2214 3307 2226 3341
rect 2168 3273 2226 3307
rect 2168 3239 2180 3273
rect 2214 3239 2226 3273
rect 2168 3205 2226 3239
rect 2168 3171 2180 3205
rect 2214 3171 2226 3205
rect 1083 3079 1095 3113
rect 1129 3079 1141 3113
rect 1083 3036 1141 3079
rect 2168 3137 2226 3171
rect 2168 3103 2180 3137
rect 2214 3103 2226 3137
rect 2168 3069 2226 3103
rect 2168 3035 2180 3069
rect 2214 3035 2226 3069
rect 1392 2964 1450 3007
rect 1392 2930 1404 2964
rect 1438 2930 1450 2964
rect 1392 2896 1450 2930
rect 1392 2862 1404 2896
rect 1438 2862 1450 2896
rect 1392 2828 1450 2862
rect 1392 2794 1404 2828
rect 1438 2794 1450 2828
rect 1392 2760 1450 2794
rect 1392 2726 1404 2760
rect 1438 2726 1450 2760
rect 1392 2692 1450 2726
rect 1392 2658 1404 2692
rect 1438 2658 1450 2692
rect 1392 2624 1450 2658
rect 1392 2590 1404 2624
rect 1438 2590 1450 2624
rect 1392 2556 1450 2590
rect 1392 2522 1404 2556
rect 1438 2522 1450 2556
rect 1392 2488 1450 2522
rect 1392 2454 1404 2488
rect 1438 2454 1450 2488
rect 1392 2420 1450 2454
rect 1392 2386 1404 2420
rect 1438 2386 1450 2420
rect 1392 2352 1450 2386
rect 1392 2318 1404 2352
rect 1438 2318 1450 2352
rect 1392 2284 1450 2318
rect 1392 2250 1404 2284
rect 1438 2250 1450 2284
rect 1392 2207 1450 2250
rect 1550 2964 1608 3007
rect 1550 2930 1562 2964
rect 1596 2930 1608 2964
rect 1550 2896 1608 2930
rect 1550 2862 1562 2896
rect 1596 2862 1608 2896
rect 1550 2828 1608 2862
rect 1550 2794 1562 2828
rect 1596 2794 1608 2828
rect 1550 2760 1608 2794
rect 1550 2726 1562 2760
rect 1596 2726 1608 2760
rect 1550 2692 1608 2726
rect 1550 2658 1562 2692
rect 1596 2658 1608 2692
rect 1550 2624 1608 2658
rect 1550 2590 1562 2624
rect 1596 2590 1608 2624
rect 1550 2556 1608 2590
rect 1550 2522 1562 2556
rect 1596 2522 1608 2556
rect 1550 2488 1608 2522
rect 1550 2454 1562 2488
rect 1596 2454 1608 2488
rect 1550 2420 1608 2454
rect 1550 2386 1562 2420
rect 1596 2386 1608 2420
rect 1550 2352 1608 2386
rect 1550 2318 1562 2352
rect 1596 2318 1608 2352
rect 1550 2284 1608 2318
rect 1550 2250 1562 2284
rect 1596 2250 1608 2284
rect 1550 2207 1608 2250
rect 1708 2964 1766 3007
rect 1708 2930 1720 2964
rect 1754 2930 1766 2964
rect 1708 2896 1766 2930
rect 1708 2862 1720 2896
rect 1754 2862 1766 2896
rect 1708 2828 1766 2862
rect 1708 2794 1720 2828
rect 1754 2794 1766 2828
rect 1708 2760 1766 2794
rect 2168 3001 2226 3035
rect 2168 2967 2180 3001
rect 2214 2967 2226 3001
rect 2168 2933 2226 2967
rect 2168 2899 2180 2933
rect 2214 2899 2226 2933
rect 2168 2865 2226 2899
rect 2168 2831 2180 2865
rect 2214 2831 2226 2865
rect 2168 2788 2226 2831
rect 2326 3545 2384 3588
rect 2326 3511 2338 3545
rect 2372 3511 2384 3545
rect 2326 3477 2384 3511
rect 2326 3443 2338 3477
rect 2372 3443 2384 3477
rect 2326 3409 2384 3443
rect 2326 3375 2338 3409
rect 2372 3375 2384 3409
rect 2326 3341 2384 3375
rect 2326 3307 2338 3341
rect 2372 3307 2384 3341
rect 2326 3273 2384 3307
rect 2326 3239 2338 3273
rect 2372 3239 2384 3273
rect 2326 3205 2384 3239
rect 2326 3171 2338 3205
rect 2372 3171 2384 3205
rect 2326 3137 2384 3171
rect 2326 3103 2338 3137
rect 2372 3103 2384 3137
rect 2326 3069 2384 3103
rect 2326 3035 2338 3069
rect 2372 3035 2384 3069
rect 2326 3001 2384 3035
rect 2326 2967 2338 3001
rect 2372 2967 2384 3001
rect 2326 2933 2384 2967
rect 2326 2899 2338 2933
rect 2372 2899 2384 2933
rect 2326 2865 2384 2899
rect 2326 2831 2338 2865
rect 2372 2831 2384 2865
rect 2326 2788 2384 2831
rect 2484 3545 2542 3588
rect 2484 3511 2496 3545
rect 2530 3511 2542 3545
rect 2484 3477 2542 3511
rect 2484 3443 2496 3477
rect 2530 3443 2542 3477
rect 2484 3409 2542 3443
rect 2484 3375 2496 3409
rect 2530 3375 2542 3409
rect 2484 3341 2542 3375
rect 2484 3307 2496 3341
rect 2530 3307 2542 3341
rect 2484 3273 2542 3307
rect 2484 3239 2496 3273
rect 2530 3239 2542 3273
rect 2484 3205 2542 3239
rect 2484 3171 2496 3205
rect 2530 3171 2542 3205
rect 2484 3137 2542 3171
rect 2484 3103 2496 3137
rect 2530 3103 2542 3137
rect 2484 3069 2542 3103
rect 2484 3035 2496 3069
rect 2530 3035 2542 3069
rect 2484 3001 2542 3035
rect 2484 2967 2496 3001
rect 2530 2967 2542 3001
rect 2484 2933 2542 2967
rect 2484 2899 2496 2933
rect 2530 2899 2542 2933
rect 2484 2865 2542 2899
rect 2484 2831 2496 2865
rect 2530 2831 2542 2865
rect 2484 2788 2542 2831
rect 2914 3576 2972 3610
rect 2914 3542 2926 3576
rect 2960 3542 2972 3576
rect 2914 3508 2972 3542
rect 2914 3474 2926 3508
rect 2960 3474 2972 3508
rect 2914 3440 2972 3474
rect 2914 3406 2926 3440
rect 2960 3406 2972 3440
rect 2914 3372 2972 3406
rect 2914 3338 2926 3372
rect 2960 3338 2972 3372
rect 2914 3304 2972 3338
rect 2914 3270 2926 3304
rect 2960 3270 2972 3304
rect 2914 3236 2972 3270
rect 2914 3202 2926 3236
rect 2960 3202 2972 3236
rect 2914 3168 2972 3202
rect 2914 3134 2926 3168
rect 2960 3134 2972 3168
rect 2914 3100 2972 3134
rect 2914 3066 2926 3100
rect 2960 3066 2972 3100
rect 2914 3032 2972 3066
rect 2914 2998 2926 3032
rect 2960 2998 2972 3032
rect 2914 2964 2972 2998
rect 2914 2930 2926 2964
rect 2960 2930 2972 2964
rect 2914 2896 2972 2930
rect 2914 2862 2926 2896
rect 2960 2862 2972 2896
rect 2914 2828 2972 2862
rect 2914 2794 2926 2828
rect 2960 2794 2972 2828
rect 1708 2726 1720 2760
rect 1754 2726 1766 2760
rect 1708 2692 1766 2726
rect 1708 2658 1720 2692
rect 1754 2658 1766 2692
rect 1708 2624 1766 2658
rect 1708 2590 1720 2624
rect 1754 2590 1766 2624
rect 2914 2760 2972 2794
rect 2914 2726 2926 2760
rect 2960 2726 2972 2760
rect 2914 2692 2972 2726
rect 2914 2658 2926 2692
rect 2960 2658 2972 2692
rect 2914 2624 2972 2658
rect 1708 2556 1766 2590
rect 1708 2522 1720 2556
rect 1754 2522 1766 2556
rect 1708 2488 1766 2522
rect 2914 2590 2926 2624
rect 2960 2590 2972 2624
rect 2914 2556 2972 2590
rect 2914 2522 2926 2556
rect 2960 2522 2972 2556
rect 1708 2454 1720 2488
rect 1754 2454 1766 2488
rect 1708 2420 1766 2454
rect 1708 2386 1720 2420
rect 1754 2386 1766 2420
rect 1708 2352 1766 2386
rect 1708 2318 1720 2352
rect 1754 2318 1766 2352
rect 1708 2284 1766 2318
rect 1708 2250 1720 2284
rect 1754 2250 1766 2284
rect 1708 2207 1766 2250
rect 2914 2488 2972 2522
rect 2914 2454 2926 2488
rect 2960 2454 2972 2488
rect 2914 2420 2972 2454
rect 2914 2386 2926 2420
rect 2960 2386 2972 2420
rect 2914 2352 2972 2386
rect 2914 2318 2926 2352
rect 2960 2318 2972 2352
rect 2914 2284 2972 2318
rect 2914 2250 2926 2284
rect 2960 2250 2972 2284
rect 2914 2216 2972 2250
rect 2914 2182 2926 2216
rect 2960 2182 2972 2216
rect 2914 2148 2972 2182
rect 2914 2114 2926 2148
rect 2960 2114 2972 2148
rect 2914 2080 2972 2114
rect 2914 2046 2926 2080
rect 2960 2046 2972 2080
rect 2914 2012 2972 2046
rect 2914 1978 2926 2012
rect 2960 1978 2972 2012
rect 2914 1944 2972 1978
rect 2914 1910 2926 1944
rect 2960 1910 2972 1944
rect 2914 1876 2972 1910
rect 2914 1842 2926 1876
rect 2960 1842 2972 1876
rect 2914 1811 2972 1842
rect 3072 3780 3130 3811
rect 3072 3746 3084 3780
rect 3118 3746 3130 3780
rect 3072 3712 3130 3746
rect 3072 3678 3084 3712
rect 3118 3678 3130 3712
rect 3072 3644 3130 3678
rect 3072 3610 3084 3644
rect 3118 3610 3130 3644
rect 3072 3576 3130 3610
rect 3072 3542 3084 3576
rect 3118 3542 3130 3576
rect 3072 3508 3130 3542
rect 3072 3474 3084 3508
rect 3118 3474 3130 3508
rect 3072 3440 3130 3474
rect 3072 3406 3084 3440
rect 3118 3406 3130 3440
rect 3072 3372 3130 3406
rect 3072 3338 3084 3372
rect 3118 3338 3130 3372
rect 3072 3304 3130 3338
rect 3072 3270 3084 3304
rect 3118 3270 3130 3304
rect 3072 3236 3130 3270
rect 3072 3202 3084 3236
rect 3118 3202 3130 3236
rect 3072 3168 3130 3202
rect 3072 3134 3084 3168
rect 3118 3134 3130 3168
rect 3072 3100 3130 3134
rect 3072 3066 3084 3100
rect 3118 3066 3130 3100
rect 3072 3032 3130 3066
rect 3072 2998 3084 3032
rect 3118 2998 3130 3032
rect 3072 2964 3130 2998
rect 3072 2930 3084 2964
rect 3118 2930 3130 2964
rect 3072 2896 3130 2930
rect 3072 2862 3084 2896
rect 3118 2862 3130 2896
rect 3072 2828 3130 2862
rect 3072 2794 3084 2828
rect 3118 2794 3130 2828
rect 3072 2760 3130 2794
rect 3072 2726 3084 2760
rect 3118 2726 3130 2760
rect 3072 2692 3130 2726
rect 3072 2658 3084 2692
rect 3118 2658 3130 2692
rect 3072 2624 3130 2658
rect 3072 2590 3084 2624
rect 3118 2590 3130 2624
rect 3072 2556 3130 2590
rect 3072 2522 3084 2556
rect 3118 2522 3130 2556
rect 3072 2488 3130 2522
rect 3072 2454 3084 2488
rect 3118 2454 3130 2488
rect 3072 2420 3130 2454
rect 3072 2386 3084 2420
rect 3118 2386 3130 2420
rect 3072 2352 3130 2386
rect 3072 2318 3084 2352
rect 3118 2318 3130 2352
rect 3072 2284 3130 2318
rect 3072 2250 3084 2284
rect 3118 2250 3130 2284
rect 3072 2216 3130 2250
rect 3072 2182 3084 2216
rect 3118 2182 3130 2216
rect 3072 2148 3130 2182
rect 3072 2114 3084 2148
rect 3118 2114 3130 2148
rect 3072 2080 3130 2114
rect 3072 2046 3084 2080
rect 3118 2046 3130 2080
rect 3072 2012 3130 2046
rect 3072 1978 3084 2012
rect 3118 1978 3130 2012
rect 3072 1944 3130 1978
rect 3072 1910 3084 1944
rect 3118 1910 3130 1944
rect 3072 1876 3130 1910
rect 3072 1842 3084 1876
rect 3118 1842 3130 1876
rect 3072 1811 3130 1842
rect 3230 3780 3288 3811
rect 3230 3746 3242 3780
rect 3276 3746 3288 3780
rect 3230 3712 3288 3746
rect 3230 3678 3242 3712
rect 3276 3678 3288 3712
rect 3230 3644 3288 3678
rect 3230 3610 3242 3644
rect 3276 3610 3288 3644
rect 3230 3576 3288 3610
rect 3230 3542 3242 3576
rect 3276 3542 3288 3576
rect 3230 3508 3288 3542
rect 3230 3474 3242 3508
rect 3276 3474 3288 3508
rect 3230 3440 3288 3474
rect 3230 3406 3242 3440
rect 3276 3406 3288 3440
rect 3230 3372 3288 3406
rect 3230 3338 3242 3372
rect 3276 3338 3288 3372
rect 3230 3304 3288 3338
rect 3230 3270 3242 3304
rect 3276 3270 3288 3304
rect 3230 3236 3288 3270
rect 3230 3202 3242 3236
rect 3276 3202 3288 3236
rect 3230 3168 3288 3202
rect 3230 3134 3242 3168
rect 3276 3134 3288 3168
rect 3230 3100 3288 3134
rect 3230 3066 3242 3100
rect 3276 3066 3288 3100
rect 3230 3032 3288 3066
rect 3230 2998 3242 3032
rect 3276 2998 3288 3032
rect 3230 2964 3288 2998
rect 3230 2930 3242 2964
rect 3276 2930 3288 2964
rect 3230 2896 3288 2930
rect 3230 2862 3242 2896
rect 3276 2862 3288 2896
rect 3230 2828 3288 2862
rect 3230 2794 3242 2828
rect 3276 2794 3288 2828
rect 3230 2760 3288 2794
rect 3230 2726 3242 2760
rect 3276 2726 3288 2760
rect 3230 2692 3288 2726
rect 3230 2658 3242 2692
rect 3276 2658 3288 2692
rect 3230 2624 3288 2658
rect 3230 2590 3242 2624
rect 3276 2590 3288 2624
rect 3230 2556 3288 2590
rect 3230 2522 3242 2556
rect 3276 2522 3288 2556
rect 3230 2488 3288 2522
rect 3230 2454 3242 2488
rect 3276 2454 3288 2488
rect 3230 2420 3288 2454
rect 3230 2386 3242 2420
rect 3276 2386 3288 2420
rect 3230 2352 3288 2386
rect 3230 2318 3242 2352
rect 3276 2318 3288 2352
rect 3230 2284 3288 2318
rect 3230 2250 3242 2284
rect 3276 2250 3288 2284
rect 3230 2216 3288 2250
rect 3230 2182 3242 2216
rect 3276 2182 3288 2216
rect 3230 2148 3288 2182
rect 3230 2114 3242 2148
rect 3276 2114 3288 2148
rect 3230 2080 3288 2114
rect 3230 2046 3242 2080
rect 3276 2046 3288 2080
rect 3230 2012 3288 2046
rect 3230 1978 3242 2012
rect 3276 1978 3288 2012
rect 3230 1944 3288 1978
rect 3230 1910 3242 1944
rect 3276 1910 3288 1944
rect 3230 1876 3288 1910
rect 3230 1842 3242 1876
rect 3276 1842 3288 1876
rect 3230 1811 3288 1842
rect 3388 3780 3446 3811
rect 3388 3746 3400 3780
rect 3434 3746 3446 3780
rect 3388 3712 3446 3746
rect 3388 3678 3400 3712
rect 3434 3678 3446 3712
rect 3388 3644 3446 3678
rect 3388 3610 3400 3644
rect 3434 3610 3446 3644
rect 3388 3576 3446 3610
rect 3388 3542 3400 3576
rect 3434 3542 3446 3576
rect 3388 3508 3446 3542
rect 3388 3474 3400 3508
rect 3434 3474 3446 3508
rect 3388 3440 3446 3474
rect 3388 3406 3400 3440
rect 3434 3406 3446 3440
rect 3388 3372 3446 3406
rect 3388 3338 3400 3372
rect 3434 3338 3446 3372
rect 3388 3304 3446 3338
rect 3388 3270 3400 3304
rect 3434 3270 3446 3304
rect 3388 3236 3446 3270
rect 3388 3202 3400 3236
rect 3434 3202 3446 3236
rect 3388 3168 3446 3202
rect 3388 3134 3400 3168
rect 3434 3134 3446 3168
rect 3388 3100 3446 3134
rect 3388 3066 3400 3100
rect 3434 3066 3446 3100
rect 3388 3032 3446 3066
rect 3388 2998 3400 3032
rect 3434 2998 3446 3032
rect 3388 2964 3446 2998
rect 3388 2930 3400 2964
rect 3434 2930 3446 2964
rect 3388 2896 3446 2930
rect 3388 2862 3400 2896
rect 3434 2862 3446 2896
rect 3388 2828 3446 2862
rect 3388 2794 3400 2828
rect 3434 2794 3446 2828
rect 3388 2760 3446 2794
rect 3388 2726 3400 2760
rect 3434 2726 3446 2760
rect 3388 2692 3446 2726
rect 3388 2658 3400 2692
rect 3434 2658 3446 2692
rect 3388 2624 3446 2658
rect 3388 2590 3400 2624
rect 3434 2590 3446 2624
rect 3388 2556 3446 2590
rect 3388 2522 3400 2556
rect 3434 2522 3446 2556
rect 3388 2488 3446 2522
rect 3388 2454 3400 2488
rect 3434 2454 3446 2488
rect 3388 2420 3446 2454
rect 3388 2386 3400 2420
rect 3434 2386 3446 2420
rect 3388 2352 3446 2386
rect 3388 2318 3400 2352
rect 3434 2318 3446 2352
rect 3388 2284 3446 2318
rect 3388 2250 3400 2284
rect 3434 2250 3446 2284
rect 3388 2216 3446 2250
rect 3388 2182 3400 2216
rect 3434 2182 3446 2216
rect 3388 2148 3446 2182
rect 3388 2114 3400 2148
rect 3434 2114 3446 2148
rect 3388 2080 3446 2114
rect 3388 2046 3400 2080
rect 3434 2046 3446 2080
rect 3388 2012 3446 2046
rect 3388 1978 3400 2012
rect 3434 1978 3446 2012
rect 3388 1944 3446 1978
rect 3388 1910 3400 1944
rect 3434 1910 3446 1944
rect 3388 1876 3446 1910
rect 3388 1842 3400 1876
rect 3434 1842 3446 1876
rect 3388 1811 3446 1842
rect 3546 3780 3604 3811
rect 3546 3746 3558 3780
rect 3592 3746 3604 3780
rect 3546 3712 3604 3746
rect 3546 3678 3558 3712
rect 3592 3678 3604 3712
rect 3546 3644 3604 3678
rect 3546 3610 3558 3644
rect 3592 3610 3604 3644
rect 3546 3576 3604 3610
rect 3546 3542 3558 3576
rect 3592 3542 3604 3576
rect 3546 3508 3604 3542
rect 3546 3474 3558 3508
rect 3592 3474 3604 3508
rect 3546 3440 3604 3474
rect 3546 3406 3558 3440
rect 3592 3406 3604 3440
rect 3546 3372 3604 3406
rect 3546 3338 3558 3372
rect 3592 3338 3604 3372
rect 3546 3304 3604 3338
rect 3546 3270 3558 3304
rect 3592 3270 3604 3304
rect 3546 3236 3604 3270
rect 3546 3202 3558 3236
rect 3592 3202 3604 3236
rect 3546 3168 3604 3202
rect 3546 3134 3558 3168
rect 3592 3134 3604 3168
rect 3546 3100 3604 3134
rect 3546 3066 3558 3100
rect 3592 3066 3604 3100
rect 3546 3032 3604 3066
rect 3546 2998 3558 3032
rect 3592 2998 3604 3032
rect 3546 2964 3604 2998
rect 3546 2930 3558 2964
rect 3592 2930 3604 2964
rect 3546 2896 3604 2930
rect 3546 2862 3558 2896
rect 3592 2862 3604 2896
rect 3546 2828 3604 2862
rect 3546 2794 3558 2828
rect 3592 2794 3604 2828
rect 3546 2760 3604 2794
rect 3546 2726 3558 2760
rect 3592 2726 3604 2760
rect 3546 2692 3604 2726
rect 3546 2658 3558 2692
rect 3592 2658 3604 2692
rect 3546 2624 3604 2658
rect 3546 2590 3558 2624
rect 3592 2590 3604 2624
rect 3546 2556 3604 2590
rect 3546 2522 3558 2556
rect 3592 2522 3604 2556
rect 3546 2488 3604 2522
rect 3546 2454 3558 2488
rect 3592 2454 3604 2488
rect 3546 2420 3604 2454
rect 3546 2386 3558 2420
rect 3592 2386 3604 2420
rect 3546 2352 3604 2386
rect 3546 2318 3558 2352
rect 3592 2318 3604 2352
rect 3546 2284 3604 2318
rect 3546 2250 3558 2284
rect 3592 2250 3604 2284
rect 3546 2216 3604 2250
rect 3546 2182 3558 2216
rect 3592 2182 3604 2216
rect 3546 2148 3604 2182
rect 3546 2114 3558 2148
rect 3592 2114 3604 2148
rect 3546 2080 3604 2114
rect 3546 2046 3558 2080
rect 3592 2046 3604 2080
rect 3546 2012 3604 2046
rect 3546 1978 3558 2012
rect 3592 1978 3604 2012
rect 3546 1944 3604 1978
rect 3546 1910 3558 1944
rect 3592 1910 3604 1944
rect 3546 1876 3604 1910
rect 3546 1842 3558 1876
rect 3592 1842 3604 1876
rect 3546 1811 3604 1842
rect 1572 1698 1630 1741
rect 1572 1664 1584 1698
rect 1618 1664 1630 1698
rect 1572 1630 1630 1664
rect 1572 1596 1584 1630
rect 1618 1596 1630 1630
rect 1572 1562 1630 1596
rect 1572 1528 1584 1562
rect 1618 1528 1630 1562
rect 1572 1494 1630 1528
rect 1572 1460 1584 1494
rect 1618 1460 1630 1494
rect 1572 1426 1630 1460
rect 1572 1392 1584 1426
rect 1618 1392 1630 1426
rect 1572 1358 1630 1392
rect 1572 1324 1584 1358
rect 1618 1324 1630 1358
rect 1572 1290 1630 1324
rect 1572 1256 1584 1290
rect 1618 1256 1630 1290
rect 1572 1222 1630 1256
rect 1572 1188 1584 1222
rect 1618 1188 1630 1222
rect 1572 1154 1630 1188
rect 1572 1120 1584 1154
rect 1618 1120 1630 1154
rect 1572 1086 1630 1120
rect 1572 1052 1584 1086
rect 1618 1052 1630 1086
rect 1572 1018 1630 1052
rect 1572 984 1584 1018
rect 1618 984 1630 1018
rect 1572 941 1630 984
rect 1730 1698 1788 1741
rect 1730 1664 1742 1698
rect 1776 1664 1788 1698
rect 1730 1630 1788 1664
rect 1730 1596 1742 1630
rect 1776 1596 1788 1630
rect 1730 1562 1788 1596
rect 1730 1528 1742 1562
rect 1776 1528 1788 1562
rect 1730 1494 1788 1528
rect 1730 1460 1742 1494
rect 1776 1460 1788 1494
rect 1730 1426 1788 1460
rect 1730 1392 1742 1426
rect 1776 1392 1788 1426
rect 1730 1358 1788 1392
rect 1730 1324 1742 1358
rect 1776 1324 1788 1358
rect 1730 1290 1788 1324
rect 1730 1256 1742 1290
rect 1776 1256 1788 1290
rect 1730 1222 1788 1256
rect 1730 1188 1742 1222
rect 1776 1188 1788 1222
rect 1730 1154 1788 1188
rect 1730 1120 1742 1154
rect 1776 1120 1788 1154
rect 1730 1086 1788 1120
rect 1730 1052 1742 1086
rect 1776 1052 1788 1086
rect 1730 1018 1788 1052
rect 1730 984 1742 1018
rect 1776 984 1788 1018
rect 1730 941 1788 984
rect 1888 1698 1946 1741
rect 1888 1664 1900 1698
rect 1934 1664 1946 1698
rect 1888 1630 1946 1664
rect 1888 1596 1900 1630
rect 1934 1596 1946 1630
rect 1888 1562 1946 1596
rect 1888 1528 1900 1562
rect 1934 1528 1946 1562
rect 1888 1494 1946 1528
rect 1888 1460 1900 1494
rect 1934 1460 1946 1494
rect 1888 1426 1946 1460
rect 1888 1392 1900 1426
rect 1934 1392 1946 1426
rect 1888 1358 1946 1392
rect 1888 1324 1900 1358
rect 1934 1324 1946 1358
rect 1888 1290 1946 1324
rect 1888 1256 1900 1290
rect 1934 1256 1946 1290
rect 1888 1222 1946 1256
rect 1888 1188 1900 1222
rect 1934 1188 1946 1222
rect 1888 1154 1946 1188
rect 1888 1120 1900 1154
rect 1934 1120 1946 1154
rect 1888 1086 1946 1120
rect 1888 1052 1900 1086
rect 1934 1052 1946 1086
rect 1888 1018 1946 1052
rect 1888 984 1900 1018
rect 1934 984 1946 1018
rect 1888 941 1946 984
rect 1473 691 1531 704
rect 1473 657 1485 691
rect 1519 657 1531 691
rect 1473 623 1531 657
rect 1473 589 1485 623
rect 1519 589 1531 623
rect 1473 555 1531 589
rect 1473 521 1485 555
rect 1519 521 1531 555
rect 1473 487 1531 521
rect 1473 453 1485 487
rect 1519 453 1531 487
rect 1473 419 1531 453
rect 1473 385 1485 419
rect 1519 385 1531 419
rect 1473 351 1531 385
rect 1473 317 1485 351
rect 1519 317 1531 351
rect 1473 304 1531 317
rect 1631 691 1689 704
rect 1631 657 1643 691
rect 1677 657 1689 691
rect 1631 623 1689 657
rect 1631 589 1643 623
rect 1677 589 1689 623
rect 1631 555 1689 589
rect 1631 521 1643 555
rect 1677 521 1689 555
rect 1631 487 1689 521
rect 1631 453 1643 487
rect 1677 453 1689 487
rect 1631 419 1689 453
rect 1631 385 1643 419
rect 1677 385 1689 419
rect 1631 351 1689 385
rect 1631 317 1643 351
rect 1677 317 1689 351
rect 1631 304 1689 317
rect 1869 691 1927 704
rect 1869 657 1881 691
rect 1915 657 1927 691
rect 1869 623 1927 657
rect 1869 589 1881 623
rect 1915 589 1927 623
rect 1869 555 1927 589
rect 1869 521 1881 555
rect 1915 521 1927 555
rect 1869 487 1927 521
rect 1869 453 1881 487
rect 1915 453 1927 487
rect 1869 419 1927 453
rect 1869 385 1881 419
rect 1915 385 1927 419
rect 1869 351 1927 385
rect 1869 317 1881 351
rect 1915 317 1927 351
rect 1869 304 1927 317
rect 2027 691 2085 704
rect 2027 657 2039 691
rect 2073 657 2085 691
rect 2027 623 2085 657
rect 2027 589 2039 623
rect 2073 589 2085 623
rect 2027 555 2085 589
rect 2027 521 2039 555
rect 2073 521 2085 555
rect 2027 487 2085 521
rect 2027 453 2039 487
rect 2073 453 2085 487
rect 2027 419 2085 453
rect 2027 385 2039 419
rect 2073 385 2085 419
rect 2027 351 2085 385
rect 2027 317 2039 351
rect 2073 317 2085 351
rect 2027 304 2085 317
<< mvndiffc >>
rect 879 2655 913 2689
rect 879 2587 913 2621
rect 879 2519 913 2553
rect 879 2451 913 2485
rect 879 2383 913 2417
rect 879 2315 913 2349
rect 1037 2655 1071 2689
rect 1037 2587 1071 2621
rect 1037 2519 1071 2553
rect 1037 2451 1071 2485
rect 1037 2383 1071 2417
rect 1037 2315 1071 2349
rect 2123 2443 2157 2477
rect 2123 2375 2157 2409
rect 2123 2307 2157 2341
rect 2123 2239 2157 2273
rect 2123 2171 2157 2205
rect 2123 2103 2157 2137
rect 2281 2443 2315 2477
rect 2281 2375 2315 2409
rect 2281 2307 2315 2341
rect 2281 2239 2315 2273
rect 2281 2171 2315 2205
rect 2281 2103 2315 2137
rect 2400 2447 2434 2481
rect 2400 2379 2434 2413
rect 2400 2311 2434 2345
rect 2400 2243 2434 2277
rect 2400 2175 2434 2209
rect 2400 2107 2434 2141
rect 2558 2447 2592 2481
rect 2558 2379 2592 2413
rect 2558 2311 2592 2345
rect 2558 2243 2592 2277
rect 2558 2175 2592 2209
rect 2558 2107 2592 2141
rect 949 1674 983 1708
rect 949 1606 983 1640
rect 949 1538 983 1572
rect 949 1470 983 1504
rect 949 1402 983 1436
rect 949 1334 983 1368
rect 1107 1674 1141 1708
rect 1107 1606 1141 1640
rect 1107 1538 1141 1572
rect 1107 1470 1141 1504
rect 1107 1402 1141 1436
rect 1107 1334 1141 1368
rect 1265 1674 1299 1708
rect 1265 1606 1299 1640
rect 1265 1538 1299 1572
rect 1265 1470 1299 1504
rect 1265 1402 1299 1436
rect 1265 1334 1299 1368
rect 953 1099 987 1133
rect 953 1031 987 1065
rect 953 963 987 997
rect 953 895 987 929
rect 953 827 987 861
rect 953 759 987 793
rect 953 691 987 725
rect 953 623 987 657
rect 953 555 987 589
rect 953 487 987 521
rect 953 419 987 453
rect 1111 1099 1145 1133
rect 1111 1031 1145 1065
rect 1111 963 1145 997
rect 2193 1642 2227 1676
rect 2193 1574 2227 1608
rect 2193 1506 2227 1540
rect 2193 1438 2227 1472
rect 2193 1370 2227 1404
rect 2193 1302 2227 1336
rect 2351 1642 2385 1676
rect 2351 1574 2385 1608
rect 2351 1506 2385 1540
rect 2351 1438 2385 1472
rect 2351 1370 2385 1404
rect 2351 1302 2385 1336
rect 2509 1642 2543 1676
rect 2509 1574 2543 1608
rect 2509 1506 2543 1540
rect 2509 1438 2543 1472
rect 2509 1370 2543 1404
rect 2509 1302 2543 1336
rect 2931 1405 2965 1439
rect 2931 1337 2965 1371
rect 2931 1269 2965 1303
rect 2931 1201 2965 1235
rect 2931 1133 2965 1167
rect 2931 1065 2965 1099
rect 2931 997 2965 1031
rect 1111 895 1145 929
rect 2931 929 2965 963
rect 1111 827 1145 861
rect 1111 759 1145 793
rect 1111 691 1145 725
rect 2931 861 2965 895
rect 2931 793 2965 827
rect 1111 623 1145 657
rect 1111 555 1145 589
rect 1111 487 1145 521
rect 1111 419 1145 453
rect 2931 725 2965 759
rect 2931 657 2965 691
rect 2350 544 2384 578
rect 2350 476 2384 510
rect 2350 408 2384 442
rect 2350 340 2384 374
rect 2350 272 2384 306
rect 2350 204 2384 238
rect 2508 544 2542 578
rect 2508 476 2542 510
rect 2508 408 2542 442
rect 2508 340 2542 374
rect 2508 272 2542 306
rect 2508 204 2542 238
rect 2666 544 2700 578
rect 2666 476 2700 510
rect 2666 408 2700 442
rect 2666 340 2700 374
rect 2666 272 2700 306
rect 2931 589 2965 623
rect 2931 521 2965 555
rect 2931 453 2965 487
rect 2931 385 2965 419
rect 2931 317 2965 351
rect 3089 1405 3123 1439
rect 3089 1337 3123 1371
rect 3089 1269 3123 1303
rect 3089 1201 3123 1235
rect 3089 1133 3123 1167
rect 3089 1065 3123 1099
rect 3089 997 3123 1031
rect 3089 929 3123 963
rect 3089 861 3123 895
rect 3089 793 3123 827
rect 3089 725 3123 759
rect 3089 657 3123 691
rect 3089 589 3123 623
rect 3089 521 3123 555
rect 3089 453 3123 487
rect 3089 385 3123 419
rect 3089 317 3123 351
rect 3247 1405 3281 1439
rect 3247 1337 3281 1371
rect 3247 1269 3281 1303
rect 3247 1201 3281 1235
rect 3247 1133 3281 1167
rect 3247 1065 3281 1099
rect 3247 997 3281 1031
rect 3247 929 3281 963
rect 3247 861 3281 895
rect 3247 793 3281 827
rect 3247 725 3281 759
rect 3247 657 3281 691
rect 3247 589 3281 623
rect 3247 521 3281 555
rect 3247 453 3281 487
rect 3247 385 3281 419
rect 3247 317 3281 351
rect 3405 1405 3439 1439
rect 3405 1337 3439 1371
rect 3405 1269 3439 1303
rect 3405 1201 3439 1235
rect 3405 1133 3439 1167
rect 3405 1065 3439 1099
rect 3405 997 3439 1031
rect 3405 929 3439 963
rect 3405 861 3439 895
rect 3405 793 3439 827
rect 3405 725 3439 759
rect 3405 657 3439 691
rect 3405 589 3439 623
rect 3405 521 3439 555
rect 3405 453 3439 487
rect 3405 385 3439 419
rect 3405 317 3439 351
rect 3563 1405 3597 1439
rect 3563 1337 3597 1371
rect 3563 1269 3597 1303
rect 3563 1201 3597 1235
rect 3563 1133 3597 1167
rect 3563 1065 3597 1099
rect 3563 997 3597 1031
rect 3563 929 3597 963
rect 3563 861 3597 895
rect 3563 793 3597 827
rect 3563 725 3597 759
rect 3563 657 3597 691
rect 3563 589 3597 623
rect 3563 521 3597 555
rect 3563 453 3597 487
rect 3563 385 3597 419
rect 3563 317 3597 351
rect 2666 204 2700 238
<< mvpdiffc >>
rect 779 3759 813 3793
rect 779 3691 813 3725
rect 779 3623 813 3657
rect 779 3555 813 3589
rect 779 3487 813 3521
rect 779 3419 813 3453
rect 779 3351 813 3385
rect 779 3283 813 3317
rect 779 3215 813 3249
rect 779 3147 813 3181
rect 779 3079 813 3113
rect 937 3759 971 3793
rect 937 3691 971 3725
rect 937 3623 971 3657
rect 937 3555 971 3589
rect 937 3487 971 3521
rect 937 3419 971 3453
rect 937 3351 971 3385
rect 937 3283 971 3317
rect 937 3215 971 3249
rect 937 3147 971 3181
rect 937 3079 971 3113
rect 1095 3759 1129 3793
rect 1095 3691 1129 3725
rect 1095 3623 1129 3657
rect 2926 3746 2960 3780
rect 2926 3678 2960 3712
rect 1095 3555 1129 3589
rect 2926 3610 2960 3644
rect 1095 3487 1129 3521
rect 1095 3419 1129 3453
rect 1095 3351 1129 3385
rect 1095 3283 1129 3317
rect 1095 3215 1129 3249
rect 1095 3147 1129 3181
rect 1403 3493 1437 3527
rect 1403 3425 1437 3459
rect 1403 3357 1437 3391
rect 1403 3289 1437 3323
rect 1403 3221 1437 3255
rect 1403 3153 1437 3187
rect 1561 3493 1595 3527
rect 1561 3425 1595 3459
rect 1561 3357 1595 3391
rect 1561 3289 1595 3323
rect 1561 3221 1595 3255
rect 1561 3153 1595 3187
rect 2180 3511 2214 3545
rect 2180 3443 2214 3477
rect 2180 3375 2214 3409
rect 2180 3307 2214 3341
rect 2180 3239 2214 3273
rect 2180 3171 2214 3205
rect 1095 3079 1129 3113
rect 2180 3103 2214 3137
rect 2180 3035 2214 3069
rect 1404 2930 1438 2964
rect 1404 2862 1438 2896
rect 1404 2794 1438 2828
rect 1404 2726 1438 2760
rect 1404 2658 1438 2692
rect 1404 2590 1438 2624
rect 1404 2522 1438 2556
rect 1404 2454 1438 2488
rect 1404 2386 1438 2420
rect 1404 2318 1438 2352
rect 1404 2250 1438 2284
rect 1562 2930 1596 2964
rect 1562 2862 1596 2896
rect 1562 2794 1596 2828
rect 1562 2726 1596 2760
rect 1562 2658 1596 2692
rect 1562 2590 1596 2624
rect 1562 2522 1596 2556
rect 1562 2454 1596 2488
rect 1562 2386 1596 2420
rect 1562 2318 1596 2352
rect 1562 2250 1596 2284
rect 1720 2930 1754 2964
rect 1720 2862 1754 2896
rect 1720 2794 1754 2828
rect 2180 2967 2214 3001
rect 2180 2899 2214 2933
rect 2180 2831 2214 2865
rect 2338 3511 2372 3545
rect 2338 3443 2372 3477
rect 2338 3375 2372 3409
rect 2338 3307 2372 3341
rect 2338 3239 2372 3273
rect 2338 3171 2372 3205
rect 2338 3103 2372 3137
rect 2338 3035 2372 3069
rect 2338 2967 2372 3001
rect 2338 2899 2372 2933
rect 2338 2831 2372 2865
rect 2496 3511 2530 3545
rect 2496 3443 2530 3477
rect 2496 3375 2530 3409
rect 2496 3307 2530 3341
rect 2496 3239 2530 3273
rect 2496 3171 2530 3205
rect 2496 3103 2530 3137
rect 2496 3035 2530 3069
rect 2496 2967 2530 3001
rect 2496 2899 2530 2933
rect 2496 2831 2530 2865
rect 2926 3542 2960 3576
rect 2926 3474 2960 3508
rect 2926 3406 2960 3440
rect 2926 3338 2960 3372
rect 2926 3270 2960 3304
rect 2926 3202 2960 3236
rect 2926 3134 2960 3168
rect 2926 3066 2960 3100
rect 2926 2998 2960 3032
rect 2926 2930 2960 2964
rect 2926 2862 2960 2896
rect 2926 2794 2960 2828
rect 1720 2726 1754 2760
rect 1720 2658 1754 2692
rect 1720 2590 1754 2624
rect 2926 2726 2960 2760
rect 2926 2658 2960 2692
rect 1720 2522 1754 2556
rect 2926 2590 2960 2624
rect 2926 2522 2960 2556
rect 1720 2454 1754 2488
rect 1720 2386 1754 2420
rect 1720 2318 1754 2352
rect 1720 2250 1754 2284
rect 2926 2454 2960 2488
rect 2926 2386 2960 2420
rect 2926 2318 2960 2352
rect 2926 2250 2960 2284
rect 2926 2182 2960 2216
rect 2926 2114 2960 2148
rect 2926 2046 2960 2080
rect 2926 1978 2960 2012
rect 2926 1910 2960 1944
rect 2926 1842 2960 1876
rect 3084 3746 3118 3780
rect 3084 3678 3118 3712
rect 3084 3610 3118 3644
rect 3084 3542 3118 3576
rect 3084 3474 3118 3508
rect 3084 3406 3118 3440
rect 3084 3338 3118 3372
rect 3084 3270 3118 3304
rect 3084 3202 3118 3236
rect 3084 3134 3118 3168
rect 3084 3066 3118 3100
rect 3084 2998 3118 3032
rect 3084 2930 3118 2964
rect 3084 2862 3118 2896
rect 3084 2794 3118 2828
rect 3084 2726 3118 2760
rect 3084 2658 3118 2692
rect 3084 2590 3118 2624
rect 3084 2522 3118 2556
rect 3084 2454 3118 2488
rect 3084 2386 3118 2420
rect 3084 2318 3118 2352
rect 3084 2250 3118 2284
rect 3084 2182 3118 2216
rect 3084 2114 3118 2148
rect 3084 2046 3118 2080
rect 3084 1978 3118 2012
rect 3084 1910 3118 1944
rect 3084 1842 3118 1876
rect 3242 3746 3276 3780
rect 3242 3678 3276 3712
rect 3242 3610 3276 3644
rect 3242 3542 3276 3576
rect 3242 3474 3276 3508
rect 3242 3406 3276 3440
rect 3242 3338 3276 3372
rect 3242 3270 3276 3304
rect 3242 3202 3276 3236
rect 3242 3134 3276 3168
rect 3242 3066 3276 3100
rect 3242 2998 3276 3032
rect 3242 2930 3276 2964
rect 3242 2862 3276 2896
rect 3242 2794 3276 2828
rect 3242 2726 3276 2760
rect 3242 2658 3276 2692
rect 3242 2590 3276 2624
rect 3242 2522 3276 2556
rect 3242 2454 3276 2488
rect 3242 2386 3276 2420
rect 3242 2318 3276 2352
rect 3242 2250 3276 2284
rect 3242 2182 3276 2216
rect 3242 2114 3276 2148
rect 3242 2046 3276 2080
rect 3242 1978 3276 2012
rect 3242 1910 3276 1944
rect 3242 1842 3276 1876
rect 3400 3746 3434 3780
rect 3400 3678 3434 3712
rect 3400 3610 3434 3644
rect 3400 3542 3434 3576
rect 3400 3474 3434 3508
rect 3400 3406 3434 3440
rect 3400 3338 3434 3372
rect 3400 3270 3434 3304
rect 3400 3202 3434 3236
rect 3400 3134 3434 3168
rect 3400 3066 3434 3100
rect 3400 2998 3434 3032
rect 3400 2930 3434 2964
rect 3400 2862 3434 2896
rect 3400 2794 3434 2828
rect 3400 2726 3434 2760
rect 3400 2658 3434 2692
rect 3400 2590 3434 2624
rect 3400 2522 3434 2556
rect 3400 2454 3434 2488
rect 3400 2386 3434 2420
rect 3400 2318 3434 2352
rect 3400 2250 3434 2284
rect 3400 2182 3434 2216
rect 3400 2114 3434 2148
rect 3400 2046 3434 2080
rect 3400 1978 3434 2012
rect 3400 1910 3434 1944
rect 3400 1842 3434 1876
rect 3558 3746 3592 3780
rect 3558 3678 3592 3712
rect 3558 3610 3592 3644
rect 3558 3542 3592 3576
rect 3558 3474 3592 3508
rect 3558 3406 3592 3440
rect 3558 3338 3592 3372
rect 3558 3270 3592 3304
rect 3558 3202 3592 3236
rect 3558 3134 3592 3168
rect 3558 3066 3592 3100
rect 3558 2998 3592 3032
rect 3558 2930 3592 2964
rect 3558 2862 3592 2896
rect 3558 2794 3592 2828
rect 3558 2726 3592 2760
rect 3558 2658 3592 2692
rect 3558 2590 3592 2624
rect 3558 2522 3592 2556
rect 3558 2454 3592 2488
rect 3558 2386 3592 2420
rect 3558 2318 3592 2352
rect 3558 2250 3592 2284
rect 3558 2182 3592 2216
rect 3558 2114 3592 2148
rect 3558 2046 3592 2080
rect 3558 1978 3592 2012
rect 3558 1910 3592 1944
rect 3558 1842 3592 1876
rect 1584 1664 1618 1698
rect 1584 1596 1618 1630
rect 1584 1528 1618 1562
rect 1584 1460 1618 1494
rect 1584 1392 1618 1426
rect 1584 1324 1618 1358
rect 1584 1256 1618 1290
rect 1584 1188 1618 1222
rect 1584 1120 1618 1154
rect 1584 1052 1618 1086
rect 1584 984 1618 1018
rect 1742 1664 1776 1698
rect 1742 1596 1776 1630
rect 1742 1528 1776 1562
rect 1742 1460 1776 1494
rect 1742 1392 1776 1426
rect 1742 1324 1776 1358
rect 1742 1256 1776 1290
rect 1742 1188 1776 1222
rect 1742 1120 1776 1154
rect 1742 1052 1776 1086
rect 1742 984 1776 1018
rect 1900 1664 1934 1698
rect 1900 1596 1934 1630
rect 1900 1528 1934 1562
rect 1900 1460 1934 1494
rect 1900 1392 1934 1426
rect 1900 1324 1934 1358
rect 1900 1256 1934 1290
rect 1900 1188 1934 1222
rect 1900 1120 1934 1154
rect 1900 1052 1934 1086
rect 1900 984 1934 1018
rect 1485 657 1519 691
rect 1485 589 1519 623
rect 1485 521 1519 555
rect 1485 453 1519 487
rect 1485 385 1519 419
rect 1485 317 1519 351
rect 1643 657 1677 691
rect 1643 589 1677 623
rect 1643 521 1677 555
rect 1643 453 1677 487
rect 1643 385 1677 419
rect 1643 317 1677 351
rect 1881 657 1915 691
rect 1881 589 1915 623
rect 1881 521 1915 555
rect 1881 453 1915 487
rect 1881 385 1915 419
rect 1881 317 1915 351
rect 2039 657 2073 691
rect 2039 589 2073 623
rect 2039 521 2073 555
rect 2039 453 2073 487
rect 2039 385 2073 419
rect 2039 317 2073 351
<< psubdiff >>
rect -464 93 1213 131
rect -464 59 -398 93
rect -364 59 -167 93
rect -133 59 116 93
rect 150 59 305 93
rect 339 59 479 93
rect 513 59 662 93
rect 696 59 849 93
rect 883 59 1052 93
rect 1086 59 1213 93
rect -464 22 1213 59
<< mvnsubdiff >>
rect 1202 3868 1886 3877
rect 1202 3863 2734 3868
rect 1202 3829 1271 3863
rect 1305 3829 1409 3863
rect 1202 3795 1409 3829
rect 1202 3761 1271 3795
rect 1305 3761 1409 3795
rect 1511 3761 1678 3863
rect 1780 3831 2734 3863
rect 1780 3797 1996 3831
rect 2030 3797 2185 3831
rect 2219 3797 2379 3831
rect 2413 3797 2584 3831
rect 2618 3797 2734 3831
rect 1780 3761 2734 3797
rect 1202 3760 2734 3761
rect 1202 3748 1886 3760
<< psubdiffcont >>
rect -398 59 -364 93
rect -167 59 -133 93
rect 116 59 150 93
rect 305 59 339 93
rect 479 59 513 93
rect 662 59 696 93
rect 849 59 883 93
rect 1052 59 1086 93
<< mvnsubdiffcont >>
rect 1271 3829 1305 3863
rect 1271 3761 1305 3795
rect 1409 3761 1511 3863
rect 1678 3761 1780 3863
rect 1996 3797 2030 3831
rect 2185 3797 2219 3831
rect 2379 3797 2413 3831
rect 2584 3797 2618 3831
<< poly >>
rect -156 3860 -90 3876
rect -156 3826 -140 3860
rect -106 3826 -90 3860
rect -156 3446 -90 3826
rect -804 1768 -738 2148
rect -804 1734 -788 1768
rect -754 1734 -738 1768
rect -804 1718 -738 1734
rect -180 2032 -114 2048
rect -180 1998 -164 2032
rect -130 1998 -114 2032
rect -180 1618 -114 1998
rect 10 1341 76 1721
rect 10 1307 26 1341
rect 60 1307 76 1341
rect 10 1291 76 1307
rect 825 3836 925 3862
rect 983 3836 1083 3862
rect 2972 3811 3072 3837
rect 3130 3811 3230 3837
rect 3288 3811 3388 3837
rect 3446 3811 3546 3837
rect 2226 3588 2326 3614
rect 2384 3588 2484 3614
rect 1449 3540 1549 3566
rect 1230 3121 1284 3134
rect 1449 3121 1549 3140
rect 1230 3118 1549 3121
rect 1230 3084 1240 3118
rect 1274 3114 1549 3118
rect 1274 3084 1520 3114
rect 1230 3081 1520 3084
rect 1230 3068 1284 3081
rect 825 3010 925 3036
rect 983 3010 1083 3036
rect 716 2935 770 2950
rect 854 2935 891 3010
rect 1012 2944 1049 3010
rect 1450 3007 1550 3033
rect 1608 3007 1708 3033
rect 986 2935 1052 2944
rect 716 2934 1052 2935
rect 716 2900 726 2934
rect 760 2900 1002 2934
rect 1036 2900 1052 2934
rect 716 2898 1052 2900
rect 716 2884 770 2898
rect 986 2890 1052 2898
rect 940 2818 1006 2828
rect 940 2784 956 2818
rect 990 2784 1006 2818
rect 940 2774 1006 2784
rect 958 2732 988 2774
rect 958 2728 992 2732
rect 925 2702 1025 2728
rect 925 2276 1025 2302
rect 2226 2762 2326 2788
rect 2384 2762 2484 2788
rect 2258 2647 2304 2762
rect 2248 2643 2314 2647
rect 2421 2643 2467 2762
rect 2248 2637 2467 2643
rect 2248 2603 2264 2637
rect 2298 2603 2467 2637
rect 2248 2597 2467 2603
rect 2248 2593 2314 2597
rect 2169 2490 2269 2516
rect 2446 2494 2546 2520
rect 1450 2181 1550 2207
rect 1608 2181 1708 2207
rect 1478 2063 1518 2181
rect 1638 2064 1675 2181
rect 2169 2064 2269 2090
rect 2446 2068 2546 2094
rect 1471 2047 1525 2063
rect 1471 2013 1481 2047
rect 1515 2013 1525 2047
rect 1471 1997 1525 2013
rect 1630 2048 1684 2064
rect 1630 2014 1640 2048
rect 1674 2014 1684 2048
rect 1630 1998 1684 2014
rect 2203 2019 2246 2064
rect 2483 2019 2526 2068
rect 2203 1976 2693 2019
rect 2650 1895 2693 1976
rect 2645 1879 2699 1895
rect 1014 1845 1068 1861
rect 1014 1811 1024 1845
rect 1058 1811 1068 1845
rect 1014 1795 1068 1811
rect 1177 1841 1231 1857
rect 1177 1807 1187 1841
rect 1221 1807 1231 1841
rect 1020 1747 1062 1795
rect 1177 1791 1231 1807
rect 2337 1842 2391 1858
rect 2337 1808 2347 1842
rect 2381 1808 2391 1842
rect 2645 1845 2655 1879
rect 2689 1845 2699 1879
rect 2645 1829 2699 1845
rect 2337 1798 2391 1808
rect 1184 1747 1223 1791
rect 995 1721 1095 1747
rect 1153 1721 1253 1747
rect 1630 1741 1730 1767
rect 1788 1741 1888 1767
rect 2274 1758 2457 1798
rect 550 1341 616 1721
rect 550 1307 566 1341
rect 600 1307 616 1341
rect 550 1291 616 1307
rect 995 1295 1095 1321
rect 1153 1295 1253 1321
rect 999 1176 1099 1202
rect -612 110 -546 490
rect 2274 1715 2314 1758
rect 2417 1715 2457 1758
rect 2972 1764 3072 1811
rect 2972 1730 3005 1764
rect 3039 1730 3072 1764
rect 2239 1689 2339 1715
rect 2397 1689 2497 1715
rect 2972 1714 3072 1730
rect 3130 1764 3230 1811
rect 3130 1730 3163 1764
rect 3197 1730 3230 1764
rect 3130 1714 3230 1730
rect 3288 1764 3388 1811
rect 3288 1730 3321 1764
rect 3355 1730 3388 1764
rect 3288 1714 3388 1730
rect 3446 1764 3546 1811
rect 3446 1730 3479 1764
rect 3513 1730 3546 1764
rect 3446 1714 3546 1730
rect 2977 1550 3077 1566
rect 2977 1516 3010 1550
rect 3044 1516 3077 1550
rect 2977 1478 3077 1516
rect 3135 1550 3235 1566
rect 3135 1516 3168 1550
rect 3202 1516 3235 1550
rect 3135 1478 3235 1516
rect 3293 1550 3393 1566
rect 3293 1516 3326 1550
rect 3360 1516 3393 1550
rect 3293 1478 3393 1516
rect 3451 1550 3551 1566
rect 3451 1516 3484 1550
rect 3518 1516 3551 1550
rect 3451 1478 3551 1516
rect 2239 1263 2339 1289
rect 2397 1263 2497 1289
rect 1630 915 1730 941
rect 1788 915 1888 941
rect 1662 831 1712 915
rect 1814 831 1864 915
rect 1379 781 1864 831
rect 1379 720 1429 781
rect 2280 770 2346 778
rect 2280 768 2626 770
rect 2280 734 2296 768
rect 2330 734 2626 768
rect 2280 731 2626 734
rect 1371 710 1437 720
rect 1371 676 1387 710
rect 1421 676 1437 710
rect 1531 704 1631 730
rect 1927 704 2027 730
rect 2280 724 2346 731
rect 1371 666 1437 676
rect 999 350 1099 376
rect 1033 259 1073 350
rect 2423 617 2462 731
rect 2587 617 2626 731
rect 2396 591 2496 617
rect 2554 591 2654 617
rect 1531 278 1631 304
rect 1927 278 2027 304
rect 1026 243 1080 259
rect 1026 209 1036 243
rect 1070 209 1080 243
rect 1026 193 1080 209
rect 1351 208 1417 218
rect 1567 208 1601 278
rect 1961 208 1995 278
rect 2113 208 2179 218
rect 1351 174 1367 208
rect 1401 174 2129 208
rect 2163 174 2179 208
rect 2977 252 3077 278
rect 3135 252 3235 278
rect 3293 252 3393 278
rect 3451 252 3551 278
rect 1351 164 1417 174
rect 2113 164 2179 174
rect 2396 165 2496 191
rect 2554 165 2654 191
rect -612 76 -596 110
rect -562 76 -546 110
rect -612 60 -546 76
<< polycont >>
rect -140 3826 -106 3860
rect -788 1734 -754 1768
rect -164 1998 -130 2032
rect 26 1307 60 1341
rect 1240 3084 1274 3118
rect 726 2900 760 2934
rect 1002 2900 1036 2934
rect 956 2784 990 2818
rect 2264 2603 2298 2637
rect 1481 2013 1515 2047
rect 1640 2014 1674 2048
rect 1024 1811 1058 1845
rect 1187 1807 1221 1841
rect 2347 1808 2381 1842
rect 2655 1845 2689 1879
rect 566 1307 600 1341
rect 3005 1730 3039 1764
rect 3163 1730 3197 1764
rect 3321 1730 3355 1764
rect 3479 1730 3513 1764
rect 3010 1516 3044 1550
rect 3168 1516 3202 1550
rect 3326 1516 3360 1550
rect 3484 1516 3518 1550
rect 2296 734 2330 768
rect 1387 676 1421 710
rect 1036 209 1070 243
rect 1367 174 1401 208
rect 2129 174 2163 208
rect -596 76 -562 110
<< npolyres >>
rect 10 3919 184 3985
rect -804 3276 -630 3342
rect -804 2148 -738 3276
rect -696 2318 -630 3276
rect -588 3276 -414 3342
rect -588 2318 -522 3276
rect -696 2252 -522 2318
rect -480 2318 -414 3276
rect -372 3276 -198 3342
rect -372 2318 -306 3276
rect -480 2252 -306 2318
rect -264 2318 -198 3276
rect -156 2318 -90 3446
rect -264 2252 -90 2318
rect -612 1448 -438 1514
rect -612 490 -546 1448
rect -504 660 -438 1448
rect -396 1448 -222 1514
rect -396 660 -330 1448
rect -504 594 -330 660
rect -288 660 -222 1448
rect -180 660 -114 1618
rect 10 1721 76 3919
rect 118 1891 184 3919
rect 226 3919 400 3985
rect 226 1891 292 3919
rect 118 1825 292 1891
rect 334 1891 400 3919
rect 442 3919 616 3985
rect 442 1891 508 3919
rect 334 1825 508 1891
rect 550 1721 616 3919
rect -288 594 -114 660
<< locali >>
rect 1862 3900 2788 3933
rect -162 3860 -88 3878
rect -162 3858 -140 3860
rect -162 3824 -142 3858
rect -106 3826 -88 3860
rect 1172 3863 2788 3900
rect -108 3824 -88 3826
rect -162 3786 -88 3824
rect 779 3813 813 3840
rect 779 3741 813 3759
rect 779 3669 813 3691
rect 779 3597 813 3623
rect 779 3525 813 3555
rect 779 3453 813 3487
rect 779 3385 813 3419
rect 779 3317 813 3347
rect 779 3249 813 3275
rect 779 3181 813 3203
rect 779 3113 813 3131
rect 775 3059 779 3088
rect 775 3032 813 3059
rect 937 3813 971 3840
rect 937 3741 971 3759
rect 937 3669 971 3691
rect 937 3597 971 3623
rect 937 3525 971 3555
rect 937 3453 971 3487
rect 937 3385 971 3419
rect 937 3317 971 3347
rect 937 3249 971 3275
rect 937 3181 971 3203
rect 937 3113 971 3131
rect 937 3032 971 3059
rect 1095 3813 1129 3840
rect 1095 3741 1129 3759
rect 1172 3829 1271 3863
rect 1305 3836 1409 3863
rect 1305 3829 1353 3836
rect 1172 3802 1353 3829
rect 1387 3802 1409 3836
rect 1172 3795 1409 3802
rect 1172 3761 1271 3795
rect 1305 3761 1409 3795
rect 1511 3831 1678 3863
rect 1511 3797 1577 3831
rect 1611 3797 1678 3831
rect 1511 3761 1678 3797
rect 1780 3833 2788 3863
rect 1780 3831 2537 3833
rect 1780 3828 1996 3831
rect 1780 3794 1820 3828
rect 1854 3797 1996 3828
rect 2030 3830 2185 3831
rect 2030 3797 2043 3830
rect 1854 3796 2043 3797
rect 2077 3796 2115 3830
rect 2149 3797 2185 3830
rect 2219 3828 2379 3831
rect 2219 3797 2278 3828
rect 2149 3796 2278 3797
rect 1854 3794 2278 3796
rect 2312 3794 2350 3828
rect 2413 3799 2537 3831
rect 2571 3831 2609 3833
rect 2571 3799 2584 3831
rect 2643 3799 2788 3833
rect 2413 3797 2584 3799
rect 2618 3797 2788 3799
rect 2384 3794 2788 3797
rect 1780 3761 2788 3794
rect 2919 3916 3596 3923
rect 2919 3882 2926 3916
rect 2960 3882 3596 3916
rect 2919 3875 3596 3882
rect 2919 3783 2967 3875
rect 1172 3718 2788 3761
rect 1862 3717 2788 3718
rect 2926 3780 2960 3783
rect 1095 3669 1129 3691
rect 1095 3597 1129 3623
rect 2926 3712 2960 3730
rect 2926 3644 2960 3658
rect 1095 3525 1129 3555
rect 2180 3565 2214 3592
rect 1095 3453 1129 3487
rect 1095 3385 1129 3419
rect 1095 3317 1129 3347
rect 1095 3249 1129 3275
rect 1095 3181 1129 3203
rect 1403 3527 1437 3544
rect 1403 3459 1437 3467
rect 1403 3391 1437 3395
rect 1403 3285 1437 3289
rect 1403 3213 1437 3221
rect 1403 3136 1437 3153
rect 1561 3527 1595 3544
rect 1561 3459 1595 3467
rect 1561 3391 1595 3395
rect 1561 3285 1595 3289
rect 1561 3213 1595 3221
rect 1561 3136 1595 3153
rect 2180 3493 2214 3511
rect 2180 3421 2214 3443
rect 2180 3349 2214 3375
rect 2180 3277 2214 3307
rect 2180 3205 2214 3239
rect 2180 3137 2214 3171
rect 1095 3113 1129 3131
rect 1237 3118 1277 3121
rect 1224 3084 1240 3118
rect 1274 3084 1290 3118
rect 1237 3081 1277 3084
rect 775 3022 812 3032
rect 725 2985 812 3022
rect 725 2950 762 2985
rect 660 2934 770 2950
rect 1002 2936 1036 2950
rect 1001 2934 1038 2936
rect 660 2900 726 2934
rect 760 2900 776 2934
rect 1001 2900 1002 2934
rect 1036 2900 1038 2934
rect 660 2867 770 2900
rect 1001 2899 1038 2900
rect 1002 2884 1036 2899
rect -185 2032 -119 2047
rect -185 1998 -164 2032
rect -130 1998 -114 2032
rect -185 1788 -119 1998
rect -812 1768 -119 1788
rect -812 1734 -788 1768
rect -754 1734 -119 1768
rect -812 1722 -119 1734
rect -187 340 -121 1722
rect 660 1359 724 2867
rect 956 2818 990 2834
rect 1095 2818 1129 3059
rect 2180 3069 2214 3099
rect 990 2784 1129 2818
rect 1404 2984 1438 3011
rect 1404 2912 1438 2930
rect 1404 2840 1438 2862
rect 956 2768 990 2784
rect 879 2689 913 2706
rect 879 2621 913 2629
rect 879 2553 913 2557
rect 1037 2704 1072 2784
rect 1404 2768 1438 2794
rect 1037 2689 1071 2704
rect 1037 2621 1071 2629
rect 1037 2553 1071 2557
rect 879 2447 913 2451
rect 879 2375 913 2383
rect 879 2298 913 2315
rect 1030 2451 1037 2509
rect 1030 2447 1071 2451
rect 1030 2383 1037 2447
rect 1030 2375 1071 2383
rect 1030 2315 1037 2375
rect 1030 2298 1071 2315
rect 1404 2696 1438 2726
rect 1404 2624 1438 2658
rect 1404 2556 1438 2590
rect 1404 2488 1438 2518
rect 1404 2420 1438 2446
rect 1404 2352 1438 2374
rect 1030 2146 1067 2298
rect 1404 2284 1438 2302
rect 1404 2203 1438 2230
rect 1562 2984 1596 3011
rect 1562 2912 1596 2930
rect 1562 2840 1596 2862
rect 1562 2768 1596 2794
rect 1562 2696 1596 2726
rect 1562 2624 1596 2658
rect 1562 2556 1596 2590
rect 1562 2488 1596 2518
rect 1562 2420 1596 2446
rect 1562 2352 1596 2374
rect 1562 2284 1596 2302
rect 1562 2203 1596 2230
rect 1720 2984 1754 3011
rect 1720 2912 1754 2930
rect 2180 3001 2214 3027
rect 2180 2933 2214 2955
rect 2180 2879 2214 2883
rect 2338 3565 2372 3592
rect 2338 3493 2372 3511
rect 2338 3421 2372 3443
rect 2338 3349 2372 3375
rect 2338 3277 2372 3307
rect 2338 3205 2372 3239
rect 2338 3137 2372 3171
rect 2338 3069 2372 3099
rect 2338 3001 2372 3027
rect 2338 2933 2372 2955
rect 1720 2840 1754 2862
rect 1720 2768 1754 2794
rect 1720 2696 1754 2726
rect 1720 2624 1754 2658
rect 2171 2865 2217 2879
rect 2171 2811 2180 2865
rect 2214 2811 2217 2865
rect 2171 2643 2217 2811
rect 2338 2865 2372 2883
rect 2338 2784 2372 2811
rect 2496 3565 2530 3592
rect 2496 3493 2530 3511
rect 2496 3421 2530 3443
rect 2496 3349 2530 3375
rect 2496 3277 2530 3307
rect 2496 3205 2530 3239
rect 2496 3137 2530 3171
rect 2496 3069 2530 3099
rect 2496 3001 2530 3027
rect 2496 2933 2530 2955
rect 2496 2865 2530 2883
rect 2496 2784 2530 2811
rect 2926 3576 2960 3586
rect 2926 3508 2960 3514
rect 2926 3440 2960 3442
rect 2926 3404 2960 3406
rect 2926 3332 2960 3338
rect 2926 3260 2960 3270
rect 2926 3188 2960 3202
rect 2926 3116 2960 3134
rect 2926 3044 2960 3066
rect 2926 2972 2960 2998
rect 2926 2900 2960 2930
rect 2926 2828 2960 2862
rect 2926 2760 2960 2794
rect 2926 2692 2960 2722
rect 2264 2643 2298 2653
rect 2613 2645 2783 2651
rect 2171 2637 2304 2643
rect 2171 2603 2264 2637
rect 2298 2603 2304 2637
rect 2613 2611 2618 2645
rect 2652 2611 2783 2645
rect 2613 2606 2783 2611
rect 2670 2604 2783 2606
rect 2171 2597 2304 2603
rect 1720 2556 1754 2590
rect 2264 2587 2298 2597
rect 1720 2488 1754 2518
rect 1720 2420 1754 2446
rect 1720 2352 1754 2374
rect 1720 2301 1754 2302
rect 2123 2477 2157 2494
rect 2123 2409 2157 2417
rect 2123 2341 2157 2345
rect 1720 2284 2048 2301
rect 1754 2258 2048 2284
rect 1720 2203 1754 2230
rect 1030 2106 1918 2146
rect 1030 2076 1067 2106
rect 0 1341 171 1354
rect 0 1307 26 1341
rect 60 1340 171 1341
rect 60 1307 123 1340
rect 0 1306 123 1307
rect 157 1306 171 1340
rect 0 1293 171 1306
rect 542 1341 724 1359
rect 542 1307 566 1341
rect 600 1307 724 1341
rect 542 1276 724 1307
rect 765 2039 1067 2076
rect 1478 2047 1518 2050
rect 1639 2048 1676 2050
rect 163 990 567 993
rect 163 956 165 990
rect 199 956 530 990
rect 564 956 567 990
rect 163 954 567 956
rect 619 711 669 1276
rect 619 677 627 711
rect 661 677 669 711
rect 619 669 669 677
rect 682 340 716 343
rect -187 306 682 340
rect 682 303 716 306
rect 765 244 802 2039
rect 1465 2013 1481 2047
rect 1515 2013 1531 2047
rect 1624 2014 1640 2048
rect 1674 2014 1690 2048
rect 1478 1958 1518 2013
rect 1020 1956 1518 1958
rect 1020 1922 1417 1956
rect 1451 1922 1518 1956
rect 1020 1918 1518 1922
rect 1020 1882 1060 1918
rect 1639 1884 1676 2014
rect 1020 1845 1062 1882
rect 1185 1845 1676 1884
rect 1878 1903 1918 2106
rect 2005 2029 2048 2258
rect 2123 2235 2157 2239
rect 2123 2163 2157 2171
rect 2123 2086 2157 2103
rect 2281 2477 2315 2494
rect 2281 2409 2315 2417
rect 2281 2341 2315 2345
rect 2281 2235 2315 2239
rect 2281 2163 2315 2171
rect 2281 2086 2315 2103
rect 2400 2481 2434 2498
rect 2400 2413 2434 2421
rect 2400 2345 2434 2349
rect 2400 2239 2434 2243
rect 2400 2167 2434 2175
rect 2400 2090 2434 2107
rect 2558 2481 2592 2498
rect 2558 2413 2592 2421
rect 2558 2345 2592 2349
rect 2736 2362 2783 2604
rect 2736 2328 2742 2362
rect 2776 2328 2783 2362
rect 2736 2322 2783 2328
rect 2926 2624 2960 2650
rect 2926 2556 2960 2578
rect 2926 2488 2960 2506
rect 2926 2420 2960 2434
rect 2926 2352 2960 2362
rect 2558 2239 2592 2243
rect 2558 2167 2592 2175
rect 2558 2090 2592 2107
rect 2926 2284 2960 2290
rect 2926 2216 2960 2218
rect 2926 2180 2960 2182
rect 2926 2108 2960 2114
rect 2926 2036 2960 2046
rect 2005 1999 2560 2029
rect 2005 1986 2521 1999
rect 2555 1986 2560 1999
rect 2926 1964 2960 1978
rect 2834 1911 2883 1919
rect 2344 1903 2384 1904
rect 1878 1863 2384 1903
rect 2651 1879 2694 1884
rect 1008 1811 1024 1845
rect 1058 1811 1074 1845
rect 1185 1841 1237 1845
rect 1020 1807 1062 1811
rect 1171 1807 1187 1841
rect 1221 1807 1237 1841
rect 1185 1805 1224 1807
rect 949 1708 983 1725
rect 949 1640 983 1648
rect 949 1572 983 1576
rect 949 1466 983 1470
rect 949 1394 983 1402
rect 949 1317 983 1334
rect 1107 1708 1141 1725
rect 1107 1640 1141 1648
rect 1107 1572 1141 1576
rect 1107 1466 1141 1470
rect 1107 1394 1141 1402
rect 1107 1317 1141 1334
rect 1265 1708 1299 1725
rect 1265 1640 1299 1648
rect 1265 1572 1299 1576
rect 1265 1466 1299 1470
rect 1366 1443 1405 1845
rect 2331 1842 2384 1863
rect 2639 1845 2655 1879
rect 2689 1845 2705 1879
rect 2834 1877 2841 1911
rect 2875 1877 2883 1911
rect 2331 1808 2347 1842
rect 2381 1808 2397 1842
rect 2344 1805 2384 1808
rect 1366 1409 1368 1443
rect 1402 1409 1405 1443
rect 1366 1407 1405 1409
rect 1584 1718 1618 1745
rect 1584 1646 1618 1664
rect 1584 1574 1618 1596
rect 1584 1502 1618 1528
rect 1584 1430 1618 1460
rect 1265 1394 1299 1402
rect 1265 1317 1299 1334
rect 1584 1358 1618 1392
rect 1584 1290 1618 1324
rect 1584 1222 1618 1252
rect 1312 1186 1361 1194
rect 953 1153 987 1180
rect 953 1081 987 1099
rect 953 1009 987 1031
rect 953 937 987 963
rect 953 865 987 895
rect 953 793 987 827
rect 953 725 987 759
rect 953 657 987 687
rect 953 589 987 615
rect 953 521 987 543
rect 953 453 987 471
rect 953 372 987 399
rect 1111 1153 1145 1180
rect 1111 1081 1145 1099
rect 1111 1009 1145 1031
rect 1111 937 1145 963
rect 1111 865 1145 895
rect 1111 793 1145 827
rect 1312 1152 1319 1186
rect 1353 1152 1361 1186
rect 1312 853 1361 1152
rect 1584 1154 1618 1180
rect 1584 1086 1618 1108
rect 1584 1018 1618 1036
rect 1584 937 1618 964
rect 1742 1718 1776 1745
rect 1742 1646 1776 1664
rect 1742 1574 1776 1596
rect 1742 1502 1776 1528
rect 1742 1430 1776 1460
rect 1742 1358 1776 1392
rect 1742 1290 1776 1324
rect 1742 1222 1776 1252
rect 1742 1154 1776 1180
rect 1742 1086 1776 1108
rect 1742 1018 1776 1036
rect 1742 937 1776 964
rect 1900 1718 1934 1745
rect 1900 1646 1934 1664
rect 1900 1574 1934 1596
rect 1900 1502 1934 1528
rect 1900 1430 1934 1460
rect 1900 1358 1934 1392
rect 1900 1290 1934 1324
rect 2193 1676 2227 1693
rect 2193 1608 2227 1616
rect 2193 1540 2227 1544
rect 2193 1434 2227 1438
rect 2193 1362 2227 1370
rect 2193 1285 2227 1302
rect 2351 1676 2385 1693
rect 2351 1608 2385 1616
rect 2351 1540 2385 1544
rect 2351 1434 2385 1438
rect 2351 1362 2385 1370
rect 2351 1285 2385 1302
rect 2509 1676 2543 1693
rect 2509 1608 2543 1616
rect 2509 1540 2543 1544
rect 2509 1434 2543 1438
rect 2509 1362 2543 1370
rect 2509 1285 2543 1302
rect 1900 1222 1934 1252
rect 2651 1246 2694 1845
rect 2834 1676 2883 1877
rect 2926 1892 2960 1910
rect 2926 1807 2960 1842
rect 3084 3780 3118 3815
rect 3234 3780 3282 3875
rect 3548 3846 3596 3875
rect 3548 3823 3598 3846
rect 3234 3778 3242 3780
rect 3084 3712 3118 3730
rect 3084 3644 3118 3658
rect 3084 3576 3118 3586
rect 3084 3508 3118 3514
rect 3084 3440 3118 3442
rect 3084 3404 3118 3406
rect 3084 3332 3118 3338
rect 3084 3260 3118 3270
rect 3084 3188 3118 3202
rect 3084 3116 3118 3134
rect 3084 3044 3118 3066
rect 3084 2972 3118 2998
rect 3084 2900 3118 2930
rect 3084 2828 3118 2862
rect 3084 2760 3118 2794
rect 3084 2692 3118 2722
rect 3084 2624 3118 2650
rect 3084 2556 3118 2578
rect 3084 2488 3118 2506
rect 3084 2420 3118 2434
rect 3084 2352 3118 2362
rect 3084 2284 3118 2290
rect 3084 2216 3118 2218
rect 3084 2180 3118 2182
rect 3084 2108 3118 2114
rect 3084 2036 3118 2046
rect 3084 1964 3118 1978
rect 3084 1892 3118 1910
rect 3084 1807 3118 1842
rect 3276 3778 3282 3780
rect 3400 3780 3434 3815
rect 3242 3712 3276 3730
rect 3242 3644 3276 3658
rect 3242 3576 3276 3586
rect 3242 3508 3276 3514
rect 3242 3440 3276 3442
rect 3242 3404 3276 3406
rect 3242 3332 3276 3338
rect 3242 3260 3276 3270
rect 3242 3188 3276 3202
rect 3242 3116 3276 3134
rect 3242 3044 3276 3066
rect 3242 2972 3276 2998
rect 3242 2900 3276 2930
rect 3242 2828 3276 2862
rect 3242 2760 3276 2794
rect 3242 2692 3276 2722
rect 3242 2624 3276 2650
rect 3242 2556 3276 2578
rect 3242 2488 3276 2506
rect 3242 2420 3276 2434
rect 3242 2352 3276 2362
rect 3242 2284 3276 2290
rect 3242 2216 3276 2218
rect 3242 2180 3276 2182
rect 3242 2108 3276 2114
rect 3242 2036 3276 2046
rect 3242 1964 3276 1978
rect 3242 1892 3276 1910
rect 3242 1807 3276 1842
rect 3550 3780 3598 3823
rect 3550 3778 3558 3780
rect 3400 3712 3434 3730
rect 3400 3644 3434 3658
rect 3400 3576 3434 3586
rect 3400 3508 3434 3514
rect 3400 3440 3434 3442
rect 3400 3404 3434 3406
rect 3400 3332 3434 3338
rect 3400 3260 3434 3270
rect 3400 3188 3434 3202
rect 3400 3116 3434 3134
rect 3400 3044 3434 3066
rect 3400 2972 3434 2998
rect 3400 2900 3434 2930
rect 3400 2828 3434 2862
rect 3400 2760 3434 2794
rect 3400 2692 3434 2722
rect 3400 2624 3434 2650
rect 3400 2556 3434 2578
rect 3400 2488 3434 2506
rect 3400 2420 3434 2434
rect 3400 2352 3434 2362
rect 3400 2284 3434 2290
rect 3400 2216 3434 2218
rect 3400 2180 3434 2182
rect 3400 2108 3434 2114
rect 3400 2036 3434 2046
rect 3400 1964 3434 1978
rect 3400 1892 3434 1910
rect 3400 1807 3434 1842
rect 3592 3778 3598 3780
rect 3558 3712 3592 3730
rect 3558 3644 3592 3658
rect 3558 3576 3592 3586
rect 3558 3508 3592 3514
rect 3558 3440 3592 3442
rect 3558 3404 3592 3406
rect 3558 3332 3592 3338
rect 3558 3260 3592 3270
rect 3558 3188 3592 3202
rect 3558 3116 3592 3134
rect 3558 3044 3592 3066
rect 3558 2972 3592 2998
rect 3558 2900 3592 2930
rect 3558 2828 3592 2862
rect 3558 2760 3592 2794
rect 3558 2692 3592 2722
rect 3558 2624 3592 2650
rect 3558 2556 3592 2578
rect 3558 2488 3592 2506
rect 3558 2420 3592 2434
rect 3558 2352 3592 2362
rect 3558 2284 3592 2290
rect 3558 2216 3592 2218
rect 3558 2180 3592 2182
rect 3558 2108 3592 2114
rect 3558 2036 3592 2046
rect 3558 1964 3592 1978
rect 3558 1892 3592 1910
rect 3558 1807 3592 1842
rect 2972 1730 3005 1764
rect 3039 1730 3072 1764
rect 3130 1730 3163 1764
rect 3197 1730 3230 1764
rect 3288 1730 3321 1764
rect 3355 1730 3388 1764
rect 3446 1730 3479 1764
rect 3513 1730 3546 1764
rect 2834 1668 3662 1676
rect 2834 1665 3620 1668
rect 2730 1662 3620 1665
rect 2730 1628 2733 1662
rect 2767 1634 3620 1662
rect 3654 1634 3662 1668
rect 2767 1628 3662 1634
rect 2730 1627 3662 1628
rect 2730 1625 2873 1627
rect 1900 1154 1934 1180
rect 1900 1086 1934 1108
rect 1900 1018 1934 1036
rect 1900 937 1934 964
rect 2114 1203 2694 1246
rect 2807 1558 2850 1563
rect 2807 1524 2811 1558
rect 2845 1524 2850 1558
rect 1312 844 1878 853
rect 1312 810 1836 844
rect 1870 810 1878 844
rect 1312 804 1878 810
rect 1111 725 1145 759
rect 1387 718 1421 726
rect 1111 657 1145 687
rect 1379 710 1429 718
rect 1379 676 1387 710
rect 1421 676 1429 710
rect 1379 668 1429 676
rect 1485 691 1519 708
rect 1387 660 1421 668
rect 1111 589 1145 615
rect 1111 521 1145 543
rect 1111 453 1145 471
rect 1111 372 1145 399
rect 1485 623 1519 631
rect 1485 555 1519 559
rect 1485 449 1519 453
rect 1485 377 1519 385
rect 1485 300 1519 317
rect 1643 691 1677 708
rect 1643 623 1677 631
rect 1643 555 1677 559
rect 1643 449 1677 453
rect 1643 377 1677 385
rect 1643 300 1677 317
rect 1881 691 1915 708
rect 1881 623 1915 631
rect 1881 555 1915 559
rect 1881 449 1915 453
rect 1881 377 1915 385
rect 1881 300 1915 317
rect 2039 691 2073 708
rect 2039 623 2073 631
rect 2039 555 2073 559
rect 2039 449 2073 453
rect 2039 377 2073 385
rect 2039 300 2073 317
rect 876 244 1073 246
rect 765 243 1073 244
rect 765 209 1036 243
rect 1070 209 1086 243
rect 2114 226 2157 1203
rect 2208 771 2260 774
rect 2296 771 2330 784
rect 2208 768 2333 771
rect 2208 734 2296 768
rect 2330 734 2333 768
rect 2208 732 2333 734
rect 2208 594 2260 732
rect 2296 718 2330 732
rect 2807 713 2850 1524
rect 2977 1516 3010 1550
rect 3044 1516 3077 1550
rect 3135 1516 3168 1550
rect 3202 1516 3235 1550
rect 3293 1516 3326 1550
rect 3360 1516 3393 1550
rect 3451 1516 3484 1550
rect 3518 1516 3551 1550
rect 2373 708 2850 713
rect 2373 674 2377 708
rect 2411 674 2850 708
rect 2373 670 2850 674
rect 2931 1439 2965 1482
rect 2931 1371 2965 1401
rect 2931 1303 2965 1329
rect 2931 1235 2965 1257
rect 2931 1167 2965 1185
rect 2931 1099 2965 1113
rect 2931 1031 2965 1041
rect 2931 963 2965 969
rect 2931 895 2965 897
rect 2931 859 2965 861
rect 2931 787 2965 793
rect 2931 715 2965 725
rect 2350 594 2384 595
rect 2208 578 2389 594
rect 2208 542 2350 578
rect 2384 542 2389 578
rect 2508 578 2542 595
rect 2350 510 2384 518
rect 2350 442 2384 446
rect 2350 336 2384 340
rect 2350 264 2384 272
rect 765 207 1073 209
rect 1367 208 1401 224
rect 876 206 1073 207
rect 1331 174 1367 208
rect 1367 158 1401 174
rect 2114 208 2186 226
rect 2114 174 2129 208
rect 2163 174 2186 208
rect 2350 187 2384 204
rect 2665 578 2708 670
rect 2665 535 2666 578
rect 2508 510 2542 518
rect 2508 442 2542 446
rect 2508 336 2542 340
rect 2508 264 2542 272
rect 2508 187 2542 204
rect 2700 535 2708 578
rect 2931 643 2965 657
rect 2931 571 2965 589
rect 2666 510 2700 518
rect 2666 442 2700 446
rect 2931 499 2965 521
rect 2931 427 2965 453
rect 2931 355 2965 385
rect 2666 336 2700 340
rect 2666 264 2700 272
rect 2666 187 2700 204
rect 2805 347 2845 350
rect 2805 313 2808 347
rect 2842 313 2845 347
rect 2114 164 2186 174
rect -692 157 66 158
rect 2117 157 2186 164
rect 2805 177 2845 313
rect 3089 1439 3123 1482
rect 3089 1371 3123 1401
rect 3089 1303 3123 1329
rect 3089 1235 3123 1257
rect 3089 1167 3123 1185
rect 3089 1099 3123 1113
rect 3089 1031 3123 1041
rect 3089 963 3123 969
rect 3089 895 3123 897
rect 3089 859 3123 861
rect 3089 787 3123 793
rect 3089 715 3123 725
rect 3089 643 3123 657
rect 3089 571 3123 589
rect 3089 499 3123 521
rect 3089 427 3123 453
rect 3089 355 3123 385
rect 2931 274 2965 317
rect 3084 317 3089 322
rect 3247 1439 3281 1482
rect 3247 1371 3281 1401
rect 3247 1303 3281 1329
rect 3247 1235 3281 1257
rect 3247 1167 3281 1185
rect 3247 1099 3281 1113
rect 3247 1031 3281 1041
rect 3247 963 3281 969
rect 3247 895 3281 897
rect 3247 859 3281 861
rect 3247 787 3281 793
rect 3247 715 3281 725
rect 3247 643 3281 657
rect 3247 571 3281 589
rect 3247 499 3281 521
rect 3247 427 3281 453
rect 3247 355 3281 385
rect 3123 317 3124 322
rect 3084 177 3124 317
rect 3247 274 3281 317
rect 3405 1439 3439 1482
rect 3405 1371 3439 1401
rect 3405 1303 3439 1329
rect 3405 1235 3439 1257
rect 3405 1167 3439 1185
rect 3405 1099 3439 1113
rect 3405 1031 3439 1041
rect 3405 963 3439 969
rect 3405 895 3439 897
rect 3405 859 3439 861
rect 3405 787 3439 793
rect 3405 715 3439 725
rect 3405 643 3439 657
rect 3405 571 3439 589
rect 3405 499 3439 521
rect 3405 427 3439 453
rect 3405 355 3439 385
rect 3405 313 3439 317
rect 3563 1439 3597 1482
rect 3563 1371 3597 1401
rect 3563 1303 3597 1329
rect 3563 1235 3597 1257
rect 3563 1167 3597 1185
rect 3563 1099 3597 1113
rect 3563 1031 3597 1041
rect 3563 963 3597 969
rect 3563 895 3597 897
rect 3563 859 3597 861
rect 3563 787 3597 793
rect 3563 715 3597 725
rect 3563 643 3597 657
rect 3563 571 3597 589
rect 3563 499 3597 521
rect 3563 427 3597 453
rect 3563 355 3597 385
rect 3402 177 3442 313
rect 3563 274 3597 317
rect -692 110 1251 157
rect 2805 137 3442 177
rect -692 76 -596 110
rect -562 99 1251 110
rect -561 95 757 99
rect -561 93 72 95
rect -692 65 -595 76
rect -561 65 -398 93
rect -692 59 -398 65
rect -364 89 -167 93
rect -364 59 -271 89
rect -692 55 -271 59
rect -237 59 -167 89
rect -133 85 72 93
rect -133 59 -49 85
rect -237 55 -49 59
rect -692 51 -49 55
rect -15 61 72 85
rect 106 93 578 95
rect 106 61 116 93
rect -15 59 116 61
rect 150 59 240 93
rect 274 59 305 93
rect 339 59 409 93
rect 443 59 479 93
rect 513 61 578 93
rect 612 93 757 95
rect 612 61 662 93
rect 513 59 662 61
rect 696 65 757 93
rect 791 93 944 99
rect 791 65 849 93
rect 696 59 849 65
rect 883 65 944 93
rect 978 97 1251 99
rect 978 93 1145 97
rect 978 65 1052 93
rect 883 59 1052 65
rect 1086 63 1145 93
rect 1179 63 1251 97
rect 1086 59 1251 63
rect -15 51 1251 59
rect -692 0 1251 51
rect -692 -4 66 0
<< viali >>
rect -142 3826 -140 3858
rect -140 3826 -108 3858
rect -142 3824 -108 3826
rect 779 3793 813 3813
rect 779 3779 813 3793
rect 779 3725 813 3741
rect 779 3707 813 3725
rect 779 3657 813 3669
rect 779 3635 813 3657
rect 779 3589 813 3597
rect 779 3563 813 3589
rect 779 3521 813 3525
rect 779 3491 813 3521
rect 779 3419 813 3453
rect 779 3351 813 3381
rect 779 3347 813 3351
rect 779 3283 813 3309
rect 779 3275 813 3283
rect 779 3215 813 3237
rect 779 3203 813 3215
rect 779 3147 813 3165
rect 779 3131 813 3147
rect 779 3079 813 3093
rect 779 3059 813 3079
rect 937 3793 971 3813
rect 937 3779 971 3793
rect 937 3725 971 3741
rect 937 3707 971 3725
rect 937 3657 971 3669
rect 937 3635 971 3657
rect 937 3589 971 3597
rect 937 3563 971 3589
rect 937 3521 971 3525
rect 937 3491 971 3521
rect 937 3419 971 3453
rect 937 3351 971 3381
rect 937 3347 971 3351
rect 937 3283 971 3309
rect 937 3275 971 3283
rect 937 3215 971 3237
rect 937 3203 971 3215
rect 937 3147 971 3165
rect 937 3131 971 3147
rect 937 3079 971 3093
rect 937 3059 971 3079
rect 1095 3793 1129 3813
rect 1095 3779 1129 3793
rect 1095 3725 1129 3741
rect 1095 3707 1129 3725
rect 1353 3802 1387 3836
rect 1577 3797 1611 3831
rect 1820 3794 1854 3828
rect 2043 3796 2077 3830
rect 2115 3796 2149 3830
rect 2278 3794 2312 3828
rect 2350 3797 2379 3828
rect 2379 3797 2384 3828
rect 2537 3799 2571 3833
rect 2609 3831 2643 3833
rect 2609 3799 2618 3831
rect 2618 3799 2643 3831
rect 2350 3794 2384 3797
rect 2926 3882 2960 3916
rect 2926 3746 2960 3764
rect 2926 3730 2960 3746
rect 1095 3657 1129 3669
rect 1095 3635 1129 3657
rect 1095 3589 1129 3597
rect 2926 3678 2960 3692
rect 2926 3658 2960 3678
rect 2926 3610 2960 3620
rect 1095 3563 1129 3589
rect 2180 3545 2214 3565
rect 1095 3521 1129 3525
rect 1095 3491 1129 3521
rect 1095 3419 1129 3453
rect 1095 3351 1129 3381
rect 1095 3347 1129 3351
rect 1095 3283 1129 3309
rect 1095 3275 1129 3283
rect 1095 3215 1129 3237
rect 1095 3203 1129 3215
rect 1095 3147 1129 3165
rect 1095 3131 1129 3147
rect 1403 3493 1437 3501
rect 1403 3467 1437 3493
rect 1403 3425 1437 3429
rect 1403 3395 1437 3425
rect 1403 3323 1437 3357
rect 1403 3255 1437 3285
rect 1403 3251 1437 3255
rect 1403 3187 1437 3213
rect 1403 3179 1437 3187
rect 1561 3493 1595 3501
rect 1561 3467 1595 3493
rect 1561 3425 1595 3429
rect 1561 3395 1595 3425
rect 1561 3323 1595 3357
rect 1561 3255 1595 3285
rect 1561 3251 1595 3255
rect 1561 3187 1595 3213
rect 1561 3179 1595 3187
rect 2180 3531 2214 3545
rect 2180 3477 2214 3493
rect 2180 3459 2214 3477
rect 2180 3409 2214 3421
rect 2180 3387 2214 3409
rect 2180 3341 2214 3349
rect 2180 3315 2214 3341
rect 2180 3273 2214 3277
rect 2180 3243 2214 3273
rect 2180 3171 2214 3205
rect 1095 3079 1129 3093
rect 1240 3084 1274 3118
rect 2180 3103 2214 3133
rect 2180 3099 2214 3103
rect 1095 3059 1129 3079
rect 1002 2900 1036 2934
rect 2180 3035 2214 3061
rect 2180 3027 2214 3035
rect 1404 2964 1438 2984
rect 1404 2950 1438 2964
rect 1404 2896 1438 2912
rect 1404 2878 1438 2896
rect 1404 2828 1438 2840
rect 1404 2806 1438 2828
rect 879 2655 913 2663
rect 879 2629 913 2655
rect 879 2587 913 2591
rect 879 2557 913 2587
rect 879 2485 913 2519
rect 1404 2760 1438 2768
rect 1404 2734 1438 2760
rect 1037 2655 1071 2663
rect 1037 2629 1071 2655
rect 1037 2587 1071 2591
rect 1037 2557 1071 2587
rect 879 2417 913 2447
rect 879 2413 913 2417
rect 879 2349 913 2375
rect 879 2341 913 2349
rect 1037 2485 1071 2519
rect 1037 2417 1071 2447
rect 1037 2413 1071 2417
rect 1037 2349 1071 2375
rect 1037 2341 1071 2349
rect 1404 2692 1438 2696
rect 1404 2662 1438 2692
rect 1404 2590 1438 2624
rect 1404 2522 1438 2552
rect 1404 2518 1438 2522
rect 1404 2454 1438 2480
rect 1404 2446 1438 2454
rect 1404 2386 1438 2408
rect 1404 2374 1438 2386
rect 1404 2318 1438 2336
rect 1404 2302 1438 2318
rect 1404 2250 1438 2264
rect 1404 2230 1438 2250
rect 1562 2964 1596 2984
rect 1562 2950 1596 2964
rect 1562 2896 1596 2912
rect 1562 2878 1596 2896
rect 1562 2828 1596 2840
rect 1562 2806 1596 2828
rect 1562 2760 1596 2768
rect 1562 2734 1596 2760
rect 1562 2692 1596 2696
rect 1562 2662 1596 2692
rect 1562 2590 1596 2624
rect 1562 2522 1596 2552
rect 1562 2518 1596 2522
rect 1562 2454 1596 2480
rect 1562 2446 1596 2454
rect 1562 2386 1596 2408
rect 1562 2374 1596 2386
rect 1562 2318 1596 2336
rect 1562 2302 1596 2318
rect 1562 2250 1596 2264
rect 1562 2230 1596 2250
rect 1720 2964 1754 2984
rect 1720 2950 1754 2964
rect 1720 2896 1754 2912
rect 1720 2878 1754 2896
rect 2180 2967 2214 2989
rect 2180 2955 2214 2967
rect 2180 2899 2214 2917
rect 2180 2883 2214 2899
rect 2338 3545 2372 3565
rect 2338 3531 2372 3545
rect 2338 3477 2372 3493
rect 2338 3459 2372 3477
rect 2338 3409 2372 3421
rect 2338 3387 2372 3409
rect 2338 3341 2372 3349
rect 2338 3315 2372 3341
rect 2338 3273 2372 3277
rect 2338 3243 2372 3273
rect 2338 3171 2372 3205
rect 2338 3103 2372 3133
rect 2338 3099 2372 3103
rect 2338 3035 2372 3061
rect 2338 3027 2372 3035
rect 2338 2967 2372 2989
rect 2338 2955 2372 2967
rect 2338 2899 2372 2917
rect 2338 2883 2372 2899
rect 1720 2828 1754 2840
rect 1720 2806 1754 2828
rect 1720 2760 1754 2768
rect 1720 2734 1754 2760
rect 1720 2692 1754 2696
rect 1720 2662 1754 2692
rect 1720 2590 1754 2624
rect 2180 2831 2214 2845
rect 2180 2811 2214 2831
rect 2338 2831 2372 2845
rect 2338 2811 2372 2831
rect 2496 3545 2530 3565
rect 2496 3531 2530 3545
rect 2496 3477 2530 3493
rect 2496 3459 2530 3477
rect 2496 3409 2530 3421
rect 2496 3387 2530 3409
rect 2496 3341 2530 3349
rect 2496 3315 2530 3341
rect 2496 3273 2530 3277
rect 2496 3243 2530 3273
rect 2496 3171 2530 3205
rect 2496 3103 2530 3133
rect 2496 3099 2530 3103
rect 2496 3035 2530 3061
rect 2496 3027 2530 3035
rect 2496 2967 2530 2989
rect 2496 2955 2530 2967
rect 2496 2899 2530 2917
rect 2496 2883 2530 2899
rect 2496 2831 2530 2845
rect 2496 2811 2530 2831
rect 2926 3586 2960 3610
rect 2926 3542 2960 3548
rect 2926 3514 2960 3542
rect 2926 3474 2960 3476
rect 2926 3442 2960 3474
rect 2926 3372 2960 3404
rect 2926 3370 2960 3372
rect 2926 3304 2960 3332
rect 2926 3298 2960 3304
rect 2926 3236 2960 3260
rect 2926 3226 2960 3236
rect 2926 3168 2960 3188
rect 2926 3154 2960 3168
rect 2926 3100 2960 3116
rect 2926 3082 2960 3100
rect 2926 3032 2960 3044
rect 2926 3010 2960 3032
rect 2926 2964 2960 2972
rect 2926 2938 2960 2964
rect 2926 2896 2960 2900
rect 2926 2866 2960 2896
rect 2926 2794 2960 2828
rect 2926 2726 2960 2756
rect 2926 2722 2960 2726
rect 2926 2658 2960 2684
rect 2618 2611 2652 2645
rect 1720 2522 1754 2552
rect 1720 2518 1754 2522
rect 1720 2454 1754 2480
rect 1720 2446 1754 2454
rect 1720 2386 1754 2408
rect 1720 2374 1754 2386
rect 1720 2318 1754 2336
rect 1720 2302 1754 2318
rect 2123 2443 2157 2451
rect 2123 2417 2157 2443
rect 2123 2375 2157 2379
rect 2123 2345 2157 2375
rect 1720 2250 1754 2264
rect 1720 2230 1754 2250
rect 123 1306 157 1340
rect 165 956 199 990
rect 530 956 564 990
rect 627 677 661 711
rect 682 306 716 340
rect 1417 1922 1451 1956
rect 2123 2273 2157 2307
rect 2123 2205 2157 2235
rect 2123 2201 2157 2205
rect 2123 2137 2157 2163
rect 2123 2129 2157 2137
rect 2281 2443 2315 2451
rect 2281 2417 2315 2443
rect 2281 2375 2315 2379
rect 2281 2345 2315 2375
rect 2281 2273 2315 2307
rect 2281 2205 2315 2235
rect 2281 2201 2315 2205
rect 2281 2137 2315 2163
rect 2281 2129 2315 2137
rect 2400 2447 2434 2455
rect 2400 2421 2434 2447
rect 2400 2379 2434 2383
rect 2400 2349 2434 2379
rect 2400 2277 2434 2311
rect 2400 2209 2434 2239
rect 2400 2205 2434 2209
rect 2400 2141 2434 2167
rect 2400 2133 2434 2141
rect 2558 2447 2592 2455
rect 2558 2421 2592 2447
rect 2558 2379 2592 2383
rect 2558 2349 2592 2379
rect 2742 2328 2776 2362
rect 2926 2650 2960 2658
rect 2926 2590 2960 2612
rect 2926 2578 2960 2590
rect 2926 2522 2960 2540
rect 2926 2506 2960 2522
rect 2926 2454 2960 2468
rect 2926 2434 2960 2454
rect 2926 2386 2960 2396
rect 2926 2362 2960 2386
rect 2558 2277 2592 2311
rect 2558 2209 2592 2239
rect 2558 2205 2592 2209
rect 2558 2141 2592 2167
rect 2558 2133 2592 2141
rect 2926 2318 2960 2324
rect 2926 2290 2960 2318
rect 2926 2250 2960 2252
rect 2926 2218 2960 2250
rect 2926 2148 2960 2180
rect 2926 2146 2960 2148
rect 2926 2080 2960 2108
rect 2926 2074 2960 2080
rect 2521 1965 2555 1999
rect 2926 2012 2960 2036
rect 2926 2002 2960 2012
rect 2926 1944 2960 1964
rect 2926 1930 2960 1944
rect 949 1674 983 1682
rect 949 1648 983 1674
rect 949 1606 983 1610
rect 949 1576 983 1606
rect 949 1504 983 1538
rect 949 1436 983 1466
rect 949 1432 983 1436
rect 949 1368 983 1394
rect 949 1360 983 1368
rect 1107 1674 1141 1682
rect 1107 1648 1141 1674
rect 1107 1606 1141 1610
rect 1107 1576 1141 1606
rect 1107 1504 1141 1538
rect 1107 1436 1141 1466
rect 1107 1432 1141 1436
rect 1107 1368 1141 1394
rect 1107 1360 1141 1368
rect 1265 1674 1299 1682
rect 1265 1648 1299 1674
rect 1265 1606 1299 1610
rect 1265 1576 1299 1606
rect 1265 1504 1299 1538
rect 1265 1436 1299 1466
rect 1265 1432 1299 1436
rect 2841 1877 2875 1911
rect 1368 1409 1402 1443
rect 1584 1698 1618 1718
rect 1584 1684 1618 1698
rect 1584 1630 1618 1646
rect 1584 1612 1618 1630
rect 1584 1562 1618 1574
rect 1584 1540 1618 1562
rect 1584 1494 1618 1502
rect 1584 1468 1618 1494
rect 1584 1426 1618 1430
rect 1265 1368 1299 1394
rect 1265 1360 1299 1368
rect 1584 1396 1618 1426
rect 1584 1324 1618 1358
rect 1584 1256 1618 1286
rect 1584 1252 1618 1256
rect 953 1133 987 1153
rect 953 1119 987 1133
rect 953 1065 987 1081
rect 953 1047 987 1065
rect 953 997 987 1009
rect 953 975 987 997
rect 953 929 987 937
rect 953 903 987 929
rect 953 861 987 865
rect 953 831 987 861
rect 953 759 987 793
rect 953 691 987 721
rect 953 687 987 691
rect 953 623 987 649
rect 953 615 987 623
rect 953 555 987 577
rect 953 543 987 555
rect 953 487 987 505
rect 953 471 987 487
rect 953 419 987 433
rect 953 399 987 419
rect 1111 1133 1145 1153
rect 1111 1119 1145 1133
rect 1111 1065 1145 1081
rect 1111 1047 1145 1065
rect 1111 997 1145 1009
rect 1111 975 1145 997
rect 1111 929 1145 937
rect 1111 903 1145 929
rect 1111 861 1145 865
rect 1111 831 1145 861
rect 1319 1152 1353 1186
rect 1584 1188 1618 1214
rect 1584 1180 1618 1188
rect 1584 1120 1618 1142
rect 1584 1108 1618 1120
rect 1584 1052 1618 1070
rect 1584 1036 1618 1052
rect 1584 984 1618 998
rect 1584 964 1618 984
rect 1742 1698 1776 1718
rect 1742 1684 1776 1698
rect 1742 1630 1776 1646
rect 1742 1612 1776 1630
rect 1742 1562 1776 1574
rect 1742 1540 1776 1562
rect 1742 1494 1776 1502
rect 1742 1468 1776 1494
rect 1742 1426 1776 1430
rect 1742 1396 1776 1426
rect 1742 1324 1776 1358
rect 1742 1256 1776 1286
rect 1742 1252 1776 1256
rect 1742 1188 1776 1214
rect 1742 1180 1776 1188
rect 1742 1120 1776 1142
rect 1742 1108 1776 1120
rect 1742 1052 1776 1070
rect 1742 1036 1776 1052
rect 1742 984 1776 998
rect 1742 964 1776 984
rect 1900 1698 1934 1718
rect 1900 1684 1934 1698
rect 1900 1630 1934 1646
rect 1900 1612 1934 1630
rect 1900 1562 1934 1574
rect 1900 1540 1934 1562
rect 1900 1494 1934 1502
rect 1900 1468 1934 1494
rect 1900 1426 1934 1430
rect 1900 1396 1934 1426
rect 1900 1324 1934 1358
rect 1900 1256 1934 1286
rect 2193 1642 2227 1650
rect 2193 1616 2227 1642
rect 2193 1574 2227 1578
rect 2193 1544 2227 1574
rect 2193 1472 2227 1506
rect 2193 1404 2227 1434
rect 2193 1400 2227 1404
rect 2193 1336 2227 1362
rect 2193 1328 2227 1336
rect 2351 1642 2385 1650
rect 2351 1616 2385 1642
rect 2351 1574 2385 1578
rect 2351 1544 2385 1574
rect 2351 1472 2385 1506
rect 2351 1404 2385 1434
rect 2351 1400 2385 1404
rect 2351 1336 2385 1362
rect 2351 1328 2385 1336
rect 2509 1642 2543 1650
rect 2509 1616 2543 1642
rect 2509 1574 2543 1578
rect 2509 1544 2543 1574
rect 2509 1472 2543 1506
rect 2509 1404 2543 1434
rect 2509 1400 2543 1404
rect 2509 1336 2543 1362
rect 2509 1328 2543 1336
rect 1900 1252 1934 1256
rect 2926 1876 2960 1892
rect 2926 1858 2960 1876
rect 3084 3746 3118 3764
rect 3084 3730 3118 3746
rect 3084 3678 3118 3692
rect 3084 3658 3118 3678
rect 3084 3610 3118 3620
rect 3084 3586 3118 3610
rect 3084 3542 3118 3548
rect 3084 3514 3118 3542
rect 3084 3474 3118 3476
rect 3084 3442 3118 3474
rect 3084 3372 3118 3404
rect 3084 3370 3118 3372
rect 3084 3304 3118 3332
rect 3084 3298 3118 3304
rect 3084 3236 3118 3260
rect 3084 3226 3118 3236
rect 3084 3168 3118 3188
rect 3084 3154 3118 3168
rect 3084 3100 3118 3116
rect 3084 3082 3118 3100
rect 3084 3032 3118 3044
rect 3084 3010 3118 3032
rect 3084 2964 3118 2972
rect 3084 2938 3118 2964
rect 3084 2896 3118 2900
rect 3084 2866 3118 2896
rect 3084 2794 3118 2828
rect 3084 2726 3118 2756
rect 3084 2722 3118 2726
rect 3084 2658 3118 2684
rect 3084 2650 3118 2658
rect 3084 2590 3118 2612
rect 3084 2578 3118 2590
rect 3084 2522 3118 2540
rect 3084 2506 3118 2522
rect 3084 2454 3118 2468
rect 3084 2434 3118 2454
rect 3084 2386 3118 2396
rect 3084 2362 3118 2386
rect 3084 2318 3118 2324
rect 3084 2290 3118 2318
rect 3084 2250 3118 2252
rect 3084 2218 3118 2250
rect 3084 2148 3118 2180
rect 3084 2146 3118 2148
rect 3084 2080 3118 2108
rect 3084 2074 3118 2080
rect 3084 2012 3118 2036
rect 3084 2002 3118 2012
rect 3084 1944 3118 1964
rect 3084 1930 3118 1944
rect 3084 1876 3118 1892
rect 3084 1858 3118 1876
rect 3242 3746 3276 3764
rect 3242 3730 3276 3746
rect 3242 3678 3276 3692
rect 3242 3658 3276 3678
rect 3242 3610 3276 3620
rect 3242 3586 3276 3610
rect 3242 3542 3276 3548
rect 3242 3514 3276 3542
rect 3242 3474 3276 3476
rect 3242 3442 3276 3474
rect 3242 3372 3276 3404
rect 3242 3370 3276 3372
rect 3242 3304 3276 3332
rect 3242 3298 3276 3304
rect 3242 3236 3276 3260
rect 3242 3226 3276 3236
rect 3242 3168 3276 3188
rect 3242 3154 3276 3168
rect 3242 3100 3276 3116
rect 3242 3082 3276 3100
rect 3242 3032 3276 3044
rect 3242 3010 3276 3032
rect 3242 2964 3276 2972
rect 3242 2938 3276 2964
rect 3242 2896 3276 2900
rect 3242 2866 3276 2896
rect 3242 2794 3276 2828
rect 3242 2726 3276 2756
rect 3242 2722 3276 2726
rect 3242 2658 3276 2684
rect 3242 2650 3276 2658
rect 3242 2590 3276 2612
rect 3242 2578 3276 2590
rect 3242 2522 3276 2540
rect 3242 2506 3276 2522
rect 3242 2454 3276 2468
rect 3242 2434 3276 2454
rect 3242 2386 3276 2396
rect 3242 2362 3276 2386
rect 3242 2318 3276 2324
rect 3242 2290 3276 2318
rect 3242 2250 3276 2252
rect 3242 2218 3276 2250
rect 3242 2148 3276 2180
rect 3242 2146 3276 2148
rect 3242 2080 3276 2108
rect 3242 2074 3276 2080
rect 3242 2012 3276 2036
rect 3242 2002 3276 2012
rect 3242 1944 3276 1964
rect 3242 1930 3276 1944
rect 3242 1876 3276 1892
rect 3242 1858 3276 1876
rect 3400 3746 3434 3764
rect 3400 3730 3434 3746
rect 3400 3678 3434 3692
rect 3400 3658 3434 3678
rect 3400 3610 3434 3620
rect 3400 3586 3434 3610
rect 3400 3542 3434 3548
rect 3400 3514 3434 3542
rect 3400 3474 3434 3476
rect 3400 3442 3434 3474
rect 3400 3372 3434 3404
rect 3400 3370 3434 3372
rect 3400 3304 3434 3332
rect 3400 3298 3434 3304
rect 3400 3236 3434 3260
rect 3400 3226 3434 3236
rect 3400 3168 3434 3188
rect 3400 3154 3434 3168
rect 3400 3100 3434 3116
rect 3400 3082 3434 3100
rect 3400 3032 3434 3044
rect 3400 3010 3434 3032
rect 3400 2964 3434 2972
rect 3400 2938 3434 2964
rect 3400 2896 3434 2900
rect 3400 2866 3434 2896
rect 3400 2794 3434 2828
rect 3400 2726 3434 2756
rect 3400 2722 3434 2726
rect 3400 2658 3434 2684
rect 3400 2650 3434 2658
rect 3400 2590 3434 2612
rect 3400 2578 3434 2590
rect 3400 2522 3434 2540
rect 3400 2506 3434 2522
rect 3400 2454 3434 2468
rect 3400 2434 3434 2454
rect 3400 2386 3434 2396
rect 3400 2362 3434 2386
rect 3400 2318 3434 2324
rect 3400 2290 3434 2318
rect 3400 2250 3434 2252
rect 3400 2218 3434 2250
rect 3400 2148 3434 2180
rect 3400 2146 3434 2148
rect 3400 2080 3434 2108
rect 3400 2074 3434 2080
rect 3400 2012 3434 2036
rect 3400 2002 3434 2012
rect 3400 1944 3434 1964
rect 3400 1930 3434 1944
rect 3400 1876 3434 1892
rect 3400 1858 3434 1876
rect 3558 3746 3592 3764
rect 3558 3730 3592 3746
rect 3558 3678 3592 3692
rect 3558 3658 3592 3678
rect 3558 3610 3592 3620
rect 3558 3586 3592 3610
rect 3558 3542 3592 3548
rect 3558 3514 3592 3542
rect 3558 3474 3592 3476
rect 3558 3442 3592 3474
rect 3558 3372 3592 3404
rect 3558 3370 3592 3372
rect 3558 3304 3592 3332
rect 3558 3298 3592 3304
rect 3558 3236 3592 3260
rect 3558 3226 3592 3236
rect 3558 3168 3592 3188
rect 3558 3154 3592 3168
rect 3558 3100 3592 3116
rect 3558 3082 3592 3100
rect 3558 3032 3592 3044
rect 3558 3010 3592 3032
rect 3558 2964 3592 2972
rect 3558 2938 3592 2964
rect 3558 2896 3592 2900
rect 3558 2866 3592 2896
rect 3558 2794 3592 2828
rect 3558 2726 3592 2756
rect 3558 2722 3592 2726
rect 3558 2658 3592 2684
rect 3558 2650 3592 2658
rect 3558 2590 3592 2612
rect 3558 2578 3592 2590
rect 3558 2522 3592 2540
rect 3558 2506 3592 2522
rect 3558 2454 3592 2468
rect 3558 2434 3592 2454
rect 3558 2386 3592 2396
rect 3558 2362 3592 2386
rect 3558 2318 3592 2324
rect 3558 2290 3592 2318
rect 3558 2250 3592 2252
rect 3558 2218 3592 2250
rect 3558 2148 3592 2180
rect 3558 2146 3592 2148
rect 3558 2080 3592 2108
rect 3558 2074 3592 2080
rect 3558 2012 3592 2036
rect 3558 2002 3592 2012
rect 3558 1944 3592 1964
rect 3558 1930 3592 1944
rect 3558 1876 3592 1892
rect 3558 1858 3592 1876
rect 3005 1730 3039 1764
rect 3163 1730 3197 1764
rect 3321 1730 3355 1764
rect 3479 1730 3513 1764
rect 2733 1628 2767 1662
rect 3620 1634 3654 1668
rect 1900 1188 1934 1214
rect 1900 1180 1934 1188
rect 1900 1120 1934 1142
rect 1900 1108 1934 1120
rect 1900 1052 1934 1070
rect 1900 1036 1934 1052
rect 1900 984 1934 998
rect 1900 964 1934 984
rect 2811 1524 2845 1558
rect 1836 810 1870 844
rect 1111 759 1145 793
rect 1111 691 1145 721
rect 1111 687 1145 691
rect 1387 676 1421 710
rect 1111 623 1145 649
rect 1111 615 1145 623
rect 1111 555 1145 577
rect 1111 543 1145 555
rect 1111 487 1145 505
rect 1111 471 1145 487
rect 1111 419 1145 433
rect 1111 399 1145 419
rect 1485 657 1519 665
rect 1485 631 1519 657
rect 1485 589 1519 593
rect 1485 559 1519 589
rect 1485 487 1519 521
rect 1485 419 1519 449
rect 1485 415 1519 419
rect 1485 351 1519 377
rect 1485 343 1519 351
rect 1643 657 1677 665
rect 1643 631 1677 657
rect 1643 589 1677 593
rect 1643 559 1677 589
rect 1643 487 1677 521
rect 1643 419 1677 449
rect 1643 415 1677 419
rect 1643 351 1677 377
rect 1643 343 1677 351
rect 1881 657 1915 665
rect 1881 631 1915 657
rect 1881 589 1915 593
rect 1881 559 1915 589
rect 1881 487 1915 521
rect 1881 419 1915 449
rect 1881 415 1915 419
rect 1881 351 1915 377
rect 1881 343 1915 351
rect 2039 657 2073 665
rect 2039 631 2073 657
rect 2039 589 2073 593
rect 2039 559 2073 589
rect 2039 487 2073 521
rect 2039 419 2073 449
rect 2039 415 2073 419
rect 2039 351 2073 377
rect 2039 343 2073 351
rect 3010 1516 3044 1550
rect 3168 1516 3202 1550
rect 3326 1516 3360 1550
rect 3484 1516 3518 1550
rect 2377 674 2411 708
rect 2931 1405 2965 1435
rect 2931 1401 2965 1405
rect 2931 1337 2965 1363
rect 2931 1329 2965 1337
rect 2931 1269 2965 1291
rect 2931 1257 2965 1269
rect 2931 1201 2965 1219
rect 2931 1185 2965 1201
rect 2931 1133 2965 1147
rect 2931 1113 2965 1133
rect 2931 1065 2965 1075
rect 2931 1041 2965 1065
rect 2931 997 2965 1003
rect 2931 969 2965 997
rect 2931 929 2965 931
rect 2931 897 2965 929
rect 2931 827 2965 859
rect 2931 825 2965 827
rect 2931 759 2965 787
rect 2931 753 2965 759
rect 2931 691 2965 715
rect 2931 681 2965 691
rect 2350 544 2384 552
rect 2350 518 2384 544
rect 2508 544 2542 552
rect 2350 476 2384 480
rect 2350 446 2384 476
rect 2350 374 2384 408
rect 2350 306 2384 336
rect 2350 302 2384 306
rect 2350 238 2384 264
rect 2350 230 2384 238
rect 1297 174 1331 208
rect 2508 518 2542 544
rect 2666 544 2700 552
rect 2508 476 2542 480
rect 2508 446 2542 476
rect 2508 374 2542 408
rect 2508 306 2542 336
rect 2508 302 2542 306
rect 2508 238 2542 264
rect 2508 230 2542 238
rect 2666 518 2700 544
rect 2931 623 2965 643
rect 2931 609 2965 623
rect 2931 555 2965 571
rect 2931 537 2965 555
rect 2666 476 2700 480
rect 2666 446 2700 476
rect 2666 374 2700 408
rect 2931 487 2965 499
rect 2931 465 2965 487
rect 2931 419 2965 427
rect 2931 393 2965 419
rect 2931 351 2965 355
rect 2666 306 2700 336
rect 2666 302 2700 306
rect 2666 238 2700 264
rect 2666 230 2700 238
rect 2808 313 2842 347
rect 2931 321 2965 351
rect 3089 1405 3123 1435
rect 3089 1401 3123 1405
rect 3089 1337 3123 1363
rect 3089 1329 3123 1337
rect 3089 1269 3123 1291
rect 3089 1257 3123 1269
rect 3089 1201 3123 1219
rect 3089 1185 3123 1201
rect 3089 1133 3123 1147
rect 3089 1113 3123 1133
rect 3089 1065 3123 1075
rect 3089 1041 3123 1065
rect 3089 997 3123 1003
rect 3089 969 3123 997
rect 3089 929 3123 931
rect 3089 897 3123 929
rect 3089 827 3123 859
rect 3089 825 3123 827
rect 3089 759 3123 787
rect 3089 753 3123 759
rect 3089 691 3123 715
rect 3089 681 3123 691
rect 3089 623 3123 643
rect 3089 609 3123 623
rect 3089 555 3123 571
rect 3089 537 3123 555
rect 3089 487 3123 499
rect 3089 465 3123 487
rect 3089 419 3123 427
rect 3089 393 3123 419
rect 3089 351 3123 355
rect 3089 321 3123 351
rect 3247 1405 3281 1435
rect 3247 1401 3281 1405
rect 3247 1337 3281 1363
rect 3247 1329 3281 1337
rect 3247 1269 3281 1291
rect 3247 1257 3281 1269
rect 3247 1201 3281 1219
rect 3247 1185 3281 1201
rect 3247 1133 3281 1147
rect 3247 1113 3281 1133
rect 3247 1065 3281 1075
rect 3247 1041 3281 1065
rect 3247 997 3281 1003
rect 3247 969 3281 997
rect 3247 929 3281 931
rect 3247 897 3281 929
rect 3247 827 3281 859
rect 3247 825 3281 827
rect 3247 759 3281 787
rect 3247 753 3281 759
rect 3247 691 3281 715
rect 3247 681 3281 691
rect 3247 623 3281 643
rect 3247 609 3281 623
rect 3247 555 3281 571
rect 3247 537 3281 555
rect 3247 487 3281 499
rect 3247 465 3281 487
rect 3247 419 3281 427
rect 3247 393 3281 419
rect 3247 351 3281 355
rect 3247 321 3281 351
rect 3405 1405 3439 1435
rect 3405 1401 3439 1405
rect 3405 1337 3439 1363
rect 3405 1329 3439 1337
rect 3405 1269 3439 1291
rect 3405 1257 3439 1269
rect 3405 1201 3439 1219
rect 3405 1185 3439 1201
rect 3405 1133 3439 1147
rect 3405 1113 3439 1133
rect 3405 1065 3439 1075
rect 3405 1041 3439 1065
rect 3405 997 3439 1003
rect 3405 969 3439 997
rect 3405 929 3439 931
rect 3405 897 3439 929
rect 3405 827 3439 859
rect 3405 825 3439 827
rect 3405 759 3439 787
rect 3405 753 3439 759
rect 3405 691 3439 715
rect 3405 681 3439 691
rect 3405 623 3439 643
rect 3405 609 3439 623
rect 3405 555 3439 571
rect 3405 537 3439 555
rect 3405 487 3439 499
rect 3405 465 3439 487
rect 3405 419 3439 427
rect 3405 393 3439 419
rect 3405 351 3439 355
rect 3405 321 3439 351
rect 3563 1405 3597 1435
rect 3563 1401 3597 1405
rect 3563 1337 3597 1363
rect 3563 1329 3597 1337
rect 3563 1269 3597 1291
rect 3563 1257 3597 1269
rect 3563 1201 3597 1219
rect 3563 1185 3597 1201
rect 3563 1133 3597 1147
rect 3563 1113 3597 1133
rect 3563 1065 3597 1075
rect 3563 1041 3597 1065
rect 3563 997 3597 1003
rect 3563 969 3597 997
rect 3563 929 3597 931
rect 3563 897 3597 929
rect 3563 827 3597 859
rect 3563 825 3597 827
rect 3563 759 3597 787
rect 3563 753 3597 759
rect 3563 691 3597 715
rect 3563 681 3597 691
rect 3563 623 3597 643
rect 3563 609 3597 623
rect 3563 555 3597 571
rect 3563 537 3597 555
rect 3563 487 3597 499
rect 3563 465 3597 487
rect 3563 419 3597 427
rect 3563 393 3597 419
rect 3563 351 3597 355
rect 3563 321 3597 351
rect -595 76 -562 99
rect -562 76 -561 99
rect -595 65 -561 76
rect -271 55 -237 89
rect -49 51 -15 85
rect 72 61 106 95
rect 240 59 274 93
rect 409 59 443 93
rect 578 61 612 95
rect 757 65 791 99
rect 944 65 978 99
rect 1145 63 1179 97
<< metal1 >>
rect 1862 3932 2788 3933
rect -157 3931 2788 3932
rect -162 3923 2788 3931
rect 2913 3923 2973 3935
rect -162 3916 2973 3923
rect -162 3885 2926 3916
rect -162 3884 -76 3885
rect -174 3858 -76 3884
rect -174 3824 -142 3858
rect -108 3824 -76 3858
rect -174 3798 -76 3824
rect 773 3813 819 3836
rect 773 3779 779 3813
rect 813 3779 819 3813
rect 773 3741 819 3779
rect 773 3707 779 3741
rect 813 3707 819 3741
rect 773 3669 819 3707
rect 773 3635 779 3669
rect 813 3635 819 3669
rect 773 3597 819 3635
rect 773 3563 779 3597
rect 813 3563 819 3597
rect 773 3525 819 3563
rect 773 3491 779 3525
rect 813 3491 819 3525
rect 773 3453 819 3491
rect 773 3419 779 3453
rect 813 3419 819 3453
rect 773 3381 819 3419
rect 773 3347 779 3381
rect 813 3347 819 3381
rect 773 3309 819 3347
rect 773 3275 779 3309
rect 813 3275 819 3309
rect 773 3237 819 3275
rect 773 3203 779 3237
rect 813 3203 819 3237
rect 773 3165 819 3203
rect 773 3131 779 3165
rect 813 3131 819 3165
rect 773 3093 819 3131
rect 773 3059 779 3093
rect 813 3059 819 3093
rect 773 3036 819 3059
rect 931 3813 978 3885
rect 1166 3882 2926 3885
rect 2960 3882 2973 3916
rect 1166 3875 2973 3882
rect 1166 3836 2788 3875
rect 2913 3863 2973 3875
rect 3068 3872 3074 3924
rect 3126 3875 3445 3924
rect 3126 3872 3132 3875
rect 931 3779 937 3813
rect 971 3811 978 3813
rect 1089 3813 1135 3836
rect 971 3779 977 3811
rect 931 3741 977 3779
rect 931 3707 937 3741
rect 971 3707 977 3741
rect 931 3669 977 3707
rect 931 3635 937 3669
rect 971 3635 977 3669
rect 931 3597 977 3635
rect 931 3563 937 3597
rect 971 3563 977 3597
rect 931 3525 977 3563
rect 931 3491 937 3525
rect 971 3491 977 3525
rect 931 3453 977 3491
rect 931 3419 937 3453
rect 971 3419 977 3453
rect 931 3381 977 3419
rect 931 3347 937 3381
rect 971 3347 977 3381
rect 931 3309 977 3347
rect 931 3275 937 3309
rect 971 3275 977 3309
rect 931 3237 977 3275
rect 931 3203 937 3237
rect 971 3203 977 3237
rect 931 3165 977 3203
rect 931 3131 937 3165
rect 971 3131 977 3165
rect 931 3093 977 3131
rect 931 3059 937 3093
rect 971 3059 977 3093
rect 931 3036 977 3059
rect 1089 3779 1095 3813
rect 1129 3779 1135 3813
rect 1089 3741 1135 3779
rect 1089 3707 1095 3741
rect 1129 3707 1135 3741
rect 1166 3802 1353 3836
rect 1387 3833 2788 3836
rect 1387 3831 2537 3833
rect 1387 3802 1577 3831
rect 1166 3797 1577 3802
rect 1611 3830 2537 3831
rect 1611 3828 2043 3830
rect 1611 3797 1820 3828
rect 1166 3794 1820 3797
rect 1854 3796 2043 3828
rect 2077 3796 2115 3830
rect 2149 3828 2537 3830
rect 2149 3796 2278 3828
rect 1854 3794 2278 3796
rect 2312 3794 2350 3828
rect 2384 3799 2537 3828
rect 2571 3799 2609 3833
rect 2643 3799 2788 3833
rect 2384 3794 2788 3799
rect 1166 3718 2788 3794
rect 1089 3669 1135 3707
rect 1089 3635 1095 3669
rect 1129 3635 1135 3669
rect 1089 3597 1135 3635
rect 1089 3563 1095 3597
rect 1129 3563 1135 3597
rect 1089 3525 1135 3563
rect 1089 3491 1095 3525
rect 1129 3491 1135 3525
rect 1390 3522 1443 3718
rect 1862 3717 2788 3718
rect 2920 3764 2966 3811
rect 3075 3796 3124 3872
rect 2920 3730 2926 3764
rect 2960 3730 2966 3764
rect 1089 3453 1135 3491
rect 1089 3419 1095 3453
rect 1129 3419 1135 3453
rect 1089 3381 1135 3419
rect 1089 3347 1095 3381
rect 1129 3347 1135 3381
rect 1089 3309 1135 3347
rect 1089 3275 1095 3309
rect 1129 3275 1135 3309
rect 1089 3237 1135 3275
rect 1089 3203 1095 3237
rect 1129 3203 1135 3237
rect 1089 3165 1135 3203
rect 1089 3131 1095 3165
rect 1129 3131 1135 3165
rect 1397 3501 1443 3522
rect 1397 3467 1403 3501
rect 1437 3467 1443 3501
rect 1397 3429 1443 3467
rect 1397 3395 1403 3429
rect 1437 3395 1443 3429
rect 1397 3357 1443 3395
rect 1397 3323 1403 3357
rect 1437 3323 1443 3357
rect 1397 3285 1443 3323
rect 1397 3251 1403 3285
rect 1437 3251 1443 3285
rect 1397 3213 1443 3251
rect 1397 3179 1403 3213
rect 1437 3179 1443 3213
rect 1397 3140 1443 3179
rect 1555 3501 1601 3540
rect 1555 3467 1561 3501
rect 1595 3467 1601 3501
rect 1555 3429 1601 3467
rect 1555 3395 1561 3429
rect 1595 3395 1601 3429
rect 1555 3357 1601 3395
rect 1555 3323 1561 3357
rect 1595 3323 1601 3357
rect 1555 3285 1601 3323
rect 1555 3251 1561 3285
rect 1595 3251 1601 3285
rect 1555 3213 1601 3251
rect 1555 3179 1561 3213
rect 1595 3179 1601 3213
rect 1555 3165 1601 3179
rect 1555 3140 1605 3165
rect 1089 3093 1135 3131
rect 1089 3059 1095 3093
rect 1129 3059 1135 3093
rect 1225 3118 1289 3127
rect 1225 3084 1240 3118
rect 1274 3084 1289 3118
rect 1225 3075 1289 3084
rect 1089 3036 1135 3059
rect 995 2937 1044 2948
rect 1237 2937 1277 3075
rect 1557 3007 1605 3140
rect 995 2934 1277 2937
rect 995 2900 1002 2934
rect 1036 2900 1277 2934
rect 1398 2984 1444 3007
rect 1398 2950 1404 2984
rect 1438 2950 1444 2984
rect 1398 2912 1444 2950
rect 995 2887 1044 2900
rect 1398 2878 1404 2912
rect 1438 2878 1444 2912
rect 1398 2840 1444 2878
rect 1398 2806 1404 2840
rect 1438 2806 1444 2840
rect 1398 2768 1444 2806
rect 1398 2734 1404 2768
rect 1438 2734 1444 2768
rect 873 2663 919 2702
rect 873 2629 879 2663
rect 913 2629 919 2663
rect 873 2591 919 2629
rect 873 2557 879 2591
rect 913 2557 919 2591
rect 873 2519 919 2557
rect 873 2485 879 2519
rect 913 2485 919 2519
rect 873 2447 919 2485
rect 873 2413 879 2447
rect 913 2413 919 2447
rect 873 2396 919 2413
rect 1031 2663 1077 2702
rect 1031 2629 1037 2663
rect 1071 2629 1077 2663
rect 1031 2591 1077 2629
rect 1031 2557 1037 2591
rect 1071 2557 1077 2591
rect 1031 2519 1077 2557
rect 1031 2485 1037 2519
rect 1071 2485 1077 2519
rect 1031 2447 1077 2485
rect 1031 2413 1037 2447
rect 1071 2413 1077 2447
rect 861 2375 922 2396
rect 861 2341 879 2375
rect 913 2341 922 2375
rect 861 2171 922 2341
rect 1031 2375 1077 2413
rect 1031 2341 1037 2375
rect 1071 2341 1077 2375
rect 1031 2302 1077 2341
rect 1398 2696 1444 2734
rect 1398 2662 1404 2696
rect 1438 2662 1444 2696
rect 1398 2624 1444 2662
rect 1398 2590 1404 2624
rect 1438 2590 1444 2624
rect 1398 2552 1444 2590
rect 1398 2518 1404 2552
rect 1438 2518 1444 2552
rect 1398 2480 1444 2518
rect 1398 2446 1404 2480
rect 1438 2446 1444 2480
rect 1398 2408 1444 2446
rect 1398 2374 1404 2408
rect 1438 2374 1444 2408
rect 1398 2336 1444 2374
rect 1398 2302 1404 2336
rect 1438 2302 1444 2336
rect 1398 2264 1444 2302
rect 1398 2257 1404 2264
rect 745 2117 922 2171
rect 1383 2230 1404 2257
rect 1438 2230 1444 2264
rect 1383 2207 1444 2230
rect 1556 2989 1605 3007
rect 1556 2984 1602 2989
rect 1556 2950 1562 2984
rect 1596 2950 1602 2984
rect 1556 2912 1602 2950
rect 1556 2878 1562 2912
rect 1596 2878 1602 2912
rect 1556 2840 1602 2878
rect 1556 2806 1562 2840
rect 1596 2806 1602 2840
rect 1556 2768 1602 2806
rect 1556 2734 1562 2768
rect 1596 2734 1602 2768
rect 1556 2696 1602 2734
rect 1556 2662 1562 2696
rect 1596 2662 1602 2696
rect 1556 2624 1602 2662
rect 1556 2590 1562 2624
rect 1596 2590 1602 2624
rect 1556 2552 1602 2590
rect 1556 2518 1562 2552
rect 1596 2518 1602 2552
rect 1556 2480 1602 2518
rect 1556 2446 1562 2480
rect 1596 2446 1602 2480
rect 1556 2408 1602 2446
rect 1556 2374 1562 2408
rect 1596 2374 1602 2408
rect 1556 2336 1602 2374
rect 1556 2302 1562 2336
rect 1596 2302 1602 2336
rect 1556 2264 1602 2302
rect 1556 2230 1562 2264
rect 1596 2230 1602 2264
rect 1556 2207 1602 2230
rect 1714 2984 1760 3007
rect 1714 2950 1720 2984
rect 1754 2950 1760 2984
rect 1714 2912 1760 2950
rect 1714 2878 1720 2912
rect 1754 2878 1760 2912
rect 1714 2840 1760 2878
rect 1714 2806 1720 2840
rect 1754 2806 1760 2840
rect 1714 2768 1760 2806
rect 1714 2734 1720 2768
rect 1754 2734 1760 2768
rect 1714 2696 1760 2734
rect 1714 2662 1720 2696
rect 1754 2662 1760 2696
rect 1714 2624 1760 2662
rect 1714 2590 1720 2624
rect 1754 2590 1760 2624
rect 1714 2552 1760 2590
rect 1714 2518 1720 2552
rect 1754 2518 1760 2552
rect 1714 2480 1760 2518
rect 1714 2446 1720 2480
rect 1754 2446 1760 2480
rect 1714 2408 1760 2446
rect 1714 2374 1720 2408
rect 1754 2374 1760 2408
rect 1866 2399 1910 3717
rect 2174 3565 2220 3588
rect 2174 3531 2180 3565
rect 2214 3531 2220 3565
rect 2331 3565 2378 3717
rect 2920 3692 2966 3730
rect 2826 3620 2832 3672
rect 2884 3620 2890 3672
rect 2920 3658 2926 3692
rect 2960 3658 2966 3692
rect 2920 3620 2966 3658
rect 2331 3541 2338 3565
rect 2174 3493 2220 3531
rect 2174 3459 2180 3493
rect 2214 3459 2220 3493
rect 2174 3421 2220 3459
rect 2174 3387 2180 3421
rect 2214 3387 2220 3421
rect 2174 3349 2220 3387
rect 2174 3315 2180 3349
rect 2214 3315 2220 3349
rect 2174 3277 2220 3315
rect 2174 3243 2180 3277
rect 2214 3243 2220 3277
rect 2174 3205 2220 3243
rect 2174 3171 2180 3205
rect 2214 3171 2220 3205
rect 2174 3133 2220 3171
rect 2174 3099 2180 3133
rect 2214 3099 2220 3133
rect 2174 3061 2220 3099
rect 2174 3027 2180 3061
rect 2214 3027 2220 3061
rect 2174 2989 2220 3027
rect 2174 2955 2180 2989
rect 2214 2955 2220 2989
rect 2174 2917 2220 2955
rect 2174 2883 2180 2917
rect 2214 2883 2220 2917
rect 2174 2845 2220 2883
rect 2174 2811 2180 2845
rect 2214 2811 2220 2845
rect 2174 2788 2220 2811
rect 2332 3531 2338 3541
rect 2372 3531 2378 3565
rect 2332 3493 2378 3531
rect 2332 3459 2338 3493
rect 2372 3459 2378 3493
rect 2332 3421 2378 3459
rect 2332 3387 2338 3421
rect 2372 3387 2378 3421
rect 2332 3349 2378 3387
rect 2332 3315 2338 3349
rect 2372 3315 2378 3349
rect 2332 3277 2378 3315
rect 2332 3243 2338 3277
rect 2372 3243 2378 3277
rect 2332 3205 2378 3243
rect 2332 3171 2338 3205
rect 2372 3171 2378 3205
rect 2332 3133 2378 3171
rect 2332 3099 2338 3133
rect 2372 3099 2378 3133
rect 2332 3061 2378 3099
rect 2332 3027 2338 3061
rect 2372 3027 2378 3061
rect 2332 2989 2378 3027
rect 2332 2955 2338 2989
rect 2372 2955 2378 2989
rect 2332 2917 2378 2955
rect 2332 2883 2338 2917
rect 2372 2883 2378 2917
rect 2332 2845 2378 2883
rect 2332 2811 2338 2845
rect 2372 2811 2378 2845
rect 2332 2788 2378 2811
rect 2490 3565 2536 3588
rect 2490 3531 2496 3565
rect 2530 3531 2536 3565
rect 2490 3493 2536 3531
rect 2490 3459 2496 3493
rect 2530 3459 2536 3493
rect 2490 3421 2536 3459
rect 2490 3387 2496 3421
rect 2530 3387 2536 3421
rect 2490 3349 2536 3387
rect 2490 3315 2496 3349
rect 2530 3315 2536 3349
rect 2490 3277 2536 3315
rect 2490 3243 2496 3277
rect 2530 3243 2536 3277
rect 2490 3205 2536 3243
rect 2490 3171 2496 3205
rect 2530 3171 2536 3205
rect 2490 3133 2536 3171
rect 2490 3099 2496 3133
rect 2530 3099 2536 3133
rect 2490 3061 2536 3099
rect 2490 3027 2496 3061
rect 2530 3027 2536 3061
rect 2490 2989 2536 3027
rect 2490 2955 2496 2989
rect 2530 2955 2536 2989
rect 2490 2917 2536 2955
rect 2490 2883 2496 2917
rect 2530 2883 2536 2917
rect 2490 2845 2536 2883
rect 2490 2811 2496 2845
rect 2530 2831 2536 2845
rect 2530 2811 2550 2831
rect 2490 2788 2550 2811
rect 2174 2676 2219 2788
rect 2174 2631 2322 2676
rect 2277 2490 2322 2631
rect 2505 2652 2550 2788
rect 2607 2652 2664 2663
rect 2505 2645 2664 2652
rect 2505 2627 2618 2645
rect 2117 2451 2163 2490
rect 2117 2417 2123 2451
rect 2157 2417 2163 2451
rect 1714 2336 1760 2374
rect 1856 2347 1862 2399
rect 1914 2347 1920 2399
rect 2117 2379 2163 2417
rect 1714 2302 1720 2336
rect 1754 2302 1760 2336
rect 1714 2264 1760 2302
rect 1714 2230 1720 2264
rect 1754 2230 1760 2264
rect 1714 2207 1760 2230
rect 2117 2345 2123 2379
rect 2157 2345 2163 2379
rect 2117 2307 2163 2345
rect 2117 2273 2123 2307
rect 2157 2273 2163 2307
rect 2117 2235 2163 2273
rect 745 2110 921 2117
rect 745 1628 806 2110
rect 1383 2084 1426 2207
rect 2117 2201 2123 2235
rect 2157 2201 2163 2235
rect 2117 2163 2163 2201
rect 2117 2129 2123 2163
rect 2157 2129 2163 2163
rect 2117 2090 2163 2129
rect 2275 2458 2322 2490
rect 2392 2611 2618 2627
rect 2652 2611 2664 2645
rect 2392 2607 2664 2611
rect 2392 2582 2550 2607
rect 2607 2594 2664 2607
rect 2392 2494 2437 2582
rect 2392 2459 2440 2494
rect 2275 2451 2321 2458
rect 2275 2417 2281 2451
rect 2315 2417 2321 2451
rect 2275 2379 2321 2417
rect 2275 2345 2281 2379
rect 2315 2345 2321 2379
rect 2275 2307 2321 2345
rect 2275 2273 2281 2307
rect 2315 2273 2321 2307
rect 2275 2235 2321 2273
rect 2275 2201 2281 2235
rect 2315 2201 2321 2235
rect 2275 2163 2321 2201
rect 2275 2129 2281 2163
rect 2315 2129 2321 2163
rect 2275 2090 2321 2129
rect 2394 2455 2440 2459
rect 2394 2421 2400 2455
rect 2434 2421 2440 2455
rect 2394 2383 2440 2421
rect 2394 2349 2400 2383
rect 2434 2349 2440 2383
rect 2394 2311 2440 2349
rect 2394 2277 2400 2311
rect 2434 2277 2440 2311
rect 2394 2239 2440 2277
rect 2394 2205 2400 2239
rect 2434 2205 2440 2239
rect 2394 2167 2440 2205
rect 2394 2133 2400 2167
rect 2434 2133 2440 2167
rect 2394 2094 2440 2133
rect 2552 2455 2598 2494
rect 2552 2421 2558 2455
rect 2592 2421 2598 2455
rect 2552 2383 2598 2421
rect 2552 2349 2558 2383
rect 2592 2349 2598 2383
rect 2552 2311 2598 2349
rect 2724 2362 2795 2375
rect 2724 2328 2742 2362
rect 2776 2328 2795 2362
rect 2724 2316 2795 2328
rect 2552 2277 2558 2311
rect 2592 2277 2598 2311
rect 2552 2239 2598 2277
rect 2552 2205 2558 2239
rect 2592 2205 2598 2239
rect 2552 2167 2598 2205
rect 2552 2133 2558 2167
rect 2592 2133 2598 2167
rect 2552 2129 2598 2133
rect 2552 2094 2600 2129
rect 1383 2041 1990 2084
rect 1784 1983 1836 1989
rect 1403 1956 1465 1964
rect 1403 1922 1417 1956
rect 1451 1922 1465 1956
rect 1403 1914 1465 1922
rect 1740 1931 1784 1936
rect 1947 1987 1990 2041
rect 2118 1987 2161 2090
rect 2557 2005 2600 2094
rect 1947 1982 2161 1987
rect 2509 1999 2600 2005
rect 1947 1944 2235 1982
rect 2509 1965 2521 1999
rect 2555 1965 2600 1999
rect 2509 1960 2600 1965
rect 2509 1959 2567 1960
rect 2118 1939 2235 1944
rect 1740 1925 1836 1931
rect 412 1567 806 1628
rect 943 1682 989 1721
rect 943 1648 949 1682
rect 983 1648 989 1682
rect 943 1610 989 1648
rect 943 1576 949 1610
rect 983 1576 989 1610
rect 104 1355 177 1366
rect 412 1355 473 1567
rect 943 1538 989 1576
rect 943 1504 949 1538
rect 983 1504 989 1538
rect 943 1466 989 1504
rect 835 1454 887 1460
rect 670 1409 835 1448
rect 104 1340 479 1355
rect 104 1306 123 1340
rect 157 1339 479 1340
rect 157 1306 481 1339
rect 104 1294 481 1306
rect 104 1281 177 1294
rect 77 990 222 1013
rect 77 956 165 990
rect 199 956 222 990
rect 77 934 222 956
rect -692 157 66 158
rect 435 157 481 1294
rect 518 992 576 996
rect 670 992 709 1409
rect 835 1396 887 1402
rect 943 1432 949 1466
rect 983 1432 989 1466
rect 943 1394 989 1432
rect 943 1376 949 1394
rect 937 1360 949 1376
rect 983 1360 989 1394
rect 937 1321 989 1360
rect 1101 1682 1147 1721
rect 1101 1648 1107 1682
rect 1141 1648 1147 1682
rect 1101 1610 1147 1648
rect 1101 1576 1107 1610
rect 1141 1576 1147 1610
rect 1101 1538 1147 1576
rect 1101 1504 1107 1538
rect 1141 1504 1147 1538
rect 1101 1466 1147 1504
rect 1101 1432 1107 1466
rect 1141 1432 1147 1466
rect 1101 1394 1147 1432
rect 1101 1360 1107 1394
rect 1141 1360 1147 1394
rect 1101 1356 1147 1360
rect 1259 1682 1305 1721
rect 1259 1648 1265 1682
rect 1299 1648 1305 1682
rect 1259 1610 1305 1648
rect 1409 1624 1459 1914
rect 1740 1892 1832 1925
rect 1740 1741 1784 1892
rect 1578 1718 1624 1741
rect 1578 1684 1584 1718
rect 1618 1684 1624 1718
rect 1578 1646 1624 1684
rect 1259 1576 1265 1610
rect 1299 1576 1305 1610
rect 1259 1538 1305 1576
rect 1402 1572 1408 1624
rect 1460 1572 1466 1624
rect 1578 1612 1584 1646
rect 1618 1612 1624 1646
rect 1578 1574 1624 1612
rect 1259 1504 1265 1538
rect 1299 1504 1305 1538
rect 1259 1466 1305 1504
rect 1259 1432 1265 1466
rect 1299 1432 1305 1466
rect 1578 1540 1584 1574
rect 1618 1540 1624 1574
rect 1578 1502 1624 1540
rect 1578 1468 1584 1502
rect 1618 1468 1624 1502
rect 1360 1453 1411 1458
rect 1259 1394 1305 1432
rect 1354 1401 1360 1453
rect 1412 1401 1418 1453
rect 1578 1430 1624 1468
rect 1360 1395 1411 1401
rect 1578 1396 1584 1430
rect 1618 1396 1624 1430
rect 1259 1360 1265 1394
rect 1299 1360 1305 1394
rect 1101 1321 1154 1356
rect 937 1282 986 1321
rect 842 1233 986 1282
rect 842 1193 891 1233
rect 834 1141 840 1193
rect 892 1141 898 1193
rect 1106 1176 1154 1321
rect 1259 1277 1305 1360
rect 1578 1358 1624 1396
rect 1578 1324 1584 1358
rect 1618 1324 1624 1358
rect 1578 1286 1624 1324
rect 1259 1231 1364 1277
rect 1578 1252 1584 1286
rect 1618 1252 1624 1286
rect 1312 1200 1361 1231
rect 1578 1214 1624 1252
rect 947 1153 993 1176
rect 518 990 709 992
rect 518 956 530 990
rect 564 956 709 990
rect 518 953 709 956
rect 947 1119 953 1153
rect 987 1119 993 1153
rect 947 1081 993 1119
rect 947 1047 953 1081
rect 987 1047 993 1081
rect 947 1009 993 1047
rect 947 975 953 1009
rect 987 975 993 1009
rect 518 950 576 953
rect 947 937 993 975
rect 947 903 953 937
rect 987 903 993 937
rect 947 865 993 903
rect 947 831 953 865
rect 987 831 993 865
rect 947 793 993 831
rect 947 759 953 793
rect 987 759 993 793
rect 618 719 670 725
rect 947 721 993 759
rect 612 667 618 719
rect 670 667 676 719
rect 947 687 953 721
rect 987 687 993 721
rect 618 663 670 667
rect 947 649 993 687
rect 947 615 953 649
rect 987 615 993 649
rect 947 577 993 615
rect 947 543 953 577
rect 987 543 993 577
rect 947 505 993 543
rect 947 471 953 505
rect 987 471 993 505
rect 947 433 993 471
rect 947 399 953 433
rect 987 399 993 433
rect 676 349 728 355
rect 670 297 676 349
rect 676 291 728 297
rect 947 157 993 399
rect 1105 1158 1154 1176
rect 1300 1186 1373 1200
rect 1105 1153 1151 1158
rect 1105 1119 1111 1153
rect 1145 1119 1151 1153
rect 1300 1152 1319 1186
rect 1353 1152 1373 1186
rect 1300 1139 1373 1152
rect 1578 1180 1584 1214
rect 1618 1180 1624 1214
rect 1578 1142 1624 1180
rect 1105 1081 1151 1119
rect 1105 1047 1111 1081
rect 1145 1047 1151 1081
rect 1105 1009 1151 1047
rect 1105 975 1111 1009
rect 1145 975 1151 1009
rect 1578 1108 1584 1142
rect 1618 1108 1624 1142
rect 1578 1070 1624 1108
rect 1578 1036 1584 1070
rect 1618 1036 1624 1070
rect 1578 998 1624 1036
rect 1578 986 1584 998
rect 1105 937 1151 975
rect 1105 903 1111 937
rect 1145 903 1151 937
rect 1576 964 1584 986
rect 1618 986 1624 998
rect 1736 1718 1784 1741
rect 1736 1684 1742 1718
rect 1776 1712 1784 1718
rect 1894 1718 1940 1741
rect 1776 1684 1782 1712
rect 1736 1646 1782 1684
rect 1736 1612 1742 1646
rect 1776 1612 1782 1646
rect 1736 1574 1782 1612
rect 1736 1540 1742 1574
rect 1776 1540 1782 1574
rect 1736 1502 1782 1540
rect 1736 1468 1742 1502
rect 1776 1468 1782 1502
rect 1736 1430 1782 1468
rect 1736 1396 1742 1430
rect 1776 1396 1782 1430
rect 1736 1358 1782 1396
rect 1736 1324 1742 1358
rect 1776 1324 1782 1358
rect 1736 1286 1782 1324
rect 1736 1252 1742 1286
rect 1776 1252 1782 1286
rect 1736 1214 1782 1252
rect 1736 1180 1742 1214
rect 1776 1180 1782 1214
rect 1736 1142 1782 1180
rect 1736 1108 1742 1142
rect 1776 1108 1782 1142
rect 1736 1070 1782 1108
rect 1736 1036 1742 1070
rect 1776 1036 1782 1070
rect 1736 998 1782 1036
rect 1618 964 1625 986
rect 1105 865 1151 903
rect 1105 831 1111 865
rect 1145 831 1151 865
rect 1285 917 1337 923
rect 1576 915 1625 964
rect 1736 964 1742 998
rect 1776 964 1782 998
rect 1894 1684 1900 1718
rect 1934 1684 1940 1718
rect 2192 1689 2235 1939
rect 2512 1689 2555 1959
rect 2736 1773 2783 2316
rect 2834 1911 2883 3620
rect 2834 1877 2841 1911
rect 2875 1877 2883 1911
rect 2834 1864 2883 1877
rect 2920 3586 2926 3620
rect 2960 3586 2966 3620
rect 2920 3548 2966 3586
rect 2920 3514 2926 3548
rect 2960 3514 2966 3548
rect 2920 3476 2966 3514
rect 2920 3442 2926 3476
rect 2960 3442 2966 3476
rect 2920 3404 2966 3442
rect 2920 3370 2926 3404
rect 2960 3370 2966 3404
rect 2920 3332 2966 3370
rect 2920 3298 2926 3332
rect 2960 3298 2966 3332
rect 2920 3260 2966 3298
rect 2920 3226 2926 3260
rect 2960 3226 2966 3260
rect 2920 3188 2966 3226
rect 2920 3154 2926 3188
rect 2960 3154 2966 3188
rect 2920 3116 2966 3154
rect 2920 3082 2926 3116
rect 2960 3082 2966 3116
rect 2920 3044 2966 3082
rect 2920 3010 2926 3044
rect 2960 3010 2966 3044
rect 2920 2972 2966 3010
rect 2920 2938 2926 2972
rect 2960 2938 2966 2972
rect 2920 2900 2966 2938
rect 2920 2866 2926 2900
rect 2960 2866 2966 2900
rect 2920 2828 2966 2866
rect 2920 2794 2926 2828
rect 2960 2794 2966 2828
rect 2920 2756 2966 2794
rect 2920 2722 2926 2756
rect 2960 2722 2966 2756
rect 2920 2684 2966 2722
rect 2920 2650 2926 2684
rect 2960 2650 2966 2684
rect 2920 2612 2966 2650
rect 2920 2578 2926 2612
rect 2960 2578 2966 2612
rect 2920 2540 2966 2578
rect 2920 2506 2926 2540
rect 2960 2506 2966 2540
rect 2920 2468 2966 2506
rect 2920 2434 2926 2468
rect 2960 2434 2966 2468
rect 2920 2396 2966 2434
rect 2920 2362 2926 2396
rect 2960 2362 2966 2396
rect 2920 2324 2966 2362
rect 2920 2290 2926 2324
rect 2960 2290 2966 2324
rect 2920 2252 2966 2290
rect 2920 2218 2926 2252
rect 2960 2218 2966 2252
rect 2920 2180 2966 2218
rect 2920 2146 2926 2180
rect 2960 2146 2966 2180
rect 2920 2108 2966 2146
rect 2920 2074 2926 2108
rect 2960 2074 2966 2108
rect 2920 2036 2966 2074
rect 2920 2002 2926 2036
rect 2960 2002 2966 2036
rect 2920 1964 2966 2002
rect 2920 1930 2926 1964
rect 2960 1930 2966 1964
rect 2920 1892 2966 1930
rect 2920 1858 2926 1892
rect 2960 1858 2966 1892
rect 2920 1811 2966 1858
rect 3078 3764 3124 3796
rect 3078 3730 3084 3764
rect 3118 3730 3124 3764
rect 3078 3692 3124 3730
rect 3078 3658 3084 3692
rect 3118 3658 3124 3692
rect 3078 3620 3124 3658
rect 3078 3586 3084 3620
rect 3118 3586 3124 3620
rect 3078 3548 3124 3586
rect 3078 3514 3084 3548
rect 3118 3514 3124 3548
rect 3078 3476 3124 3514
rect 3078 3442 3084 3476
rect 3118 3442 3124 3476
rect 3078 3404 3124 3442
rect 3078 3370 3084 3404
rect 3118 3370 3124 3404
rect 3078 3332 3124 3370
rect 3078 3298 3084 3332
rect 3118 3298 3124 3332
rect 3078 3260 3124 3298
rect 3078 3226 3084 3260
rect 3118 3226 3124 3260
rect 3078 3188 3124 3226
rect 3078 3154 3084 3188
rect 3118 3154 3124 3188
rect 3078 3116 3124 3154
rect 3078 3082 3084 3116
rect 3118 3082 3124 3116
rect 3078 3044 3124 3082
rect 3078 3010 3084 3044
rect 3118 3010 3124 3044
rect 3078 2972 3124 3010
rect 3078 2938 3084 2972
rect 3118 2938 3124 2972
rect 3078 2900 3124 2938
rect 3078 2866 3084 2900
rect 3118 2866 3124 2900
rect 3078 2828 3124 2866
rect 3078 2794 3084 2828
rect 3118 2794 3124 2828
rect 3078 2756 3124 2794
rect 3078 2722 3084 2756
rect 3118 2722 3124 2756
rect 3078 2684 3124 2722
rect 3078 2650 3084 2684
rect 3118 2650 3124 2684
rect 3078 2612 3124 2650
rect 3078 2578 3084 2612
rect 3118 2578 3124 2612
rect 3078 2540 3124 2578
rect 3078 2506 3084 2540
rect 3118 2506 3124 2540
rect 3078 2468 3124 2506
rect 3078 2434 3084 2468
rect 3118 2434 3124 2468
rect 3078 2396 3124 2434
rect 3078 2362 3084 2396
rect 3118 2362 3124 2396
rect 3078 2324 3124 2362
rect 3078 2290 3084 2324
rect 3118 2290 3124 2324
rect 3078 2252 3124 2290
rect 3078 2218 3084 2252
rect 3118 2218 3124 2252
rect 3078 2180 3124 2218
rect 3078 2146 3084 2180
rect 3118 2146 3124 2180
rect 3078 2108 3124 2146
rect 3078 2074 3084 2108
rect 3118 2074 3124 2108
rect 3078 2036 3124 2074
rect 3078 2002 3084 2036
rect 3118 2002 3124 2036
rect 3078 1964 3124 2002
rect 3078 1930 3084 1964
rect 3118 1930 3124 1964
rect 3078 1892 3124 1930
rect 3078 1858 3084 1892
rect 3118 1858 3124 1892
rect 3078 1811 3124 1858
rect 3236 3764 3282 3811
rect 3392 3800 3441 3875
rect 3236 3730 3242 3764
rect 3276 3730 3282 3764
rect 3236 3692 3282 3730
rect 3236 3658 3242 3692
rect 3276 3658 3282 3692
rect 3236 3620 3282 3658
rect 3236 3586 3242 3620
rect 3276 3586 3282 3620
rect 3236 3548 3282 3586
rect 3236 3514 3242 3548
rect 3276 3514 3282 3548
rect 3236 3476 3282 3514
rect 3236 3442 3242 3476
rect 3276 3442 3282 3476
rect 3236 3404 3282 3442
rect 3236 3370 3242 3404
rect 3276 3370 3282 3404
rect 3236 3332 3282 3370
rect 3236 3298 3242 3332
rect 3276 3298 3282 3332
rect 3236 3260 3282 3298
rect 3236 3226 3242 3260
rect 3276 3226 3282 3260
rect 3236 3188 3282 3226
rect 3236 3154 3242 3188
rect 3276 3154 3282 3188
rect 3236 3116 3282 3154
rect 3236 3082 3242 3116
rect 3276 3082 3282 3116
rect 3236 3044 3282 3082
rect 3236 3010 3242 3044
rect 3276 3010 3282 3044
rect 3236 2972 3282 3010
rect 3236 2938 3242 2972
rect 3276 2938 3282 2972
rect 3236 2900 3282 2938
rect 3236 2866 3242 2900
rect 3276 2866 3282 2900
rect 3236 2828 3282 2866
rect 3236 2794 3242 2828
rect 3276 2794 3282 2828
rect 3236 2756 3282 2794
rect 3236 2722 3242 2756
rect 3276 2722 3282 2756
rect 3236 2684 3282 2722
rect 3236 2650 3242 2684
rect 3276 2650 3282 2684
rect 3236 2612 3282 2650
rect 3236 2578 3242 2612
rect 3276 2578 3282 2612
rect 3236 2540 3282 2578
rect 3236 2506 3242 2540
rect 3276 2506 3282 2540
rect 3236 2468 3282 2506
rect 3236 2434 3242 2468
rect 3276 2434 3282 2468
rect 3236 2396 3282 2434
rect 3236 2362 3242 2396
rect 3276 2362 3282 2396
rect 3236 2324 3282 2362
rect 3236 2290 3242 2324
rect 3276 2290 3282 2324
rect 3236 2252 3282 2290
rect 3236 2218 3242 2252
rect 3276 2218 3282 2252
rect 3236 2180 3282 2218
rect 3236 2146 3242 2180
rect 3276 2146 3282 2180
rect 3236 2108 3282 2146
rect 3236 2074 3242 2108
rect 3276 2074 3282 2108
rect 3236 2036 3282 2074
rect 3236 2002 3242 2036
rect 3276 2002 3282 2036
rect 3236 1964 3282 2002
rect 3236 1930 3242 1964
rect 3276 1930 3282 1964
rect 3236 1892 3282 1930
rect 3236 1858 3242 1892
rect 3276 1858 3282 1892
rect 3236 1811 3282 1858
rect 3394 3764 3440 3800
rect 3394 3730 3400 3764
rect 3434 3730 3440 3764
rect 3394 3692 3440 3730
rect 3394 3658 3400 3692
rect 3434 3658 3440 3692
rect 3394 3620 3440 3658
rect 3394 3586 3400 3620
rect 3434 3586 3440 3620
rect 3394 3548 3440 3586
rect 3394 3514 3400 3548
rect 3434 3514 3440 3548
rect 3394 3476 3440 3514
rect 3394 3442 3400 3476
rect 3434 3442 3440 3476
rect 3394 3404 3440 3442
rect 3394 3370 3400 3404
rect 3434 3370 3440 3404
rect 3394 3332 3440 3370
rect 3394 3298 3400 3332
rect 3434 3298 3440 3332
rect 3394 3260 3440 3298
rect 3394 3226 3400 3260
rect 3434 3226 3440 3260
rect 3394 3188 3440 3226
rect 3394 3154 3400 3188
rect 3434 3154 3440 3188
rect 3394 3116 3440 3154
rect 3394 3082 3400 3116
rect 3434 3082 3440 3116
rect 3394 3044 3440 3082
rect 3394 3010 3400 3044
rect 3434 3010 3440 3044
rect 3394 2972 3440 3010
rect 3394 2938 3400 2972
rect 3434 2938 3440 2972
rect 3394 2900 3440 2938
rect 3394 2866 3400 2900
rect 3434 2866 3440 2900
rect 3394 2828 3440 2866
rect 3394 2794 3400 2828
rect 3434 2794 3440 2828
rect 3394 2756 3440 2794
rect 3394 2722 3400 2756
rect 3434 2722 3440 2756
rect 3394 2684 3440 2722
rect 3394 2650 3400 2684
rect 3434 2650 3440 2684
rect 3394 2612 3440 2650
rect 3394 2578 3400 2612
rect 3434 2578 3440 2612
rect 3394 2540 3440 2578
rect 3394 2506 3400 2540
rect 3434 2506 3440 2540
rect 3394 2468 3440 2506
rect 3394 2434 3400 2468
rect 3434 2434 3440 2468
rect 3394 2396 3440 2434
rect 3394 2362 3400 2396
rect 3434 2362 3440 2396
rect 3394 2324 3440 2362
rect 3394 2290 3400 2324
rect 3434 2290 3440 2324
rect 3394 2252 3440 2290
rect 3394 2218 3400 2252
rect 3434 2218 3440 2252
rect 3394 2180 3440 2218
rect 3394 2146 3400 2180
rect 3434 2146 3440 2180
rect 3394 2108 3440 2146
rect 3394 2074 3400 2108
rect 3434 2074 3440 2108
rect 3394 2036 3440 2074
rect 3394 2002 3400 2036
rect 3434 2002 3440 2036
rect 3394 1964 3440 2002
rect 3394 1930 3400 1964
rect 3434 1930 3440 1964
rect 3394 1892 3440 1930
rect 3394 1858 3400 1892
rect 3434 1858 3440 1892
rect 3394 1811 3440 1858
rect 3552 3764 3598 3811
rect 3552 3730 3558 3764
rect 3592 3730 3598 3764
rect 3552 3692 3598 3730
rect 3552 3658 3558 3692
rect 3592 3658 3598 3692
rect 3552 3620 3598 3658
rect 3552 3586 3558 3620
rect 3592 3586 3598 3620
rect 3552 3548 3598 3586
rect 3552 3514 3558 3548
rect 3592 3514 3598 3548
rect 3552 3476 3598 3514
rect 3552 3442 3558 3476
rect 3592 3442 3598 3476
rect 3552 3404 3598 3442
rect 3552 3370 3558 3404
rect 3592 3370 3598 3404
rect 3552 3332 3598 3370
rect 3552 3298 3558 3332
rect 3592 3298 3598 3332
rect 3552 3260 3598 3298
rect 3552 3226 3558 3260
rect 3592 3226 3598 3260
rect 3552 3188 3598 3226
rect 3552 3154 3558 3188
rect 3592 3154 3598 3188
rect 3552 3116 3598 3154
rect 3552 3082 3558 3116
rect 3592 3082 3598 3116
rect 3552 3044 3598 3082
rect 3552 3010 3558 3044
rect 3592 3010 3598 3044
rect 3552 2972 3598 3010
rect 3552 2938 3558 2972
rect 3592 2938 3598 2972
rect 3552 2900 3598 2938
rect 3552 2866 3558 2900
rect 3592 2866 3598 2900
rect 3552 2828 3598 2866
rect 3552 2794 3558 2828
rect 3592 2794 3598 2828
rect 3552 2756 3598 2794
rect 3552 2722 3558 2756
rect 3592 2722 3598 2756
rect 3552 2684 3598 2722
rect 3552 2650 3558 2684
rect 3592 2650 3598 2684
rect 3552 2612 3598 2650
rect 3552 2578 3558 2612
rect 3592 2578 3598 2612
rect 3552 2540 3598 2578
rect 3552 2506 3558 2540
rect 3592 2506 3598 2540
rect 3552 2468 3598 2506
rect 3552 2434 3558 2468
rect 3592 2434 3598 2468
rect 3552 2396 3598 2434
rect 3552 2362 3558 2396
rect 3592 2362 3598 2396
rect 3552 2324 3598 2362
rect 3552 2290 3558 2324
rect 3592 2290 3598 2324
rect 3552 2252 3598 2290
rect 3552 2218 3558 2252
rect 3592 2218 3598 2252
rect 3552 2180 3598 2218
rect 3552 2146 3558 2180
rect 3592 2146 3598 2180
rect 3552 2108 3598 2146
rect 3552 2074 3558 2108
rect 3592 2074 3598 2108
rect 3552 2036 3598 2074
rect 3552 2002 3558 2036
rect 3592 2002 3598 2036
rect 3552 1964 3598 2002
rect 3552 1930 3558 1964
rect 3592 1930 3598 1964
rect 3552 1892 3598 1930
rect 3552 1858 3558 1892
rect 3592 1858 3598 1892
rect 3552 1811 3598 1858
rect 2736 1764 3542 1773
rect 2736 1730 3005 1764
rect 3039 1730 3163 1764
rect 3197 1730 3321 1764
rect 3355 1730 3479 1764
rect 3513 1730 3542 1764
rect 2736 1726 3542 1730
rect 2951 1718 3542 1726
rect 1894 1646 1940 1684
rect 1894 1612 1900 1646
rect 1934 1612 1940 1646
rect 1894 1574 1940 1612
rect 1894 1540 1900 1574
rect 1934 1540 1940 1574
rect 1894 1502 1940 1540
rect 1894 1468 1900 1502
rect 1934 1468 1940 1502
rect 1894 1430 1940 1468
rect 1894 1396 1900 1430
rect 1934 1396 1940 1430
rect 1894 1358 1940 1396
rect 1894 1324 1900 1358
rect 1934 1324 1940 1358
rect 1894 1286 1940 1324
rect 2187 1650 2235 1689
rect 2187 1616 2193 1650
rect 2227 1645 2235 1650
rect 2345 1650 2391 1689
rect 2227 1616 2233 1645
rect 2187 1578 2233 1616
rect 2187 1544 2193 1578
rect 2227 1544 2233 1578
rect 2187 1506 2233 1544
rect 2187 1472 2193 1506
rect 2227 1472 2233 1506
rect 2187 1434 2233 1472
rect 2187 1400 2193 1434
rect 2227 1400 2233 1434
rect 2187 1362 2233 1400
rect 2187 1328 2193 1362
rect 2227 1328 2233 1362
rect 2187 1289 2233 1328
rect 2345 1616 2351 1650
rect 2385 1616 2391 1650
rect 2345 1578 2391 1616
rect 2345 1544 2351 1578
rect 2385 1544 2391 1578
rect 2345 1506 2391 1544
rect 2345 1472 2351 1506
rect 2385 1472 2391 1506
rect 2345 1434 2391 1472
rect 2345 1400 2351 1434
rect 2385 1400 2391 1434
rect 2345 1362 2391 1400
rect 2345 1328 2351 1362
rect 2385 1328 2391 1362
rect 2345 1307 2391 1328
rect 2503 1654 2555 1689
rect 3574 1668 3699 1703
rect 2721 1662 2779 1668
rect 2503 1650 2549 1654
rect 2503 1616 2509 1650
rect 2543 1616 2549 1650
rect 2503 1578 2549 1616
rect 2503 1544 2509 1578
rect 2543 1544 2549 1578
rect 2584 1624 2636 1630
rect 2721 1628 2733 1662
rect 2767 1628 2779 1662
rect 2721 1623 2779 1628
rect 2636 1622 2779 1623
rect 3574 1634 3620 1668
rect 3654 1634 3699 1668
rect 2636 1573 2770 1622
rect 3574 1596 3699 1634
rect 2584 1566 2636 1572
rect 2503 1506 2549 1544
rect 2503 1472 2509 1506
rect 2543 1472 2549 1506
rect 2503 1434 2549 1472
rect 2503 1400 2509 1434
rect 2543 1400 2549 1434
rect 2503 1362 2549 1400
rect 2503 1328 2509 1362
rect 2543 1328 2549 1362
rect 1894 1252 1900 1286
rect 1934 1252 1940 1286
rect 1894 1214 1940 1252
rect 1894 1180 1900 1214
rect 1934 1180 1940 1214
rect 1894 1142 1940 1180
rect 1894 1108 1900 1142
rect 1934 1108 1940 1142
rect 1894 1070 1940 1108
rect 1894 1036 1900 1070
rect 1934 1036 1940 1070
rect 1894 998 1940 1036
rect 2343 1063 2393 1307
rect 2503 1289 2549 1328
rect 2730 1340 2770 1573
rect 2801 1563 2856 1575
rect 2970 1563 3561 1565
rect 2801 1558 3561 1563
rect 2801 1524 2811 1558
rect 2845 1550 3561 1558
rect 2845 1524 3010 1550
rect 2801 1520 3010 1524
rect 2801 1508 2856 1520
rect 2970 1516 3010 1520
rect 3044 1516 3168 1550
rect 3202 1516 3326 1550
rect 3360 1516 3484 1550
rect 3518 1516 3561 1550
rect 2970 1510 3561 1516
rect 2925 1435 2971 1478
rect 2925 1401 2931 1435
rect 2965 1401 2971 1435
rect 2925 1363 2971 1401
rect 2730 1300 2845 1340
rect 2343 1013 2551 1063
rect 2343 1009 2393 1013
rect 1894 965 1900 998
rect 1736 941 1782 964
rect 1892 964 1900 965
rect 1934 965 1940 998
rect 1934 964 1941 965
rect 1337 866 1625 915
rect 1285 859 1337 865
rect 1105 793 1151 831
rect 1576 846 1625 866
rect 1892 852 1941 964
rect 1576 797 1689 846
rect 1823 844 1941 852
rect 1823 810 1836 844
rect 1870 810 1941 844
rect 1823 803 1941 810
rect 1105 759 1111 793
rect 1145 759 1151 793
rect 1105 721 1151 759
rect 1373 724 1435 730
rect 1105 687 1111 721
rect 1145 687 1151 721
rect 1105 649 1151 687
rect 1367 719 1435 724
rect 1367 667 1373 719
rect 1425 667 1435 719
rect 1640 704 1689 797
rect 1829 796 1926 803
rect 1367 662 1435 667
rect 1373 656 1435 662
rect 1479 665 1525 704
rect 1105 615 1111 649
rect 1145 615 1151 649
rect 1105 577 1151 615
rect 1105 543 1111 577
rect 1145 543 1151 577
rect 1105 505 1151 543
rect 1105 471 1111 505
rect 1145 471 1151 505
rect 1105 433 1151 471
rect 1105 399 1111 433
rect 1145 399 1151 433
rect 1105 376 1151 399
rect 1479 631 1485 665
rect 1519 631 1525 665
rect 1479 593 1525 631
rect 1479 559 1485 593
rect 1519 559 1525 593
rect 1479 521 1525 559
rect 1479 487 1485 521
rect 1519 487 1525 521
rect 1479 449 1525 487
rect 1479 415 1485 449
rect 1519 415 1525 449
rect 1479 377 1525 415
rect 1479 358 1485 377
rect 1473 343 1485 358
rect 1519 343 1525 377
rect 1473 304 1525 343
rect 1637 672 1689 704
rect 1865 689 1926 796
rect 2365 712 2423 714
rect 2216 708 2423 712
rect 1637 665 1683 672
rect 1637 631 1643 665
rect 1677 631 1683 665
rect 1637 593 1683 631
rect 1637 559 1643 593
rect 1677 559 1683 593
rect 1637 521 1683 559
rect 1637 487 1643 521
rect 1677 487 1683 521
rect 1637 449 1683 487
rect 1637 415 1643 449
rect 1677 415 1683 449
rect 1637 377 1683 415
rect 1637 343 1643 377
rect 1677 343 1683 377
rect 1637 304 1683 343
rect 1875 665 1921 689
rect 1875 631 1881 665
rect 1915 631 1921 665
rect 1875 593 1921 631
rect 1875 559 1881 593
rect 1915 559 1921 593
rect 1875 521 1921 559
rect 1875 487 1881 521
rect 1915 487 1921 521
rect 1875 449 1921 487
rect 1875 415 1881 449
rect 1915 415 1921 449
rect 1875 377 1921 415
rect 1875 343 1881 377
rect 1915 343 1921 377
rect 1875 304 1921 343
rect 2033 665 2079 704
rect 2033 631 2039 665
rect 2073 631 2079 665
rect 2033 593 2079 631
rect 2033 559 2039 593
rect 2073 559 2079 593
rect 2033 521 2079 559
rect 2033 487 2039 521
rect 2073 487 2079 521
rect 2033 449 2079 487
rect 2033 415 2039 449
rect 2073 415 2079 449
rect 2033 377 2079 415
rect 2033 343 2039 377
rect 2073 343 2079 377
rect 2033 338 2079 343
rect 2216 674 2377 708
rect 2411 674 2423 708
rect 2216 669 2423 674
rect 2033 304 2112 338
rect 1291 217 1337 220
rect 1282 165 1288 217
rect 1340 165 1346 217
rect 1291 162 1337 165
rect -692 129 1251 157
rect 1473 150 1511 304
rect 2036 290 2112 304
rect 2216 290 2259 669
rect 2365 668 2423 669
rect 2036 247 2259 290
rect 2344 552 2390 591
rect 2344 518 2350 552
rect 2384 518 2390 552
rect 2501 552 2551 1013
rect 2501 538 2508 552
rect 2344 480 2390 518
rect 2344 446 2350 480
rect 2384 446 2390 480
rect 2344 408 2390 446
rect 2344 374 2350 408
rect 2384 374 2390 408
rect 2344 336 2390 374
rect 2344 302 2350 336
rect 2384 302 2390 336
rect 2344 264 2390 302
rect 2344 230 2350 264
rect 2384 230 2390 264
rect 2344 191 2390 230
rect 2502 518 2508 538
rect 2542 538 2551 552
rect 2660 552 2706 591
rect 2542 518 2548 538
rect 2502 480 2548 518
rect 2502 446 2508 480
rect 2542 446 2548 480
rect 2502 408 2548 446
rect 2502 374 2508 408
rect 2542 374 2548 408
rect 2502 336 2548 374
rect 2502 302 2508 336
rect 2542 302 2548 336
rect 2502 264 2548 302
rect 2502 230 2508 264
rect 2542 256 2548 264
rect 2660 518 2666 552
rect 2700 518 2706 552
rect 2660 480 2706 518
rect 2660 446 2666 480
rect 2700 446 2706 480
rect 2660 408 2706 446
rect 2660 374 2666 408
rect 2700 374 2706 408
rect 2660 336 2706 374
rect 2805 356 2845 1300
rect 2925 1329 2931 1363
rect 2965 1329 2971 1363
rect 2925 1291 2971 1329
rect 2925 1257 2931 1291
rect 2965 1257 2971 1291
rect 2925 1219 2971 1257
rect 2925 1185 2931 1219
rect 2965 1185 2971 1219
rect 2925 1147 2971 1185
rect 2925 1113 2931 1147
rect 2965 1113 2971 1147
rect 2925 1075 2971 1113
rect 2925 1041 2931 1075
rect 2965 1041 2971 1075
rect 2925 1003 2971 1041
rect 2925 969 2931 1003
rect 2965 969 2971 1003
rect 2925 931 2971 969
rect 2925 897 2931 931
rect 2965 897 2971 931
rect 2925 859 2971 897
rect 2925 825 2931 859
rect 2965 825 2971 859
rect 2925 787 2971 825
rect 2925 753 2931 787
rect 2965 753 2971 787
rect 2925 715 2971 753
rect 2925 681 2931 715
rect 2965 681 2971 715
rect 2925 643 2971 681
rect 2925 609 2931 643
rect 2965 609 2971 643
rect 2925 571 2971 609
rect 2925 537 2931 571
rect 2965 537 2971 571
rect 2925 499 2971 537
rect 2925 465 2931 499
rect 2965 465 2971 499
rect 2925 427 2971 465
rect 2925 393 2931 427
rect 2965 393 2971 427
rect 2660 302 2666 336
rect 2700 302 2706 336
rect 2793 347 2857 356
rect 2793 313 2808 347
rect 2842 313 2857 347
rect 2793 304 2857 313
rect 2925 355 2971 393
rect 2925 321 2931 355
rect 2965 321 2971 355
rect 2660 264 2706 302
rect 2542 230 2553 256
rect 2502 191 2553 230
rect 2660 230 2666 264
rect 2700 230 2706 264
rect 2925 287 2971 321
rect 3083 1435 3129 1478
rect 3083 1401 3089 1435
rect 3123 1401 3129 1435
rect 3083 1363 3129 1401
rect 3083 1329 3089 1363
rect 3123 1329 3129 1363
rect 3083 1291 3129 1329
rect 3083 1257 3089 1291
rect 3123 1257 3129 1291
rect 3083 1219 3129 1257
rect 3083 1185 3089 1219
rect 3123 1185 3129 1219
rect 3083 1147 3129 1185
rect 3083 1113 3089 1147
rect 3123 1113 3129 1147
rect 3083 1075 3129 1113
rect 3083 1041 3089 1075
rect 3123 1041 3129 1075
rect 3083 1003 3129 1041
rect 3083 969 3089 1003
rect 3123 969 3129 1003
rect 3083 931 3129 969
rect 3083 897 3089 931
rect 3123 897 3129 931
rect 3083 859 3129 897
rect 3083 825 3089 859
rect 3123 825 3129 859
rect 3083 787 3129 825
rect 3083 753 3089 787
rect 3123 753 3129 787
rect 3083 715 3129 753
rect 3083 681 3089 715
rect 3123 681 3129 715
rect 3083 643 3129 681
rect 3083 609 3089 643
rect 3123 609 3129 643
rect 3083 571 3129 609
rect 3083 537 3089 571
rect 3123 537 3129 571
rect 3083 499 3129 537
rect 3083 465 3089 499
rect 3123 465 3129 499
rect 3083 427 3129 465
rect 3083 393 3089 427
rect 3123 393 3129 427
rect 3083 355 3129 393
rect 3083 321 3089 355
rect 3123 321 3129 355
rect 2925 286 2972 287
rect 2925 255 2978 286
rect 3083 278 3129 321
rect 3241 1435 3287 1478
rect 3241 1401 3247 1435
rect 3281 1401 3287 1435
rect 3241 1363 3287 1401
rect 3241 1329 3247 1363
rect 3281 1329 3287 1363
rect 3241 1291 3287 1329
rect 3241 1257 3247 1291
rect 3281 1257 3287 1291
rect 3241 1219 3287 1257
rect 3241 1185 3247 1219
rect 3281 1185 3287 1219
rect 3241 1147 3287 1185
rect 3241 1113 3247 1147
rect 3281 1113 3287 1147
rect 3241 1075 3287 1113
rect 3241 1041 3247 1075
rect 3281 1041 3287 1075
rect 3241 1003 3287 1041
rect 3241 969 3247 1003
rect 3281 969 3287 1003
rect 3241 931 3287 969
rect 3241 897 3247 931
rect 3281 897 3287 931
rect 3241 859 3287 897
rect 3241 825 3247 859
rect 3281 825 3287 859
rect 3241 787 3287 825
rect 3241 753 3247 787
rect 3281 753 3287 787
rect 3241 715 3287 753
rect 3241 681 3247 715
rect 3281 681 3287 715
rect 3241 643 3287 681
rect 3241 609 3247 643
rect 3281 609 3287 643
rect 3241 571 3287 609
rect 3241 537 3247 571
rect 3281 537 3287 571
rect 3241 499 3287 537
rect 3241 465 3247 499
rect 3281 465 3287 499
rect 3241 427 3287 465
rect 3241 393 3247 427
rect 3281 393 3287 427
rect 3241 355 3287 393
rect 3241 321 3247 355
rect 3281 321 3287 355
rect 3241 320 3287 321
rect 3399 1435 3445 1478
rect 3399 1401 3405 1435
rect 3439 1401 3445 1435
rect 3399 1363 3445 1401
rect 3399 1329 3405 1363
rect 3439 1329 3445 1363
rect 3399 1291 3445 1329
rect 3399 1257 3405 1291
rect 3439 1257 3445 1291
rect 3399 1219 3445 1257
rect 3399 1185 3405 1219
rect 3439 1185 3445 1219
rect 3399 1147 3445 1185
rect 3399 1113 3405 1147
rect 3439 1113 3445 1147
rect 3399 1075 3445 1113
rect 3399 1041 3405 1075
rect 3439 1041 3445 1075
rect 3399 1003 3445 1041
rect 3399 969 3405 1003
rect 3439 969 3445 1003
rect 3399 931 3445 969
rect 3399 897 3405 931
rect 3439 897 3445 931
rect 3399 859 3445 897
rect 3399 825 3405 859
rect 3439 825 3445 859
rect 3399 787 3445 825
rect 3399 753 3405 787
rect 3439 753 3445 787
rect 3399 715 3445 753
rect 3399 681 3405 715
rect 3439 681 3445 715
rect 3399 643 3445 681
rect 3399 609 3405 643
rect 3439 609 3445 643
rect 3399 571 3445 609
rect 3399 537 3405 571
rect 3439 537 3445 571
rect 3399 499 3445 537
rect 3399 465 3405 499
rect 3439 465 3445 499
rect 3399 427 3445 465
rect 3399 393 3405 427
rect 3439 393 3445 427
rect 3399 355 3445 393
rect 3399 321 3405 355
rect 3439 321 3445 355
rect 3241 278 3292 320
rect 3399 278 3445 321
rect 3557 1435 3603 1478
rect 3557 1401 3563 1435
rect 3597 1401 3603 1435
rect 3557 1363 3603 1401
rect 3557 1329 3563 1363
rect 3597 1329 3603 1363
rect 3557 1291 3603 1329
rect 3557 1257 3563 1291
rect 3597 1257 3603 1291
rect 3557 1219 3603 1257
rect 3557 1185 3563 1219
rect 3597 1185 3603 1219
rect 3557 1147 3603 1185
rect 3557 1113 3563 1147
rect 3597 1113 3603 1147
rect 3557 1075 3603 1113
rect 3557 1041 3563 1075
rect 3597 1041 3603 1075
rect 3557 1003 3603 1041
rect 3557 969 3563 1003
rect 3597 969 3603 1003
rect 3557 931 3603 969
rect 3557 897 3563 931
rect 3597 897 3603 931
rect 3557 859 3603 897
rect 3557 825 3563 859
rect 3597 825 3603 859
rect 3557 787 3603 825
rect 3557 753 3563 787
rect 3597 753 3603 787
rect 3557 715 3603 753
rect 3557 681 3563 715
rect 3597 681 3603 715
rect 3557 643 3603 681
rect 3557 609 3563 643
rect 3597 609 3603 643
rect 3557 571 3603 609
rect 3557 537 3563 571
rect 3597 537 3603 571
rect 3557 499 3603 537
rect 3557 465 3563 499
rect 3597 465 3603 499
rect 3557 427 3603 465
rect 3557 393 3563 427
rect 3597 393 3603 427
rect 3557 355 3603 393
rect 3557 321 3563 355
rect 3597 335 3603 355
rect 3597 321 3607 335
rect 3557 278 3607 321
rect 2660 191 2706 230
rect 2932 201 2978 255
rect 3246 201 3292 278
rect 3561 201 3607 278
rect 2348 150 2386 191
rect -692 99 1260 129
rect 1473 112 2386 150
rect -692 65 -595 99
rect -561 95 757 99
rect -561 89 72 95
rect -561 65 -271 89
rect -692 55 -271 65
rect -237 85 72 89
rect -237 55 -49 85
rect -692 51 -49 55
rect -15 61 72 85
rect 106 93 578 95
rect 106 61 240 93
rect -15 59 240 61
rect 274 59 409 93
rect 443 61 578 93
rect 612 65 757 95
rect 791 65 944 99
rect 978 97 1260 99
rect 978 65 1145 97
rect 612 63 1145 65
rect 1179 75 1260 97
rect 2507 75 2553 191
rect 2932 155 3607 201
rect 2932 75 2978 155
rect 1179 63 2978 75
rect 612 61 2978 63
rect 443 59 2978 61
rect -15 51 2978 59
rect -692 29 2978 51
rect -692 0 1260 29
rect -692 -4 66 0
<< via1 >>
rect 3074 3872 3126 3924
rect 2832 3620 2884 3672
rect 1862 2347 1914 2399
rect 1784 1931 1836 1983
rect 835 1402 887 1454
rect 1408 1572 1460 1624
rect 1360 1443 1412 1453
rect 1360 1409 1368 1443
rect 1368 1409 1402 1443
rect 1402 1409 1412 1443
rect 1360 1401 1412 1409
rect 840 1141 892 1193
rect 618 711 670 719
rect 618 677 627 711
rect 627 677 661 711
rect 661 677 670 711
rect 618 667 670 677
rect 676 340 728 349
rect 676 306 682 340
rect 682 306 716 340
rect 716 306 728 340
rect 676 297 728 306
rect 1285 865 1337 917
rect 2584 1572 2636 1624
rect 1373 710 1425 719
rect 1373 676 1387 710
rect 1387 676 1421 710
rect 1421 676 1425 710
rect 1373 667 1425 676
rect 1288 208 1340 217
rect 1288 174 1297 208
rect 1297 174 1331 208
rect 1331 174 1340 208
rect 1288 165 1340 174
<< metal2 >>
rect 3074 3924 3126 3930
rect 2833 3874 3074 3923
rect 2833 3678 2882 3874
rect 3074 3866 3126 3872
rect 2832 3672 2884 3678
rect 2832 3614 2884 3620
rect 1862 2399 1914 2405
rect 1788 2351 1862 2395
rect 1788 1983 1832 2351
rect 1862 2341 1914 2347
rect 1778 1931 1784 1983
rect 1836 1931 1842 1983
rect 1408 1624 1460 1630
rect 1405 1573 1408 1623
rect 2576 1623 2584 1624
rect 1460 1573 2584 1623
rect 2576 1572 2584 1573
rect 2636 1572 2642 1624
rect 1408 1566 1460 1572
rect 829 1402 835 1454
rect 887 1447 893 1454
rect 1360 1453 1412 1459
rect 887 1408 1360 1447
rect 887 1402 893 1408
rect 1360 1395 1412 1401
rect 840 1193 892 1199
rect 892 1189 1328 1191
rect 892 1142 1336 1189
rect 840 1135 892 1141
rect 1287 917 1336 1142
rect 1279 865 1285 917
rect 1337 865 1343 917
rect 618 719 670 725
rect 1373 719 1425 730
rect 670 668 1373 718
rect 618 661 670 667
rect 1373 656 1425 667
rect 670 297 676 349
rect 728 297 734 349
rect 685 208 719 297
rect 1288 217 1340 223
rect 685 179 1288 208
rect 759 174 1288 179
rect 1288 159 1340 165
<< labels >>
flabel metal1 s 1627 3894 1627 3894 0 FreeSans 3906 0 0 0 VDD
flabel metal1 s 3680 1652 3680 1652 0 FreeSans 3906 0 0 0 OUT
flabel metal1 s 976 79 976 79 0 FreeSans 3906 0 0 0 GND
flabel metal1 s 116 974 116 974 0 FreeSans 2500 0 0 0 VIN
<< end >>
