magic
tech sky130A
magscale 1 2
timestamp 1686021299
<< metal1 >>
rect 4911 2416 4963 2422
rect 4963 2375 6897 2405
rect 4911 2358 4963 2364
rect 6744 2327 6750 2334
rect 6398 2288 6750 2327
rect 6744 2282 6750 2288
rect 6802 2282 6808 2334
rect 6867 2293 6897 2375
rect 4993 1797 4999 1849
rect 5051 1842 5057 1849
rect 5051 1803 5483 1842
rect 5051 1797 5057 1803
rect 4993 1343 4999 1395
rect 5051 1388 5057 1395
rect 5051 1349 5454 1388
rect 6228 1376 6818 1404
rect 5051 1343 5057 1349
rect 4917 1225 4969 1231
rect 6228 1213 6256 1376
rect 4969 1185 6256 1213
rect 4917 1167 4969 1173
<< via1 >>
rect 4911 2364 4963 2416
rect 6750 2282 6802 2334
rect 4999 1797 5051 1849
rect 4999 1343 5051 1395
rect 4917 1173 4969 1225
<< metal2 >>
rect 156 2333 211 2456
rect 260 2327 315 2456
rect 3446 2306 3487 2456
rect 4905 2364 4911 2416
rect 4963 2364 4969 2416
rect 4918 2289 4957 2364
rect 5004 2315 5045 2456
rect 5164 2328 5205 2456
rect 5244 2328 5285 2456
rect 5324 2315 5365 2456
rect 5404 2328 5445 2456
rect 6750 2334 6802 2340
rect 6802 2289 7029 2328
rect 6750 2276 6802 2282
rect -76 2234 -8 2243
rect -76 1028 -8 2166
rect 4999 1849 5051 1855
rect 4999 1791 5051 1797
rect 5084 1631 5125 1787
rect 5164 1642 5205 1796
rect 5244 1624 5285 1793
rect 5324 1650 5365 1793
rect 5404 1640 5445 1793
rect -76 951 -8 960
rect 26 1558 94 1567
rect 26 322 94 1490
rect 5004 1401 5045 1431
rect 4999 1395 5051 1401
rect 4999 1337 5051 1343
rect 5004 1272 5045 1337
rect 4911 1173 4917 1225
rect 4969 1173 4975 1225
rect 4929 1061 4957 1173
rect 26 245 94 254
rect 159 0 214 91
rect 260 0 315 91
rect 3446 0 3487 116
<< via2 >>
rect -76 2166 -8 2234
rect -76 960 -8 1028
rect 26 1490 94 1558
rect 26 254 94 322
<< metal3 >>
rect -118 2234 140 2278
rect -118 2166 -76 2234
rect -8 2166 140 2234
rect -118 2138 140 2166
rect -118 1558 196 1588
rect -118 1490 26 1558
rect 94 1490 196 1558
rect -118 1448 196 1490
rect -118 1028 186 1050
rect -118 960 -76 1028
rect -8 960 186 1028
rect -118 910 186 960
rect -118 322 184 360
rect -118 254 26 322
rect 94 254 184 322
rect -118 220 184 254
use 2_bit_dac  2_bit_dac_0
array 0 0 5006 0 1 1228
timestamp 1685863011
transform 1 0 408 0 1 182
box -408 -182 4598 1046
use switch_n_3v3  switch_n_3v3_1
timestamp 1686019770
transform 1 0 11886 0 1 2132
box -6932 -991 -4922 237
<< labels >>
rlabel metal3 -100 2234 -100 2234 7 VCC
rlabel metal3 -92 1522 -92 1522 7 VSS
rlabel metal2 184 2430 184 2430 7 D0
rlabel metal2 288 2432 288 2432 7 VREFL
rlabel metal2 186 20 186 20 7 D0_BUF
rlabel metal2 282 12 282 12 7 VREFH
rlabel metal2 3468 2450 3468 2450 7 D1
rlabel metal2 3468 12 3468 12 7 D1_BUF
rlabel metal2 5023 2436 5023 2436 7 D2
rlabel metal2 5023 1290 5023 1290 7 D2_BUF
rlabel metal2 7021 2310 7021 2310 7 VOUT
<< end >>
