magic
tech sky130A
magscale 1 2
timestamp 1687539450
<< metal1 >>
rect 6968 10970 6974 11022
rect 7026 10970 7032 11022
rect 6829 10923 6835 10930
rect 6516 10884 6835 10923
rect 6829 10878 6835 10884
rect 6887 10878 6893 10930
rect 6985 10889 7015 10970
rect 5350 10393 5356 10445
rect 5408 10438 5414 10445
rect 5408 10399 5627 10438
rect 5408 10393 5414 10399
rect 7079 9998 7085 10010
rect 5348 9939 5354 9991
rect 5406 9984 5412 9991
rect 5406 9945 5603 9984
rect 6908 9970 7085 9998
rect 7079 9958 7085 9970
rect 7137 9958 7143 10010
rect 5406 9939 5412 9945
<< via1 >>
rect 6974 10970 7026 11022
rect 6835 10878 6887 10930
rect 5356 10393 5408 10445
rect 5354 9939 5406 9991
rect 7085 9958 7137 10010
<< metal2 >>
rect 274 19481 329 19646
rect 378 19471 433 19648
rect 3564 19508 3605 19648
rect 5122 19510 5163 19648
rect 5202 19496 5243 19648
rect 5282 19508 5323 19648
rect 5362 19510 5403 19648
rect 7154 14887 7337 14926
rect 42 9320 110 10974
rect 5122 10923 5164 11015
rect 5202 10923 5244 11027
rect 6974 11022 7026 11028
rect 5282 10915 5324 11009
rect 5362 10929 5404 11008
rect 5442 10923 5484 11008
rect 5522 10917 5564 11008
rect 7298 11011 7337 14887
rect 7026 10981 7337 11011
rect 6974 10964 7026 10970
rect 6835 10930 6887 10936
rect 6887 10885 7150 10924
rect 6835 10872 6887 10878
rect 7111 10802 7150 10885
rect 7111 10763 7360 10802
rect 5356 10445 5408 10451
rect 144 8690 212 10332
rect 5122 10218 5163 10389
rect 5202 10222 5243 10389
rect 5282 10242 5323 10389
rect 5356 10387 5408 10393
rect 5442 10222 5483 10389
rect 5522 10232 5563 10389
rect 7085 10010 7137 10016
rect 5354 9991 5406 9997
rect 7137 9970 7322 9998
rect 7085 9952 7137 9958
rect 5354 9933 5406 9939
rect 5122 9689 5164 9825
rect 5202 9683 5244 9815
rect 5282 9697 5324 9829
rect 5362 9675 5404 9825
rect 5442 9699 5484 9827
rect 5522 9689 5564 9827
rect 7283 5102 7322 9970
rect 7154 5063 7322 5102
rect 5122 1272 5163 1404
rect 5202 1272 5243 1394
rect 5282 1272 5323 1356
rect 5362 1272 5403 1374
rect 277 0 332 225
rect 378 0 433 211
rect 3564 0 3605 92
use 5_bit_dac  5_bit_dac_0
array 0 0 7252 0 1 9824
timestamp 1687539450
transform 1 0 0 0 1 0
box -2 0 7724 9824
use switch_n_3v3  switch_n_3v3_0
timestamp 1687539450
transform 1 0 12004 0 1 10728
box -6932 -990 -4922 236
<< labels >>
rlabel metal2 82 9906 82 9906 3 VCC
rlabel metal2 180 9904 180 9904 3 VSS
rlabel metal2 290 19592 290 19592 3 D0
rlabel metal2 392 19600 392 19600 3 VREFL
rlabel metal2 3576 19606 3576 19606 3 D1
rlabel metal2 5136 19622 5136 19622 3 D2
rlabel metal2 5230 19628 5230 19628 3 D3
rlabel metal2 5310 19634 5310 19634 3 D4
rlabel metal2 5386 19634 5386 19634 3 D5
rlabel metal2 282 42 282 42 3 D0_BUF
rlabel metal2 418 36 418 36 3 VREFH
rlabel metal2 3588 24 3588 24 3 D1_BUF
rlabel metal2 5128 1298 5128 1298 3 D2_BUF
rlabel metal2 5210 1312 5210 1312 3 D3_BUF
rlabel metal2 5288 1292 5288 1292 3 D4_BUF
rlabel metal2 5374 1294 5374 1294 3 D5_BUF
rlabel metal2 7344 10781 7344 10781 3 VOUT
<< end >>
