* SPICE3 file created from 7_bit_dac.ext - technology: sky130A

.subckt x7_bit_dac VCC VSS D0 VREFL D1 D2 D3 D4 D5 D6 D0_BUF VREFH D1_BUF D2_BUF D3_BUF
+ D4_BUF D5_BUF D6_BUF VOUT
X0 6_bit_dac_0[0]/VOUT D5_BUF 6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X1 6_bit_dac_0[0]/switch_n_3v3_0/DX_ switch_n_3v3_1/D5 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X2 D5_BUF 6_bit_dac_0[0]/switch_n_3v3_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X3 6_bit_dac_0[0]/VOUT D5_BUF 6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X4 6_bit_dac_0[0]/switch_n_3v3_0/DX_ switch_n_3v3_1/D5 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X5 6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/switch_n_3v3_0/DX_ 6_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6 D5_BUF 6_bit_dac_0[0]/switch_n_3v3_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X7 6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/switch_n_3v3_0/DX_ 6_bit_dac_0[0]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X8 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT D1_BUF 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X9 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X10 D1_BUF 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X11 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT D1_BUF 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X12 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X13 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X14 D1_BUF 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X15 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X16 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X17 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH D0_BUF 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X18 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X19 D0_BUF 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X20 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH D0_BUF 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X21 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X22 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X23 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X24 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X25 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H D0_BUF 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X26 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X27 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X28 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L D0_BUF 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X29 D0_BUF 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X30 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X31 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X32 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X33 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=55.1 ps=490 w=1 l=0.5
X34 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X35 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X36 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=27.5 ps=300 w=0.5 l=0.5
X37 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X38 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X39 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X40 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X41 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X42 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X43 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X44 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X45 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X46 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X47 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X48 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X49 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X50 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X51 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X52 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X53 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X54 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X55 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X56 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT D2_BUF 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X57 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X58 D2_BUF 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X59 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT D2_BUF 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X60 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X61 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X62 D2_BUF 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X63 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X64 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X65 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X66 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X67 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X68 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X69 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X70 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X71 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X72 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X73 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X74 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X75 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X76 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X77 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X78 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X79 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X80 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X81 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X82 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X83 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X84 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X85 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X86 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X87 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X88 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X89 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X90 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X91 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X92 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X93 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X94 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X95 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X96 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X97 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X98 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X99 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X100 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X101 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X102 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X103 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X104 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X105 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X106 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X107 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X108 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X109 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X110 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X111 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X112 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X113 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X114 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X115 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X116 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X117 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X118 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X119 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X120 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT D3_BUF 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X121 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X122 D3_BUF 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X123 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT D3_BUF 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X124 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X125 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X126 D3_BUF 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X127 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X128 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X129 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X130 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X131 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X132 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X133 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X134 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X135 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X136 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X137 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X138 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X139 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X140 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X141 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X142 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X143 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X144 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X145 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X146 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X147 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X148 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X149 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X150 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X151 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X152 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X153 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X154 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X155 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X156 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X157 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X158 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X159 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X160 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X161 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X162 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X163 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X164 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X165 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X166 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X167 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X168 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X169 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X170 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X171 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X172 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X173 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X174 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X175 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X176 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X177 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X178 6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X179 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X180 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X181 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X182 6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D2 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X183 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X184 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X185 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X186 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X187 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X188 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X189 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X190 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X191 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X192 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X193 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X194 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X195 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X196 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X197 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X198 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X199 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X200 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X201 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X202 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X203 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X204 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X205 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X206 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X207 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X208 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X209 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X210 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X211 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X212 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/D1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X213 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X214 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X215 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X216 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X217 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X218 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X219 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X220 6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X221 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X222 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X223 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X224 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X225 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X226 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X227 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X228 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X229 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X230 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/D0 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X231 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X232 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X233 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 6_bit_dac_0[0]/switch_n_3v3_0/D2 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X234 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X235 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X236 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 6_bit_dac_0[0]/switch_n_3v3_0/D2 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X237 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X238 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X239 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X240 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X241 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 6_bit_dac_0[0]/switch_n_3v3_0/D3 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X242 6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X243 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X244 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 6_bit_dac_0[0]/switch_n_3v3_0/D3 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X245 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X246 6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/D3 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X247 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X248 6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT D4_BUF 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X249 6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 6_bit_dac_0[0]/switch_n_3v3_0/D4 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X250 D4_BUF 6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X251 6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT D4_BUF 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X252 6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 6_bit_dac_0[0]/switch_n_3v3_0/D4 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X253 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X254 D4_BUF 6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X255 6_bit_dac_0[0]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[0]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X256 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X257 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X258 6_bit_dac_0[0]/5_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X259 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X260 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X261 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X262 6_bit_dac_0[0]/5_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X263 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X264 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X265 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X266 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X267 6_bit_dac_0[0]/5_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X268 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 6_bit_dac_0[0]/5_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X269 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X270 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X271 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X272 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X273 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 6_bit_dac_0[0]/5_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X274 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X275 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X276 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 6_bit_dac_0[0]/5_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X277 6_bit_dac_0[0]/5_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X278 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X279 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X280 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X281 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X282 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X283 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X284 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X285 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X286 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X287 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X288 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X289 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X290 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X291 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X292 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X293 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X294 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X295 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X296 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X297 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X298 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X299 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X300 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X301 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X302 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X303 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X304 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/switch_n_3v3_0/D2 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X305 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X306 6_bit_dac_0[0]/switch_n_3v3_0/D2 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X307 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/switch_n_3v3_0/D2 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X308 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X309 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X310 6_bit_dac_0[0]/switch_n_3v3_0/D2 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X311 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X312 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X313 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X314 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X315 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X316 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X317 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X318 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X319 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X320 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X321 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X322 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X323 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X324 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X325 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X326 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X327 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X328 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X329 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X330 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X331 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X332 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X333 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X334 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X335 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X336 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X337 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X338 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X339 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X340 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X341 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X342 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X343 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X344 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X345 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X346 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X347 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X348 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X349 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X350 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X351 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X352 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X353 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X354 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X355 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X356 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X357 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X358 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X359 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X360 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X361 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X362 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X363 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X364 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X365 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X366 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X367 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X368 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/switch_n_3v3_0/D3 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X369 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X370 6_bit_dac_0[0]/switch_n_3v3_0/D3 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X371 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/switch_n_3v3_0/D3 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X372 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X373 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X374 6_bit_dac_0[0]/switch_n_3v3_0/D3 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X375 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X376 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X377 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X378 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X379 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X380 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X381 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X382 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X383 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X384 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X385 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X386 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X387 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X388 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X389 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X390 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X391 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X392 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X393 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X394 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X395 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X396 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X397 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X398 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X399 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X400 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X401 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X402 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X403 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X404 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X405 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X406 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X407 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X408 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X409 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X410 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X411 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X412 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X413 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X414 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X415 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X416 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X417 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X418 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X419 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X420 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X421 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X422 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X423 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X424 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X425 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X426 6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X427 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X428 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X429 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X430 6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D2 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X431 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X432 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X433 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X434 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X435 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X436 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X437 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X438 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X439 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X440 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X441 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X442 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X443 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X444 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X445 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X446 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X447 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X448 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X449 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X450 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X451 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X452 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X453 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X454 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X455 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X456 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X457 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/D1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X458 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X459 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X460 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/D1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X461 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X462 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X463 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X464 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X465 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X466 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X467 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X468 6_bit_dac_0[1]/VREFH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X469 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X470 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/D0 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X471 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X472 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X473 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X474 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X475 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 6_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X476 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X477 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X478 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/D0 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X479 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X480 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X481 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ switch_n_3v3_1/D2 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X482 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X483 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X484 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ switch_n_3v3_1/D2 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X485 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X486 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X487 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X488 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X489 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ switch_n_3v3_1/D3 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X490 6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X491 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X492 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ switch_n_3v3_1/D3 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X493 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X494 6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/D3 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X495 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X496 6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/switch_n_3v3_0/D4 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X497 6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ switch_n_3v3_1/D4 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X498 6_bit_dac_0[0]/switch_n_3v3_0/D4 6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X499 6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/switch_n_3v3_0/D4 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X500 6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ switch_n_3v3_1/D4 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X501 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X502 6_bit_dac_0[0]/switch_n_3v3_0/D4 6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X503 6_bit_dac_0[0]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 6_bit_dac_0[0]/5_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X504 6_bit_dac_0[1]/VOUT switch_n_3v3_1/D5 6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X505 6_bit_dac_0[1]/switch_n_3v3_0/DX_ D5 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X506 switch_n_3v3_1/D5 6_bit_dac_0[1]/switch_n_3v3_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X507 6_bit_dac_0[1]/VOUT switch_n_3v3_1/D5 6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X508 6_bit_dac_0[1]/switch_n_3v3_0/DX_ D5 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X509 6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/switch_n_3v3_0/DX_ 6_bit_dac_0[1]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X510 switch_n_3v3_1/D5 6_bit_dac_0[1]/switch_n_3v3_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X511 6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/switch_n_3v3_0/DX_ 6_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X512 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X513 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X514 6_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X515 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X516 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X517 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X518 6_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X519 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X520 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X521 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X522 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X523 6_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X524 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 6_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X525 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X526 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X527 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X528 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X529 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 6_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X530 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X531 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X532 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 6_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X533 6_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X534 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X535 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X536 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X537 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X538 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X539 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X540 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X541 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X542 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X543 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X544 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X545 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X546 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X547 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X548 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X549 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X550 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X551 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X552 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X553 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X554 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X555 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X556 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X557 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X558 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X559 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X560 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT switch_n_3v3_1/D2 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X561 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X562 switch_n_3v3_1/D2 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X563 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT switch_n_3v3_1/D2 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X564 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X565 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X566 switch_n_3v3_1/D2 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X567 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X568 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X569 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X570 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X571 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X572 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X573 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X574 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X575 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X576 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X577 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X578 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X579 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X580 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X581 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X582 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X583 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X584 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X585 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X586 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X587 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X588 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X589 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X590 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X591 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X592 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X593 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X594 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X595 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X596 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X597 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X598 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X599 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X600 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X601 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X602 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X603 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X604 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X605 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X606 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X607 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X608 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X609 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X610 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X611 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X612 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X613 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X614 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X615 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X616 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X617 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X618 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X619 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X620 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X621 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X622 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/D2 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X623 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X624 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT switch_n_3v3_1/D3 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X625 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X626 switch_n_3v3_1/D3 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X627 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT switch_n_3v3_1/D3 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X628 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X629 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X630 switch_n_3v3_1/D3 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X631 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X632 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X633 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X634 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X635 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X636 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X637 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X638 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X639 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X640 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X641 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X642 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X643 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X644 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X645 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X646 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X647 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X648 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X649 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X650 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X651 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X652 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X653 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X654 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X655 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X656 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X657 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X658 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X659 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X660 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X661 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X662 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X663 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X664 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X665 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X666 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X667 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X668 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X669 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X670 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X671 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X672 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X673 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X674 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X675 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X676 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X677 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X678 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X679 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X680 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X681 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X682 6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X683 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X684 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X685 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X686 6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D2 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X687 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X688 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X689 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X690 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X691 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X692 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X693 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X694 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X695 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X696 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X697 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X698 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X699 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X700 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X701 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X702 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X703 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X704 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X705 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X706 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X707 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X708 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X709 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X710 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X711 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X712 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X713 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X714 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X715 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X716 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/D1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X717 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X718 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X719 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X720 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X721 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X722 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X723 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X724 6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X725 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X726 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X727 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X728 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X729 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X730 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X731 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X732 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X733 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X734 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/D0 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X735 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X736 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X737 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 6_bit_dac_0[1]/switch_n_3v3_0/D2 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X738 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X739 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X740 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 6_bit_dac_0[1]/switch_n_3v3_0/D2 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X741 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X742 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/D2 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X743 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X744 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X745 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 6_bit_dac_0[1]/switch_n_3v3_0/D3 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X746 6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X747 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X748 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 6_bit_dac_0[1]/switch_n_3v3_0/D3 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X749 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X750 6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/D3 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X751 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X752 6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT switch_n_3v3_1/D4 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X753 6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 6_bit_dac_0[1]/switch_n_3v3_0/D4 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X754 switch_n_3v3_1/D4 6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X755 6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT switch_n_3v3_1/D4 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X756 6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 6_bit_dac_0[1]/switch_n_3v3_0/D4 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X757 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X758 switch_n_3v3_1/D4 6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X759 6_bit_dac_0[1]/5_bit_dac_0[0]/4_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/switch_n_3v3_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[0]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X760 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X761 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X762 6_bit_dac_0[1]/5_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X763 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X764 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X765 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X766 6_bit_dac_0[1]/5_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X767 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X768 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X769 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X770 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X771 6_bit_dac_0[1]/5_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X772 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 6_bit_dac_0[1]/5_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X773 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X774 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X775 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X776 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X777 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 6_bit_dac_0[1]/5_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X778 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X779 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X780 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 6_bit_dac_0[1]/5_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X781 6_bit_dac_0[1]/5_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X782 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X783 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X784 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X785 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X786 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X787 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X788 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X789 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X790 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X791 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X792 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X793 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X794 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X795 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X796 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X797 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X798 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X799 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X800 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X801 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X802 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X803 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X804 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X805 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X806 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X807 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X808 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/switch_n_3v3_0/D2 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X809 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X810 6_bit_dac_0[1]/switch_n_3v3_0/D2 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X811 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/switch_n_3v3_0/D2 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X812 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X813 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X814 6_bit_dac_0[1]/switch_n_3v3_0/D2 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X815 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X816 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X817 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X818 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X819 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X820 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X821 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X822 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X823 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X824 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X825 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X826 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X827 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X828 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X829 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X830 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X831 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X832 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X833 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X834 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X835 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X836 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X837 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X838 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X839 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X840 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X841 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X842 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X843 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X844 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X845 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X846 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X847 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X848 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X849 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X850 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X851 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X852 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X853 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X854 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X855 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X856 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X857 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X858 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X859 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X860 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X861 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X862 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X863 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X864 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X865 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X866 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X867 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X868 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X869 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X870 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/D2 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X871 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X872 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/switch_n_3v3_0/D3 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X873 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X874 6_bit_dac_0[1]/switch_n_3v3_0/D3 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X875 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/switch_n_3v3_0/D3 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X876 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X877 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X878 6_bit_dac_0[1]/switch_n_3v3_0/D3 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X879 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/3_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/switch_n_3v3_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X880 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X881 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X882 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X883 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X884 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X885 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X886 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X887 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X888 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X889 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X890 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X891 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X892 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X893 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X894 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X895 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X896 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X897 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X898 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X899 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X900 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X901 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X902 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X903 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X904 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X905 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X906 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X907 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X908 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X909 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X910 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X911 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X912 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X913 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X914 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X915 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X916 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X917 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X918 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X919 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X920 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X921 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X922 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X923 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X924 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X925 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X926 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X927 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X928 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X929 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X930 6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X931 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X932 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X933 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X934 6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D2 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X935 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/switch_n_3v3_1/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X936 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X937 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X938 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X939 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X940 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X941 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X942 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X943 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X944 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X945 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X946 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X947 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X948 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X949 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X950 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X951 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X952 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X953 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X954 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_H 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X955 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X956 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X957 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X958 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X959 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/switch2n_3v3_0/R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X960 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0.435 ps=4.74 w=0.5 l=0.5
X961 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ D1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X962 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X963 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0.87 ps=7.74 w=1 l=0.5
X964 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ D1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X965 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X966 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D1 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X967 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch_n_3v3_v2_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X968 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X969 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X970 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X971 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X972 VREFL 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X973 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VREFH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VREFH VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X974 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# D0 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X975 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VREFL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.361 ps=3.45 w=0.5 l=0.5
X976 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.578 ps=5.32 w=0.5 l=0.5
X977 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X978 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_H 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X979 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VREFL VSS sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X980 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.578 pd=5.32 as=0 ps=0 w=0.5 l=0.5
X981 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/D0 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X982 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# D0 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X983 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/VOUTL 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/a_n6524_n498# 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/switch2n_3v3_0/R_L VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X984 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X985 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ D2 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X986 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X987 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X988 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ D2 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X989 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X990 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/D2 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X991 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/2_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/switch_n_3v3_1/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X992 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.435 pd=4.74 as=0 ps=0 w=0.5 l=0.5
X993 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ D3 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X994 6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X995 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
X996 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ D3 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X997 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X998 6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/D3 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X999 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/3_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/switch_n_3v3_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1000 6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/switch_n_3v3_0/D4 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1001 6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ D4 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1002 6_bit_dac_0[1]/switch_n_3v3_0/D4 6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1003 6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/switch_n_3v3_0/D4 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1004 6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ D4 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1005 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[1]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1006 6_bit_dac_0[1]/switch_n_3v3_0/D4 6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1007 6_bit_dac_0[1]/5_bit_dac_0[1]/4_bit_dac_0[0]/VOUT 6_bit_dac_0[1]/5_bit_dac_0[1]/switch_n_3v3_0/DX_ 6_bit_dac_0[1]/5_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X1008 VOUT D6_BUF 6_bit_dac_0[0]/VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=3.16 as=0.435 ps=4.74 w=0.5 l=0.5
X1009 switch_n_3v3_1/DX_ D6 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1010 D6_BUF switch_n_3v3_1/DX_ VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X1011 VOUT D6_BUF 6_bit_dac_0[1]/VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.5
X1012 switch_n_3v3_1/DX_ D6 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1013 6_bit_dac_0[1]/VOUT switch_n_3v3_1/DX_ VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=0.5 l=0.5
X1014 D6_BUF switch_n_3v3_1/DX_ VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0 ps=0 w=0.5 l=0.5
X1015 6_bit_dac_0[0]/VOUT switch_n_3v3_1/DX_ VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.87 pd=7.74 as=0 ps=0 w=1 l=0.5
.ends

X1 VCC VSS D0 VREFL D1 D2 D3 D4 D5 D6 D0_BUF VREFH D1_BUF D2_BUF D3_BUF D4_BUF D5_BUF D6_BUF VOUT x7_bit_dac
   
.param mc_mm_switch=0
.param mc_pr_switch=0
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /foss/pdks/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice


V1 VSS 0 dc 0
V2 VCC 0 dc 3.3

V3 VREFH 0 dc 3.3
V4 VREFL 0 dc 0

V5 D0 0 PULSE(0 1.8 0 1n 1n 1u 2u)
V6 D1 0 PULSE(0 1.8 0 1n 1n 2u 4u)
V7 D2 0 PULSE(0 1.8 0 1n 1n 4u 8u)
V8 D3 0 PULSE(0 1.8 0 1n 1n 8u 16u)
V9 D4 0 PULSE(0 1.8 0 1n 1n 16u 32u)
V10 D5 0 PULSE(0 1.8 0 1n 1n 32u 64u)
V11 D6 0 PULSE(0 1.8 0 1n 1n 64u 128u)

.tran 1u 130u
.control
run
plot VOUT
.endc
.end
