VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO 8_bit_dac_tx_buffer
  CLASS BLOCK ;
  FOREIGN 8_bit_dac_tx_buffer ;
  ORIGIN 12.045 0.900 ;
  SIZE 53.005 BY 429.140 ;
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -8.320 404.855 -8.150 428.240 ;
    END
  END D0
  OBS
      LAYER li1 ;
        RECT -12.045 -0.900 40.960 426.835 ;
      LAYER met1 ;
        RECT -10.635 -0.595 39.285 427.540 ;
      LAYER met2 ;
        RECT -11.255 404.575 -8.600 428.240 ;
        RECT -7.870 404.575 40.250 428.240 ;
        RECT -11.255 -0.555 40.250 404.575 ;
      LAYER met3 ;
        RECT -12.045 1.100 40.960 426.740 ;
  END
END 8_bit_dac_tx_buffer
END LIBRARY

