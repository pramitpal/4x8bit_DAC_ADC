magic
tech sky130A
magscale 1 2
timestamp 1686726141
<< viali >>
rect 0 0 140 140
<< metal1 >>
rect -6 146 146 152
rect -12 -6 -6 146
rect 134 140 146 146
rect 140 0 146 140
rect 134 -6 146 0
rect -6 -12 146 -6
<< via1 >>
rect -6 140 134 146
rect -6 0 0 140
rect 0 0 134 140
rect -6 -6 134 0
<< metal2 >>
rect 745 85774 779 86800
rect 848 85794 882 86800
rect 946 85794 980 86800
rect 1050 85794 1084 86800
rect 1158 85793 1192 86800
rect 1258 85785 1292 86800
rect 1366 85794 1400 86800
rect 1478 85782 1512 86800
rect 9265 85699 9373 86800
rect 11346 85794 11380 86800
rect 11449 85794 11483 86800
rect 11547 85794 11581 86800
rect 11651 85794 11685 86800
rect 11759 85786 11793 86800
rect 11859 85794 11893 86800
rect 11967 85794 12001 86800
rect 12079 85794 12113 86800
rect 19866 85716 19974 86800
rect 21947 85794 21981 86800
rect 22050 85788 22084 86800
rect 22148 85794 22182 86800
rect 22252 85788 22286 86800
rect 22360 85794 22394 86800
rect 22460 85794 22494 86800
rect 22568 85786 22602 86800
rect 22680 85794 22714 86800
rect 30467 85720 30575 86800
rect 32548 85794 32582 86800
rect 32651 85794 32685 86800
rect 32749 85794 32783 86800
rect 32853 85794 32887 86800
rect 32961 85794 32995 86800
rect 33061 85782 33095 86800
rect 33169 85794 33203 86800
rect 33281 85794 33315 86800
rect 41068 85720 41176 86800
rect 2561 77978 2897 78033
rect 2561 77723 2616 77978
rect -6 146 134 152
rect -800 0 -6 140
rect -6 -12 134 -6
<< metal3 >>
rect 0 85389 42404 85489
rect 0 81638 42404 81738
rect 0 80894 42404 80994
rect 0 80127 42404 80227
rect 0 79395 42404 79495
rect 0 78454 42404 78594
rect 0 77764 42404 77904
rect 0 77226 42404 77366
rect 0 76536 42404 76676
rect 0 75998 42404 76138
rect 0 75308 42404 75448
rect 0 74770 42404 74910
rect 0 74080 42404 74220
rect 0 73542 42404 73682
rect 0 72852 42404 72992
rect 0 72314 42404 72454
rect 0 71624 42404 71764
rect 0 71086 42404 71226
rect 0 70396 42404 70536
rect 0 69858 42404 69998
rect 0 69168 42404 69308
rect 0 68630 42404 68770
rect 0 67940 42404 68080
rect 0 67402 42404 67542
rect 0 66712 42404 66852
rect 0 66174 42404 66314
rect 0 65484 42404 65624
rect 0 64946 42404 65086
rect 0 64256 42404 64396
rect 0 63718 42404 63858
rect 0 63028 42404 63168
rect 0 62490 42404 62630
rect 0 61800 42404 61940
rect 0 61262 42404 61402
rect 0 60572 42404 60712
rect 0 60034 42404 60174
rect 0 59344 42404 59484
rect 0 58806 42404 58946
rect 0 58116 42404 58256
rect 0 57578 42404 57718
rect 0 56888 42404 57028
rect 0 56350 42404 56490
rect 0 55660 42404 55800
rect 0 55122 42404 55262
rect 0 54432 42404 54572
rect 0 53894 42404 54034
rect 0 53204 42404 53344
rect 0 52666 42404 52806
rect 0 51976 42404 52116
rect 0 51438 42404 51578
rect 0 50748 42404 50888
rect 0 50210 42404 50350
rect 0 49520 42404 49660
rect 0 48982 42404 49122
rect 0 48292 42404 48432
rect 0 47754 42404 47894
rect 0 47064 42404 47204
rect 0 46526 42404 46666
rect 0 45836 42404 45976
rect 0 45298 42404 45438
rect 0 44608 42404 44748
rect 0 44070 42404 44210
rect 0 43380 42404 43520
rect 0 42842 42404 42982
rect 0 42152 42404 42292
rect 0 41614 42404 41754
rect 0 40924 42404 41064
rect 0 40386 42404 40526
rect 0 39696 42404 39836
rect 0 39158 42404 39298
rect 0 38468 42404 38608
rect 0 37930 42404 38070
rect 0 37240 42404 37380
rect 0 36702 42404 36842
rect 0 36012 42404 36152
rect 0 35474 42404 35614
rect 0 34784 42404 34924
rect 0 34246 42404 34386
rect 0 33556 42404 33696
rect 0 33018 42404 33158
rect 0 32328 42404 32468
rect 0 31790 42404 31930
rect 0 31100 42404 31240
rect 0 30562 42404 30702
rect 0 29872 42404 30012
rect 0 29334 42404 29474
rect 0 28644 42404 28784
rect 0 28106 42404 28246
rect 0 27416 42404 27556
rect 0 26878 42404 27018
rect 0 26188 42404 26328
rect 0 25650 42404 25790
rect 0 24960 42404 25100
rect 0 24422 42404 24562
rect 0 23732 42404 23872
rect 0 23194 42404 23334
rect 0 22504 42404 22644
rect 0 21966 42404 22106
rect 0 21276 42404 21416
rect 0 20738 42404 20878
rect 0 20048 42404 20188
rect 0 19510 42404 19650
rect 0 18820 42404 18960
rect 0 18282 42404 18422
rect 0 17592 42404 17732
rect 0 17054 42404 17194
rect 0 16364 42404 16504
rect 0 15826 42404 15966
rect 0 15136 42404 15276
rect 0 14598 42404 14738
rect 0 13908 42404 14048
rect 0 13370 42404 13510
rect 0 12680 42404 12820
rect 0 12142 42404 12282
rect 0 11452 42404 11592
rect 0 10914 42404 11054
rect 0 10224 42404 10364
rect 0 9686 42404 9826
rect 0 8996 42404 9136
rect 0 8458 42404 8598
rect 0 7768 42404 7908
rect 0 7230 42404 7370
rect 0 6540 42404 6680
rect 0 6002 42404 6142
rect 0 5312 42404 5452
rect 0 4774 42404 4914
rect 0 4084 42404 4224
rect 0 3546 42404 3686
rect 0 2856 42404 2996
rect 0 2318 42404 2458
rect 0 1628 42404 1768
rect 0 1090 42404 1230
rect 0 400 42404 540
use 4x8bit_tx_buffer  4x8bit_tx_buffer_0
timestamp 1686560844
transform 1 0 0 0 1 0
box 0 0 42404 85828
<< labels >>
rlabel metal2 9265 86000 9373 86800 1 VOUT0
port 38 n signal output
rlabel metal2 19866 86000 19974 86800 1 VOUT1
port 39 n signal output
rlabel metal2 30467 86000 30575 86800 1 VOUT2
port 40 n signal output
rlabel metal2 41068 86000 41176 86800 1 VOUT3
port 41 n signal output
rlabel metal2 -800 0 -200 140 7 VREFH
port 5 w signal input
flabel metal2 s 745 86000 779 86800 0 FreeSans 240 0 0 0 Din0[0]
port 6 nsew signal input
flabel metal2 s 848 86000 882 86800 0 FreeSans 240 0 0 0 Din0[1]
port 7 nsew signal input
flabel metal2 s 946 86000 980 86800 0 FreeSans 240 0 0 0 Din0[2]
port 8 nsew signal input
flabel metal2 s 1050 86000 1084 86800 0 FreeSans 240 0 0 0 Din0[3]
port 9 nsew signal input
flabel metal2 s 1158 86000 1192 86800 0 FreeSans 240 0 0 0 Din0[4]
port 10 nsew signal input
flabel metal2 s 1258 86000 1292 86800 0 FreeSans 240 0 0 0 Din0[5]
port 11 nsew signal input
flabel metal2 s 1366 86000 1400 86800 0 FreeSans 240 0 0 0 Din0[6]
port 12 nsew signal input
flabel metal2 s 1478 86000 1512 86800 0 FreeSans 240 0 0 0 Din0[7]
port 13 nsew signal input
flabel metal2 s 11346 86000 11380 86800 0 FreeSans 240 0 0 0 Din1[0]
port 14 nsew signal input
flabel metal2 s 11449 86000 11483 86800 0 FreeSans 240 0 0 0 Din1[1]
port 15 nsew signal input
flabel metal2 s 11547 86000 11581 86800 0 FreeSans 240 0 0 0 Din1[2]
port 16 nsew signal input
flabel metal2 s 11651 86000 11685 86800 0 FreeSans 240 0 0 0 Din1[3]
port 17 nsew signal input
flabel metal2 s 11759 86000 11793 86800 0 FreeSans 240 0 0 0 Din1[4]
port 18 nsew signal input
flabel metal2 s 11859 86000 11893 86800 0 FreeSans 240 0 0 0 Din1[5]
port 19 nsew signal input
flabel metal2 s 11967 86000 12001 86800 0 FreeSans 240 0 0 0 Din1[6]
port 20 nsew signal input
flabel metal2 s 12079 86000 12113 86800 0 FreeSans 240 0 0 0 Din1[7]
port 21 nsew signal input
flabel metal2 s 21947 86000 21981 86800 0 FreeSans 240 0 0 0 Din2[0]
port 22 nsew signal input
flabel metal2 s 22050 86000 22084 86800 0 FreeSans 240 0 0 0 Din2[1]
port 23 nsew signal input
flabel metal2 s 22148 86000 22182 86800 0 FreeSans 240 0 0 0 Din2[2]
port 24 nsew signal input
flabel metal2 s 22252 86000 22286 86800 0 FreeSans 240 0 0 0 Din2[3]
port 25 nsew signal input
flabel metal2 s 22360 86000 22394 86800 0 FreeSans 240 0 0 0 Din2[4]
port 26 nsew signal input
flabel metal2 s 22460 86000 22494 86800 0 FreeSans 240 0 0 0 Din2[5]
port 27 nsew signal input
flabel metal2 s 22568 86000 22602 86800 0 FreeSans 240 0 0 0 Din2[6]
port 28 nsew signal input
flabel metal2 s 22680 86000 22714 86800 0 FreeSans 240 0 0 0 Din2[7]
port 29 nsew signal input
flabel metal2 s 32548 86000 32582 86800 0 FreeSans 240 0 0 0 Din3[0]
port 30 nsew signal input
flabel metal2 s 32651 86000 32685 86800 0 FreeSans 240 0 0 0 Din3[1]
port 31 nsew signal input
flabel metal2 s 32749 86000 32783 86800 0 FreeSans 240 0 0 0 Din3[2]
port 32 nsew signal input
flabel metal2 s 32853 86000 32887 86800 0 FreeSans 240 0 0 0 Din3[3]
port 33 nsew signal input
flabel metal2 s 32961 86000 32995 86800 0 FreeSans 240 0 0 0 Din3[4]
port 34 nsew signal input
flabel metal2 s 33061 86000 33095 86800 0 FreeSans 240 0 0 0 Din3[5]
port 35 nsew signal input
flabel metal2 s 33169 86000 33203 86800 0 FreeSans 240 0 0 0 Din3[6]
port 36 nsew signal input
flabel metal2 s 33281 86000 33315 86800 0 FreeSans 240 0 0 0 Din3[7]
port 37 nsew signal input
rlabel metal3 0 400 42404 540 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 1628 42404 1768 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 2856 42404 2996 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 4084 42404 4224 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 5312 42404 5452 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 6540 42404 6680 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 7768 42404 7908 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 8996 42404 9136 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 10224 42404 10364 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 11452 42404 11592 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 12680 42404 12820 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 13908 42404 14048 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 15136 42404 15276 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 16364 42404 16504 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 17592 42404 17732 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 18820 42404 18960 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 20048 42404 20188 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 21276 42404 21416 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 22504 42404 22644 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 23732 42404 23872 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 24960 42404 25100 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 26188 42404 26328 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 27416 42404 27556 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 28644 42404 28784 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 29872 42404 30012 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 31100 42404 31240 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 32328 42404 32468 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 33556 42404 33696 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 34784 42404 34924 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 36012 42404 36152 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 37240 42404 37380 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 38468 42404 38608 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 39696 42404 39836 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 40924 42404 41064 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 42152 42404 42292 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 43380 42404 43520 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 44608 42404 44748 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 45836 42404 45976 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 47064 42404 47204 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 48292 42404 48432 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 49520 42404 49660 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 50748 42404 50888 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 51976 42404 52116 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 53204 42404 53344 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 54432 42404 54572 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 55660 42404 55800 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 56888 42404 57028 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 58116 42404 58256 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 59344 42404 59484 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 60572 42404 60712 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 61800 42404 61940 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 63028 42404 63168 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 64256 42404 64396 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 65484 42404 65624 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 66712 42404 66852 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 67940 42404 68080 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 69168 42404 69308 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 70396 42404 70536 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 71624 42404 71764 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 72852 42404 72992 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 74080 42404 74220 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 75308 42404 75448 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 76536 42404 76676 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 77764 42404 77904 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 1090 42404 1230 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 2318 42404 2458 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 3546 42404 3686 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 4774 42404 4914 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 6002 42404 6142 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 7230 42404 7370 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 8458 42404 8598 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 9686 42404 9826 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 10914 42404 11054 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 12142 42404 12282 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 13370 42404 13510 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 14598 42404 14738 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 15826 42404 15966 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 17054 42404 17194 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 18282 42404 18422 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 19510 42404 19650 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 20738 42404 20878 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 21966 42404 22106 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 23194 42404 23334 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 24422 42404 24562 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 25650 42404 25790 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 26878 42404 27018 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 28106 42404 28246 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 29334 42404 29474 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 30562 42404 30702 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 31790 42404 31930 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 33018 42404 33158 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 34246 42404 34386 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 35474 42404 35614 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 36702 42404 36842 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 37930 42404 38070 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 39158 42404 39298 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 40386 42404 40526 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 41614 42404 41754 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 42842 42404 42982 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 44070 42404 44210 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 45298 42404 45438 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 46526 42404 46666 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 47754 42404 47894 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 48982 42404 49122 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 50210 42404 50350 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 51438 42404 51578 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 52666 42404 52806 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 53894 42404 54034 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 55122 42404 55262 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 56350 42404 56490 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 57578 42404 57718 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 58806 42404 58946 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 60034 42404 60174 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 61262 42404 61402 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 62490 42404 62630 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 63718 42404 63858 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 64946 42404 65086 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 66174 42404 66314 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 67402 42404 67542 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 68630 42404 68770 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 69858 42404 69998 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 71086 42404 71226 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 72314 42404 72454 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 73542 42404 73682 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 74770 42404 74910 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 75998 42404 76138 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 77226 42404 77366 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 78454 42404 78594 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 80127 42404 80227 1 VCCD
port 3 n power bidirectional
rlabel metal3 0 79395 42404 79495 1 VSSD
port 4 n ground bidirectional
rlabel metal3 0 80894 42404 80994 1 VDDA
port 1 n power bidirectional
rlabel metal3 0 81638 42404 81738 1 VSSA
port 2 n ground bidirectional
rlabel metal3 0 85389 42404 85489 1 VDDA
port 1 n power bidirectional
<< properties >>
string FIXED_BBOX -500 -500 43000 86390
<< end >>
