magic
tech sky130A
magscale 1 2
timestamp 1692504018
<< metal3 >>
rect -1092 772 -120 800
rect -1092 148 -204 772
rect -140 148 -120 772
rect -1092 120 -120 148
rect 120 772 1092 800
rect 120 148 1008 772
rect 1072 148 1092 772
rect 120 120 1092 148
rect -1092 -148 -120 -120
rect -1092 -772 -204 -148
rect -140 -772 -120 -148
rect -1092 -800 -120 -772
rect 120 -148 1092 -120
rect 120 -772 1008 -148
rect 1072 -772 1092 -148
rect 120 -800 1092 -772
<< via3 >>
rect -204 148 -140 772
rect 1008 148 1072 772
rect -204 -772 -140 -148
rect 1008 -772 1072 -148
<< mimcap >>
rect -1052 720 -452 760
rect -1052 200 -1012 720
rect -492 200 -452 720
rect -1052 160 -452 200
rect 160 720 760 760
rect 160 200 200 720
rect 720 200 760 720
rect 160 160 760 200
rect -1052 -200 -452 -160
rect -1052 -720 -1012 -200
rect -492 -720 -452 -200
rect -1052 -760 -452 -720
rect 160 -200 760 -160
rect 160 -720 200 -200
rect 720 -720 760 -200
rect 160 -760 760 -720
<< mimcapcontact >>
rect -1012 200 -492 720
rect 200 200 720 720
rect -1012 -720 -492 -200
rect 200 -720 720 -200
<< metal4 >>
rect -804 721 -700 920
rect -224 772 -120 920
rect -1013 720 -491 721
rect -1013 200 -1012 720
rect -492 200 -491 720
rect -1013 199 -491 200
rect -804 -199 -700 199
rect -224 148 -204 772
rect -140 148 -120 772
rect 408 721 512 920
rect 988 772 1092 920
rect 199 720 721 721
rect 199 200 200 720
rect 720 200 721 720
rect 199 199 721 200
rect -224 -148 -120 148
rect -1013 -200 -491 -199
rect -1013 -720 -1012 -200
rect -492 -720 -491 -200
rect -1013 -721 -491 -720
rect -804 -920 -700 -721
rect -224 -772 -204 -148
rect -140 -772 -120 -148
rect 408 -199 512 199
rect 988 148 1008 772
rect 1072 148 1092 772
rect 988 -148 1092 148
rect 199 -200 721 -199
rect 199 -720 200 -200
rect 720 -720 721 -200
rect 199 -721 721 -720
rect -224 -920 -120 -772
rect 408 -920 512 -721
rect 988 -772 1008 -148
rect 1072 -772 1092 -148
rect 988 -920 1092 -772
<< properties >>
string FIXED_BBOX 120 120 800 800
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 3.0 l 3.0 val 20.28 carea 2.00 cperi 0.19 nx 2 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
