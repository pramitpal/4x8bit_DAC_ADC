magic
tech sky130A
magscale 1 2
timestamp 1692509756
<< error_p >>
rect -174 -130 174 202
rect -144 -164 144 -130
<< nwell >>
rect -144 -164 144 198
<< mvpmos >>
rect -50 -64 50 136
<< mvpdiff >>
rect -108 124 -50 136
rect -108 -52 -96 124
rect -62 -52 -50 124
rect -108 -64 -50 -52
rect 50 124 108 136
rect 50 -52 62 124
rect 96 -52 108 124
rect 50 -64 108 -52
<< mvpdiffc >>
rect -96 -52 -62 124
rect 62 -52 96 124
<< poly >>
rect -50 136 50 162
rect -50 -111 50 -64
rect -50 -145 -34 -111
rect 34 -145 50 -111
rect -50 -161 50 -145
<< polycont >>
rect -34 -145 34 -111
<< locali >>
rect -96 124 -62 140
rect -96 -68 -62 -52
rect 62 124 96 140
rect 62 -68 96 -52
rect -50 -145 -34 -111
rect 34 -145 50 -111
<< viali >>
rect -96 -52 -62 124
rect 62 -52 96 124
rect -34 -145 34 -111
<< metal1 >>
rect -102 124 -56 136
rect -102 -52 -96 124
rect -62 -52 -56 124
rect -102 -64 -56 -52
rect 56 124 102 136
rect 56 -52 62 124
rect 96 -52 102 124
rect 56 -64 102 -52
rect -46 -111 46 -105
rect -46 -145 -34 -111
rect 34 -145 46 -111
rect -46 -151 46 -145
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
