magic
tech sky130A
magscale 1 2
timestamp 1686481404
<< locali >>
rect 0 78948 504 79088
rect 0 0 434 140
<< metal2 >>
rect 745 85723 779 85828
rect 848 85707 882 85828
rect 946 85711 980 85828
rect 1050 85719 1084 85828
rect 1158 85719 1192 85828
rect 1258 85719 1292 85828
rect 1366 85719 1400 85828
rect 1478 85711 1512 85828
rect 9265 85590 9373 85828
rect 11346 85681 11380 85828
rect 11449 85683 11483 85828
rect 11547 85675 11581 85828
rect 11651 85713 11685 85828
rect 11759 85709 11793 85828
rect 11859 85693 11893 85828
rect 11967 85703 12001 85828
rect 12079 85689 12113 85828
rect 19866 85572 19974 85828
<< metal3 >>
rect 0 85389 320 85489
rect 0 81638 366 81738
rect 0 80127 388 80227
rect 0 79395 344 79495
rect 0 78454 442 78594
rect 0 77764 464 77904
use 8_bit_dac_tx_buffer_v2  8_bit_dac_tx_buffer_v2_0
array 0 1 10601 0 0 85828
timestamp 1686479781
transform 1 0 2409 0 1 180
box -2409 -180 8192 85648
<< labels >>
rlabel metal3 90 85438 90 85438 3 VDDA
rlabel metal3 60 81698 60 81698 3 VSSA
rlabel metal3 84 80188 84 80188 3 VCCD
rlabel metal3 90 79450 90 79450 3 VSSD
rlabel metal3 84 78528 84 78528 3 VDDA
rlabel metal3 76 77838 76 77838 3 VSSA
rlabel locali 34 79024 34 79024 3 VREFL
rlabel locali 94 74 94 74 3 VREFH
rlabel metal2 760 85800 760 85800 3 D00
rlabel metal2 866 85808 866 85808 3 D01
rlabel metal2 964 85810 964 85810 3 D02
rlabel metal2 1062 85820 1062 85820 3 D03
rlabel metal2 1168 85820 1168 85820 3 D04
rlabel metal2 1272 85820 1272 85820 3 D05
rlabel metal2 1376 85820 1376 85820 3 D06
rlabel metal2 1492 85818 1492 85818 3 D07
rlabel metal2 9308 85784 9308 85784 3 VOUT0
rlabel metal2 11360 85800 11360 85800 3 D10
rlabel metal2 11470 85812 11470 85812 3 D11
rlabel metal2 11566 85812 11566 85812 3 D12
rlabel metal2 11662 85816 11662 85816 3 D13
rlabel metal2 11776 85822 11776 85822 3 D14
rlabel metal2 11868 85816 11868 85816 3 D15
rlabel metal2 11980 85818 11980 85818 3 D16
rlabel metal2 12092 85814 12092 85814 3 D17
rlabel metal2 19912 85786 19912 85786 3 VOUT1
<< end >>
