magic
tech sky130A
magscale 1 2
timestamp 1687027365
<< metal1 >>
rect 6512 3766 6564 3772
rect 6512 3708 6564 3714
rect 6523 3651 6553 3708
rect 6523 3621 7015 3651
rect 6837 3555 6843 3562
rect 6516 3516 6843 3555
rect 6837 3510 6843 3516
rect 6895 3510 6901 3562
rect 6985 3521 7015 3621
rect 5191 3025 5197 3077
rect 5249 3070 5255 3077
rect 5249 3031 5625 3070
rect 5249 3025 5255 3031
rect 5191 2571 5197 2623
rect 5249 2616 5255 2623
rect 5249 2577 5587 2616
rect 5249 2571 5255 2577
rect 6908 2524 6936 2636
rect 7107 2536 7159 2542
rect 6908 2496 7107 2524
rect 7107 2478 7159 2484
<< via1 >>
rect 6512 3714 6564 3766
rect 6843 3510 6895 3562
rect 5197 3025 5249 3077
rect 5197 2571 5249 2623
rect 7107 2484 7159 2536
<< metal2 >>
rect 274 4773 329 4912
rect 378 4775 433 4912
rect 3564 4828 3605 4912
rect 5122 4788 5163 4912
rect 5202 4794 5243 4912
rect 42 4374 110 4570
rect 144 3644 212 3856
rect 6523 3766 6553 3887
rect 6506 3714 6512 3766
rect 6564 3714 6570 3766
rect 42 2033 110 3618
rect 5122 3543 5164 3633
rect 5202 3531 5244 3649
rect 5282 3515 5324 3659
rect 5362 3527 5404 3645
rect 5442 3519 5484 3653
rect 5522 3545 5564 3651
rect 6843 3562 6895 3568
rect 6895 3517 7150 3556
rect 6843 3504 6895 3510
rect 5197 3077 5249 3083
rect 144 1318 212 2893
rect 5122 2862 5163 3041
rect 5197 3019 5249 3025
rect 5282 2868 5323 3021
rect 5362 2862 5403 3026
rect 5442 2871 5483 3029
rect 5522 2840 5563 3021
rect 5197 2623 5202 2629
rect 5243 2623 5249 2629
rect 5197 2565 5202 2571
rect 5243 2565 5249 2571
rect 7101 2484 7107 2536
rect 7159 2484 7165 2536
rect 5122 2329 5164 2447
rect 5202 2321 5244 2457
rect 5282 2305 5324 2453
rect 5362 2325 5404 2457
rect 5442 2321 5484 2457
rect 5522 2323 5564 2459
rect 7119 2290 7147 2484
rect 5122 1272 5163 1374
rect 5202 1272 5243 1374
rect 277 0 332 107
rect 378 0 433 97
rect 3564 0 3605 92
use 3_bit_dac  3_bit_dac_0
array 0 0 7147 0 1 2456
timestamp 1687027365
transform 1 0 118 0 1 0
box -120 0 7606 2456
use switch_n_3v3  switch_n_3v3_0
timestamp 1687027365
transform 1 0 12004 0 1 3360
box -6932 -990 -4922 236
<< labels >>
rlabel metal2 74 4472 74 4472 7 VCC
rlabel metal2 182 3754 182 3754 7 VSS
rlabel metal2 312 4878 312 4878 7 D0
rlabel metal2 420 4878 420 4878 7 VREFL
rlabel metal2 316 22 316 22 7 D0_BUF
rlabel metal2 416 16 416 16 3 VREFH
rlabel metal2 3592 4898 3592 4898 3 D1
rlabel metal2 3574 8 3574 8 3 D1_BUF
rlabel metal2 5150 4900 5150 4900 3 D2
rlabel metal2 5222 4898 5222 4898 3 D3
rlabel metal2 5140 1282 5140 1282 3 D2_BUF
rlabel metal2 5212 1290 5212 1290 3 D3_BUF
rlabel metal2 7142 3534 7142 3534 3 VOUT
<< end >>
