magic
tech sky130A
timestamp 1690460607
<< error_p >>
rect -87 -75 87 75
<< nwell >>
rect -72 -73 72 73
<< mvpmos >>
rect -25 -42 25 42
<< mvpdiff >>
rect -54 36 -25 42
rect -54 -36 -48 36
rect -31 -36 -25 36
rect -54 -42 -25 -36
rect 25 36 54 42
rect 25 -36 31 36
rect 48 -36 54 36
rect 25 -42 54 -36
<< mvpdiffc >>
rect -48 -36 -31 36
rect 31 -36 48 36
<< poly >>
rect -25 42 25 55
rect -25 -55 25 -42
<< locali >>
rect -48 36 -31 44
rect -48 -44 -31 -36
rect 31 36 48 44
rect 31 -44 48 -36
<< viali >>
rect -48 -36 -31 36
rect 31 -36 48 36
<< metal1 >>
rect -51 36 -28 42
rect -51 -36 -48 36
rect -31 -36 -28 36
rect -51 -42 -28 -36
rect 28 36 51 42
rect 28 -36 31 36
rect 48 -36 51 36
rect 28 -42 51 -36
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 0.84 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
