VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO dac_top
  CLASS BLOCK ;
  FOREIGN dac_top ;
  ORIGIN 2.500 2.500 ;
  SIZE 217.500 BY 434.450 ;
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.000 426.945 39.775 427.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 404.470 0.835 404.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 5.450 12.255 6.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 11.590 12.255 12.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 17.730 12.255 18.430 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 23.870 12.255 24.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 30.010 12.255 30.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 36.150 12.255 36.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 42.290 12.255 42.990 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 48.430 12.255 49.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 54.570 12.255 55.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 60.710 12.255 61.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 66.850 12.255 67.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 72.990 12.255 73.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 79.130 12.255 79.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 85.270 12.255 85.970 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 91.410 12.255 92.110 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 97.550 12.255 98.250 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 103.690 12.255 104.390 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 109.830 12.255 110.530 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 115.970 12.255 116.670 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 122.110 12.255 122.810 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 128.250 12.255 128.950 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 134.390 12.255 135.090 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 140.530 12.255 141.230 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 146.670 12.255 147.370 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 152.810 12.255 153.510 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 158.950 12.255 159.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 165.090 12.255 165.790 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 171.230 12.255 171.930 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 177.370 12.255 178.070 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 183.510 12.255 184.210 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 189.650 12.255 190.350 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 195.790 12.255 196.490 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 201.930 12.255 202.630 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 208.070 12.255 208.770 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 214.210 12.255 214.910 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 220.350 12.255 221.050 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 226.490 12.255 227.190 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 232.630 12.255 233.330 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 238.770 12.255 239.470 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 244.910 12.255 245.610 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 251.050 12.255 251.750 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 257.190 12.255 257.890 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 263.330 12.255 264.030 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 269.470 12.255 270.170 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 275.610 12.255 276.310 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 281.750 12.255 282.450 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 287.890 12.255 288.590 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 294.030 12.255 294.730 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 300.170 12.255 300.870 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 306.310 12.255 307.010 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 312.450 12.255 313.150 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 318.590 12.255 319.290 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 324.730 12.255 325.430 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 330.870 12.255 331.570 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 337.010 12.255 337.710 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 343.150 12.255 343.850 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 349.290 12.255 349.990 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 355.430 12.255 356.130 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 361.570 12.255 362.270 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 367.710 12.255 368.410 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 373.850 12.255 374.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 379.990 12.255 380.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 386.130 12.255 386.830 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 392.270 12.255 392.970 ;
    END
  END VDDA
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.190 22.800 408.690 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 2.000 12.765 2.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 8.140 12.765 8.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 14.280 12.765 14.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 20.420 12.765 21.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 26.560 12.765 27.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 32.700 12.765 33.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 38.840 12.765 39.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 44.980 12.765 45.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 51.120 12.765 51.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 57.260 12.765 57.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 63.400 12.765 64.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 69.540 12.765 70.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 75.680 12.765 76.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 81.820 12.765 82.520 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 87.960 12.765 88.660 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 94.100 12.765 94.800 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 100.240 12.765 100.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 106.380 12.765 107.080 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 112.520 12.765 113.220 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 118.660 12.765 119.360 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 124.800 12.765 125.500 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 130.940 12.765 131.640 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 137.080 12.765 137.780 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 143.220 12.765 143.920 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 149.360 12.765 150.060 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 155.500 12.765 156.200 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 161.640 12.765 162.340 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 167.780 12.765 168.480 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 173.920 12.765 174.620 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 180.060 12.765 180.760 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 186.200 12.765 186.900 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 192.340 12.765 193.040 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 198.480 12.765 199.180 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 204.620 12.765 205.320 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 210.760 12.765 211.460 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 216.900 12.765 217.600 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 223.040 12.765 223.740 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 229.180 12.765 229.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 12.765 236.020 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 241.460 12.765 242.160 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 247.600 12.765 248.300 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 253.740 12.765 254.440 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 259.880 12.765 260.580 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 266.020 12.765 266.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 272.160 12.765 272.860 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 278.300 12.765 279.000 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 284.440 12.765 285.140 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 290.580 12.765 291.280 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 296.720 12.765 297.420 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 302.860 12.765 303.560 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 309.000 12.765 309.700 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 315.140 12.765 315.840 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 321.280 12.765 321.980 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 327.420 12.765 328.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 333.560 12.765 334.260 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 339.700 12.765 340.400 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 345.840 12.765 346.540 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 351.980 12.765 352.680 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 358.120 12.765 358.820 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 364.260 12.765 364.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 370.400 12.765 371.100 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 376.540 12.765 377.240 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 382.680 12.765 383.380 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 388.820 12.765 389.520 ;
    END
  END VSSA
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT -4.000 400.635 -0.095 401.135 ;
    END
  END VCCD
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT -4.000 396.975 -0.415 397.475 ;
    END
  END VSSD
  PIN VREFL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -4.000 394.740 -0.715 395.440 ;
    END
  END VREFL
  PIN VREFH
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -4.000 0.000 -0.030 0.700 ;
    END
  END VREFH
  PIN Din0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.725 405.755 3.895 434.000 ;
    END
  END Din0[0]
  PIN Din0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.240 405.395 4.410 434.000 ;
    END
  END Din0[1]
  PIN Din0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.730 405.715 4.900 434.000 ;
    END
  END Din0[2]
  PIN Din0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.250 406.035 5.420 434.000 ;
    END
  END Din0[3]
  PIN Din0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.790 406.355 5.960 434.000 ;
    END
  END Din0[4]
  PIN Din0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.290 406.675 6.460 434.000 ;
    END
  END Din0[5]
  PIN Din0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.830 406.995 7.000 434.000 ;
    END
  END Din0[6]
  PIN Din0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.390 407.315 7.560 434.000 ;
    END
  END Din0[7]
  PIN Din1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.730 405.755 56.900 434.000 ;
    END
  END Din1[0]
  PIN Din1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.245 405.395 57.415 434.000 ;
    END
  END Din1[1]
  PIN Din1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.735 405.715 57.905 434.000 ;
    END
  END Din1[2]
  PIN Din1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.255 406.035 58.425 434.000 ;
    END
  END Din1[3]
  PIN Din1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.795 406.355 58.965 434.000 ;
    END
  END Din1[4]
  PIN Din1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.295 406.675 59.465 434.000 ;
    END
  END Din1[5]
  PIN Din1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.835 406.995 60.005 434.000 ;
    END
  END Din1[6]
  PIN Din1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.395 407.315 60.565 434.000 ;
    END
  END Din1[7]
  PIN Din2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.735 405.755 109.905 434.000 ;
    END
  END Din2[0]
  PIN Din2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.250 405.395 110.420 434.000 ;
    END
  END Din2[1]
  PIN Din2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.740 405.715 110.910 434.000 ;
    END
  END Din2[2]
  PIN Din2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.260 406.035 111.430 434.000 ;
    END
  END Din2[3]
  PIN Din2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.800 406.355 111.970 434.000 ;
    END
  END Din2[4]
  PIN Din2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.300 406.675 112.470 434.000 ;
    END
  END Din2[5]
  PIN Din2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.840 406.995 113.010 434.000 ;
    END
  END Din2[6]
  PIN Din2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.400 407.315 113.570 434.000 ;
    END
  END Din2[7]
  PIN Din3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.740 405.755 162.910 434.000 ;
    END
  END Din3[0]
  PIN Din3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.255 405.395 163.425 434.000 ;
    END
  END Din3[1]
  PIN Din3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.745 405.715 163.915 434.000 ;
    END
  END Din3[2]
  PIN Din3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.265 406.035 164.435 434.000 ;
    END
  END Din3[3]
  PIN Din3[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.805 406.355 164.975 434.000 ;
    END
  END Din3[4]
  PIN Din3[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.305 406.675 165.475 434.000 ;
    END
  END Din3[5]
  PIN Din3[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.845 406.995 166.015 434.000 ;
    END
  END Din3[6]
  PIN Din3[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.405 407.315 166.575 434.000 ;
    END
  END Din3[7]
  PIN VOUT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.325 423.830 46.865 434.000 ;
    END
  END VOUT0
  PIN VOUT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.330 423.830 99.870 434.000 ;
    END
  END VOUT1
  PIN VOUT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.335 423.830 152.875 434.000 ;
    END
  END VOUT2
  PIN VOUT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.340 423.830 205.880 434.000 ;
    END
  END VOUT3
  OBS
      LAYER li1 ;
        RECT -0.685 0.000 212.020 427.735 ;
      LAYER met1 ;
        RECT -0.765 -0.060 207.290 427.745 ;
      LAYER met2 ;
        RECT -0.765 405.475 3.445 427.720 ;
        RECT 7.840 423.550 46.045 427.720 ;
        RECT 47.145 423.550 56.450 427.720 ;
        RECT 7.840 407.035 56.450 423.550 ;
        RECT 60.845 423.550 99.050 427.720 ;
        RECT 100.150 423.550 109.455 427.720 ;
        RECT 60.845 407.035 109.455 423.550 ;
        RECT 113.850 423.550 152.055 427.720 ;
        RECT 153.155 423.550 162.460 427.720 ;
        RECT 113.850 407.035 162.460 423.550 ;
        RECT 166.855 423.550 205.060 427.720 ;
        RECT 206.160 423.550 211.310 427.720 ;
        RECT 166.855 407.035 211.310 423.550 ;
        RECT 7.280 406.715 56.450 407.035 ;
        RECT 60.285 406.715 109.455 407.035 ;
        RECT 113.290 406.715 162.460 407.035 ;
        RECT 166.295 406.715 211.310 407.035 ;
        RECT 6.740 406.395 56.450 406.715 ;
        RECT 59.745 406.395 109.455 406.715 ;
        RECT 112.750 406.395 162.460 406.715 ;
        RECT 165.755 406.395 211.310 406.715 ;
        RECT 6.240 406.075 56.450 406.395 ;
        RECT 59.245 406.075 109.455 406.395 ;
        RECT 112.250 406.075 162.460 406.395 ;
        RECT 165.255 406.075 211.310 406.395 ;
        RECT 5.700 405.755 56.450 406.075 ;
        RECT 58.705 405.755 109.455 406.075 ;
        RECT 111.710 405.755 162.460 406.075 ;
        RECT 164.715 405.755 211.310 406.075 ;
        RECT 5.180 405.475 56.450 405.755 ;
        RECT 58.185 405.475 109.455 405.755 ;
        RECT 111.190 405.475 162.460 405.755 ;
        RECT -0.765 405.115 3.960 405.475 ;
        RECT 5.180 405.435 56.965 405.475 ;
        RECT 58.185 405.435 109.970 405.475 ;
        RECT 111.190 405.435 162.975 405.475 ;
        RECT 164.195 405.435 211.310 405.755 ;
        RECT 4.690 405.115 56.965 405.435 ;
        RECT 57.695 405.115 109.970 405.435 ;
        RECT 110.700 405.115 162.975 405.435 ;
        RECT 163.705 405.115 211.310 405.435 ;
        RECT -0.765 401.415 211.310 405.115 ;
        RECT 0.185 400.355 211.310 401.415 ;
        RECT -0.765 397.755 211.310 400.355 ;
        RECT -0.135 396.695 211.310 397.755 ;
        RECT -0.765 395.720 211.310 396.695 ;
        RECT -0.435 394.460 211.310 395.720 ;
        RECT -0.765 0.980 211.310 394.460 ;
        RECT 0.250 -0.060 211.310 0.980 ;
      LAYER met3 ;
        RECT -0.440 426.545 -0.400 427.640 ;
        RECT 40.175 426.545 212.020 427.640 ;
        RECT -0.440 409.090 212.020 426.545 ;
        RECT -0.440 407.790 -0.400 409.090 ;
        RECT 23.200 407.790 212.020 409.090 ;
        RECT -0.440 405.370 212.020 407.790 ;
        RECT -0.440 404.070 -0.400 405.370 ;
        RECT 1.235 404.070 212.020 405.370 ;
        RECT -0.440 393.370 212.020 404.070 ;
        RECT -0.440 391.870 -0.400 393.370 ;
        RECT 12.655 391.870 212.020 393.370 ;
        RECT -0.440 389.920 212.020 391.870 ;
        RECT -0.440 388.420 -0.400 389.920 ;
        RECT 13.165 388.420 212.020 389.920 ;
        RECT -0.440 387.230 212.020 388.420 ;
        RECT -0.440 385.730 -0.400 387.230 ;
        RECT 12.655 385.730 212.020 387.230 ;
        RECT -0.440 383.780 212.020 385.730 ;
        RECT -0.440 382.280 -0.400 383.780 ;
        RECT 13.165 382.280 212.020 383.780 ;
        RECT -0.440 381.090 212.020 382.280 ;
        RECT -0.440 379.590 -0.400 381.090 ;
        RECT 12.655 379.590 212.020 381.090 ;
        RECT -0.440 377.640 212.020 379.590 ;
        RECT -0.440 376.140 -0.400 377.640 ;
        RECT 13.165 376.140 212.020 377.640 ;
        RECT -0.440 374.950 212.020 376.140 ;
        RECT -0.440 373.450 -0.400 374.950 ;
        RECT 12.655 373.450 212.020 374.950 ;
        RECT -0.440 371.500 212.020 373.450 ;
        RECT -0.440 370.000 -0.400 371.500 ;
        RECT 13.165 370.000 212.020 371.500 ;
        RECT -0.440 368.810 212.020 370.000 ;
        RECT -0.440 367.310 -0.400 368.810 ;
        RECT 12.655 367.310 212.020 368.810 ;
        RECT -0.440 365.360 212.020 367.310 ;
        RECT -0.440 363.860 -0.400 365.360 ;
        RECT 13.165 363.860 212.020 365.360 ;
        RECT -0.440 362.670 212.020 363.860 ;
        RECT -0.440 361.170 -0.400 362.670 ;
        RECT 12.655 361.170 212.020 362.670 ;
        RECT -0.440 359.220 212.020 361.170 ;
        RECT -0.440 357.720 -0.400 359.220 ;
        RECT 13.165 357.720 212.020 359.220 ;
        RECT -0.440 356.530 212.020 357.720 ;
        RECT -0.440 355.030 -0.400 356.530 ;
        RECT 12.655 355.030 212.020 356.530 ;
        RECT -0.440 353.080 212.020 355.030 ;
        RECT -0.440 351.580 -0.400 353.080 ;
        RECT 13.165 351.580 212.020 353.080 ;
        RECT -0.440 350.390 212.020 351.580 ;
        RECT -0.440 348.890 -0.400 350.390 ;
        RECT 12.655 348.890 212.020 350.390 ;
        RECT -0.440 346.940 212.020 348.890 ;
        RECT -0.440 345.440 -0.400 346.940 ;
        RECT 13.165 345.440 212.020 346.940 ;
        RECT -0.440 344.250 212.020 345.440 ;
        RECT -0.440 342.750 -0.400 344.250 ;
        RECT 12.655 342.750 212.020 344.250 ;
        RECT -0.440 340.800 212.020 342.750 ;
        RECT -0.440 339.300 -0.400 340.800 ;
        RECT 13.165 339.300 212.020 340.800 ;
        RECT -0.440 338.110 212.020 339.300 ;
        RECT -0.440 336.610 -0.400 338.110 ;
        RECT 12.655 336.610 212.020 338.110 ;
        RECT -0.440 334.660 212.020 336.610 ;
        RECT -0.440 333.160 -0.400 334.660 ;
        RECT 13.165 333.160 212.020 334.660 ;
        RECT -0.440 331.970 212.020 333.160 ;
        RECT -0.440 330.470 -0.400 331.970 ;
        RECT 12.655 330.470 212.020 331.970 ;
        RECT -0.440 328.520 212.020 330.470 ;
        RECT -0.440 327.020 -0.400 328.520 ;
        RECT 13.165 327.020 212.020 328.520 ;
        RECT -0.440 325.830 212.020 327.020 ;
        RECT -0.440 324.330 -0.400 325.830 ;
        RECT 12.655 324.330 212.020 325.830 ;
        RECT -0.440 322.380 212.020 324.330 ;
        RECT -0.440 320.880 -0.400 322.380 ;
        RECT 13.165 320.880 212.020 322.380 ;
        RECT -0.440 319.690 212.020 320.880 ;
        RECT -0.440 318.190 -0.400 319.690 ;
        RECT 12.655 318.190 212.020 319.690 ;
        RECT -0.440 316.240 212.020 318.190 ;
        RECT -0.440 314.740 -0.400 316.240 ;
        RECT 13.165 314.740 212.020 316.240 ;
        RECT -0.440 313.550 212.020 314.740 ;
        RECT -0.440 312.050 -0.400 313.550 ;
        RECT 12.655 312.050 212.020 313.550 ;
        RECT -0.440 310.100 212.020 312.050 ;
        RECT -0.440 308.600 -0.400 310.100 ;
        RECT 13.165 308.600 212.020 310.100 ;
        RECT -0.440 307.410 212.020 308.600 ;
        RECT -0.440 305.910 -0.400 307.410 ;
        RECT 12.655 305.910 212.020 307.410 ;
        RECT -0.440 303.960 212.020 305.910 ;
        RECT -0.440 302.460 -0.400 303.960 ;
        RECT 13.165 302.460 212.020 303.960 ;
        RECT -0.440 301.270 212.020 302.460 ;
        RECT -0.440 299.770 -0.400 301.270 ;
        RECT 12.655 299.770 212.020 301.270 ;
        RECT -0.440 297.820 212.020 299.770 ;
        RECT -0.440 296.320 -0.400 297.820 ;
        RECT 13.165 296.320 212.020 297.820 ;
        RECT -0.440 295.130 212.020 296.320 ;
        RECT -0.440 293.630 -0.400 295.130 ;
        RECT 12.655 293.630 212.020 295.130 ;
        RECT -0.440 291.680 212.020 293.630 ;
        RECT -0.440 290.180 -0.400 291.680 ;
        RECT 13.165 290.180 212.020 291.680 ;
        RECT -0.440 288.990 212.020 290.180 ;
        RECT -0.440 287.490 -0.400 288.990 ;
        RECT 12.655 287.490 212.020 288.990 ;
        RECT -0.440 285.540 212.020 287.490 ;
        RECT -0.440 284.040 -0.400 285.540 ;
        RECT 13.165 284.040 212.020 285.540 ;
        RECT -0.440 282.850 212.020 284.040 ;
        RECT -0.440 281.350 -0.400 282.850 ;
        RECT 12.655 281.350 212.020 282.850 ;
        RECT -0.440 279.400 212.020 281.350 ;
        RECT -0.440 277.900 -0.400 279.400 ;
        RECT 13.165 277.900 212.020 279.400 ;
        RECT -0.440 276.710 212.020 277.900 ;
        RECT -0.440 275.210 -0.400 276.710 ;
        RECT 12.655 275.210 212.020 276.710 ;
        RECT -0.440 273.260 212.020 275.210 ;
        RECT -0.440 271.760 -0.400 273.260 ;
        RECT 13.165 271.760 212.020 273.260 ;
        RECT -0.440 270.570 212.020 271.760 ;
        RECT -0.440 269.070 -0.400 270.570 ;
        RECT 12.655 269.070 212.020 270.570 ;
        RECT -0.440 267.120 212.020 269.070 ;
        RECT -0.440 265.620 -0.400 267.120 ;
        RECT 13.165 265.620 212.020 267.120 ;
        RECT -0.440 264.430 212.020 265.620 ;
        RECT -0.440 262.930 -0.400 264.430 ;
        RECT 12.655 262.930 212.020 264.430 ;
        RECT -0.440 260.980 212.020 262.930 ;
        RECT -0.440 259.480 -0.400 260.980 ;
        RECT 13.165 259.480 212.020 260.980 ;
        RECT -0.440 258.290 212.020 259.480 ;
        RECT -0.440 256.790 -0.400 258.290 ;
        RECT 12.655 256.790 212.020 258.290 ;
        RECT -0.440 254.840 212.020 256.790 ;
        RECT -0.440 253.340 -0.400 254.840 ;
        RECT 13.165 253.340 212.020 254.840 ;
        RECT -0.440 252.150 212.020 253.340 ;
        RECT -0.440 250.650 -0.400 252.150 ;
        RECT 12.655 250.650 212.020 252.150 ;
        RECT -0.440 248.700 212.020 250.650 ;
        RECT -0.440 247.200 -0.400 248.700 ;
        RECT 13.165 247.200 212.020 248.700 ;
        RECT -0.440 246.010 212.020 247.200 ;
        RECT -0.440 244.510 -0.400 246.010 ;
        RECT 12.655 244.510 212.020 246.010 ;
        RECT -0.440 242.560 212.020 244.510 ;
        RECT -0.440 241.060 -0.400 242.560 ;
        RECT 13.165 241.060 212.020 242.560 ;
        RECT -0.440 239.870 212.020 241.060 ;
        RECT -0.440 238.370 -0.400 239.870 ;
        RECT 12.655 238.370 212.020 239.870 ;
        RECT -0.440 236.420 212.020 238.370 ;
        RECT -0.440 234.920 -0.400 236.420 ;
        RECT 13.165 234.920 212.020 236.420 ;
        RECT -0.440 233.730 212.020 234.920 ;
        RECT -0.440 232.230 -0.400 233.730 ;
        RECT 12.655 232.230 212.020 233.730 ;
        RECT -0.440 230.280 212.020 232.230 ;
        RECT -0.440 228.780 -0.400 230.280 ;
        RECT 13.165 228.780 212.020 230.280 ;
        RECT -0.440 227.590 212.020 228.780 ;
        RECT -0.440 226.090 -0.400 227.590 ;
        RECT 12.655 226.090 212.020 227.590 ;
        RECT -0.440 224.140 212.020 226.090 ;
        RECT -0.440 222.640 -0.400 224.140 ;
        RECT 13.165 222.640 212.020 224.140 ;
        RECT -0.440 221.450 212.020 222.640 ;
        RECT -0.440 219.950 -0.400 221.450 ;
        RECT 12.655 219.950 212.020 221.450 ;
        RECT -0.440 218.000 212.020 219.950 ;
        RECT -0.440 216.500 -0.400 218.000 ;
        RECT 13.165 216.500 212.020 218.000 ;
        RECT -0.440 215.310 212.020 216.500 ;
        RECT -0.440 213.810 -0.400 215.310 ;
        RECT 12.655 213.810 212.020 215.310 ;
        RECT -0.440 211.860 212.020 213.810 ;
        RECT -0.440 210.360 -0.400 211.860 ;
        RECT 13.165 210.360 212.020 211.860 ;
        RECT -0.440 209.170 212.020 210.360 ;
        RECT -0.440 207.670 -0.400 209.170 ;
        RECT 12.655 207.670 212.020 209.170 ;
        RECT -0.440 205.720 212.020 207.670 ;
        RECT -0.440 204.220 -0.400 205.720 ;
        RECT 13.165 204.220 212.020 205.720 ;
        RECT -0.440 203.030 212.020 204.220 ;
        RECT -0.440 201.530 -0.400 203.030 ;
        RECT 12.655 201.530 212.020 203.030 ;
        RECT -0.440 199.580 212.020 201.530 ;
        RECT -0.440 198.080 -0.400 199.580 ;
        RECT 13.165 198.080 212.020 199.580 ;
        RECT -0.440 196.890 212.020 198.080 ;
        RECT -0.440 195.390 -0.400 196.890 ;
        RECT 12.655 195.390 212.020 196.890 ;
        RECT -0.440 193.440 212.020 195.390 ;
        RECT -0.440 191.940 -0.400 193.440 ;
        RECT 13.165 191.940 212.020 193.440 ;
        RECT -0.440 190.750 212.020 191.940 ;
        RECT -0.440 189.250 -0.400 190.750 ;
        RECT 12.655 189.250 212.020 190.750 ;
        RECT -0.440 187.300 212.020 189.250 ;
        RECT -0.440 185.800 -0.400 187.300 ;
        RECT 13.165 185.800 212.020 187.300 ;
        RECT -0.440 184.610 212.020 185.800 ;
        RECT -0.440 183.110 -0.400 184.610 ;
        RECT 12.655 183.110 212.020 184.610 ;
        RECT -0.440 181.160 212.020 183.110 ;
        RECT -0.440 179.660 -0.400 181.160 ;
        RECT 13.165 179.660 212.020 181.160 ;
        RECT -0.440 178.470 212.020 179.660 ;
        RECT -0.440 176.970 -0.400 178.470 ;
        RECT 12.655 176.970 212.020 178.470 ;
        RECT -0.440 175.020 212.020 176.970 ;
        RECT -0.440 173.520 -0.400 175.020 ;
        RECT 13.165 173.520 212.020 175.020 ;
        RECT -0.440 172.330 212.020 173.520 ;
        RECT -0.440 170.830 -0.400 172.330 ;
        RECT 12.655 170.830 212.020 172.330 ;
        RECT -0.440 168.880 212.020 170.830 ;
        RECT -0.440 167.380 -0.400 168.880 ;
        RECT 13.165 167.380 212.020 168.880 ;
        RECT -0.440 166.190 212.020 167.380 ;
        RECT -0.440 164.690 -0.400 166.190 ;
        RECT 12.655 164.690 212.020 166.190 ;
        RECT -0.440 162.740 212.020 164.690 ;
        RECT -0.440 161.240 -0.400 162.740 ;
        RECT 13.165 161.240 212.020 162.740 ;
        RECT -0.440 160.050 212.020 161.240 ;
        RECT -0.440 158.550 -0.400 160.050 ;
        RECT 12.655 158.550 212.020 160.050 ;
        RECT -0.440 156.600 212.020 158.550 ;
        RECT -0.440 155.100 -0.400 156.600 ;
        RECT 13.165 155.100 212.020 156.600 ;
        RECT -0.440 153.910 212.020 155.100 ;
        RECT -0.440 152.410 -0.400 153.910 ;
        RECT 12.655 152.410 212.020 153.910 ;
        RECT -0.440 150.460 212.020 152.410 ;
        RECT -0.440 148.960 -0.400 150.460 ;
        RECT 13.165 148.960 212.020 150.460 ;
        RECT -0.440 147.770 212.020 148.960 ;
        RECT -0.440 146.270 -0.400 147.770 ;
        RECT 12.655 146.270 212.020 147.770 ;
        RECT -0.440 144.320 212.020 146.270 ;
        RECT -0.440 142.820 -0.400 144.320 ;
        RECT 13.165 142.820 212.020 144.320 ;
        RECT -0.440 141.630 212.020 142.820 ;
        RECT -0.440 140.130 -0.400 141.630 ;
        RECT 12.655 140.130 212.020 141.630 ;
        RECT -0.440 138.180 212.020 140.130 ;
        RECT -0.440 136.680 -0.400 138.180 ;
        RECT 13.165 136.680 212.020 138.180 ;
        RECT -0.440 135.490 212.020 136.680 ;
        RECT -0.440 133.990 -0.400 135.490 ;
        RECT 12.655 133.990 212.020 135.490 ;
        RECT -0.440 132.040 212.020 133.990 ;
        RECT -0.440 130.540 -0.400 132.040 ;
        RECT 13.165 130.540 212.020 132.040 ;
        RECT -0.440 129.350 212.020 130.540 ;
        RECT -0.440 127.850 -0.400 129.350 ;
        RECT 12.655 127.850 212.020 129.350 ;
        RECT -0.440 125.900 212.020 127.850 ;
        RECT -0.440 124.400 -0.400 125.900 ;
        RECT 13.165 124.400 212.020 125.900 ;
        RECT -0.440 123.210 212.020 124.400 ;
        RECT -0.440 121.710 -0.400 123.210 ;
        RECT 12.655 121.710 212.020 123.210 ;
        RECT -0.440 119.760 212.020 121.710 ;
        RECT -0.440 118.260 -0.400 119.760 ;
        RECT 13.165 118.260 212.020 119.760 ;
        RECT -0.440 117.070 212.020 118.260 ;
        RECT -0.440 115.570 -0.400 117.070 ;
        RECT 12.655 115.570 212.020 117.070 ;
        RECT -0.440 113.620 212.020 115.570 ;
        RECT -0.440 112.120 -0.400 113.620 ;
        RECT 13.165 112.120 212.020 113.620 ;
        RECT -0.440 110.930 212.020 112.120 ;
        RECT -0.440 109.430 -0.400 110.930 ;
        RECT 12.655 109.430 212.020 110.930 ;
        RECT -0.440 107.480 212.020 109.430 ;
        RECT -0.440 105.980 -0.400 107.480 ;
        RECT 13.165 105.980 212.020 107.480 ;
        RECT -0.440 104.790 212.020 105.980 ;
        RECT -0.440 103.290 -0.400 104.790 ;
        RECT 12.655 103.290 212.020 104.790 ;
        RECT -0.440 101.340 212.020 103.290 ;
        RECT -0.440 99.840 -0.400 101.340 ;
        RECT 13.165 99.840 212.020 101.340 ;
        RECT -0.440 98.650 212.020 99.840 ;
        RECT -0.440 97.150 -0.400 98.650 ;
        RECT 12.655 97.150 212.020 98.650 ;
        RECT -0.440 95.200 212.020 97.150 ;
        RECT -0.440 93.700 -0.400 95.200 ;
        RECT 13.165 93.700 212.020 95.200 ;
        RECT -0.440 92.510 212.020 93.700 ;
        RECT -0.440 91.010 -0.400 92.510 ;
        RECT 12.655 91.010 212.020 92.510 ;
        RECT -0.440 89.060 212.020 91.010 ;
        RECT -0.440 87.560 -0.400 89.060 ;
        RECT 13.165 87.560 212.020 89.060 ;
        RECT -0.440 86.370 212.020 87.560 ;
        RECT -0.440 84.870 -0.400 86.370 ;
        RECT 12.655 84.870 212.020 86.370 ;
        RECT -0.440 82.920 212.020 84.870 ;
        RECT -0.440 81.420 -0.400 82.920 ;
        RECT 13.165 81.420 212.020 82.920 ;
        RECT -0.440 80.230 212.020 81.420 ;
        RECT -0.440 78.730 -0.400 80.230 ;
        RECT 12.655 78.730 212.020 80.230 ;
        RECT -0.440 76.780 212.020 78.730 ;
        RECT -0.440 75.280 -0.400 76.780 ;
        RECT 13.165 75.280 212.020 76.780 ;
        RECT -0.440 74.090 212.020 75.280 ;
        RECT -0.440 72.590 -0.400 74.090 ;
        RECT 12.655 72.590 212.020 74.090 ;
        RECT -0.440 70.640 212.020 72.590 ;
        RECT -0.440 69.140 -0.400 70.640 ;
        RECT 13.165 69.140 212.020 70.640 ;
        RECT -0.440 67.950 212.020 69.140 ;
        RECT -0.440 66.450 -0.400 67.950 ;
        RECT 12.655 66.450 212.020 67.950 ;
        RECT -0.440 64.500 212.020 66.450 ;
        RECT -0.440 63.000 -0.400 64.500 ;
        RECT 13.165 63.000 212.020 64.500 ;
        RECT -0.440 61.810 212.020 63.000 ;
        RECT -0.440 60.310 -0.400 61.810 ;
        RECT 12.655 60.310 212.020 61.810 ;
        RECT -0.440 58.360 212.020 60.310 ;
        RECT -0.440 56.860 -0.400 58.360 ;
        RECT 13.165 56.860 212.020 58.360 ;
        RECT -0.440 55.670 212.020 56.860 ;
        RECT -0.440 54.170 -0.400 55.670 ;
        RECT 12.655 54.170 212.020 55.670 ;
        RECT -0.440 52.220 212.020 54.170 ;
        RECT -0.440 50.720 -0.400 52.220 ;
        RECT 13.165 50.720 212.020 52.220 ;
        RECT -0.440 49.530 212.020 50.720 ;
        RECT -0.440 48.030 -0.400 49.530 ;
        RECT 12.655 48.030 212.020 49.530 ;
        RECT -0.440 46.080 212.020 48.030 ;
        RECT -0.440 44.580 -0.400 46.080 ;
        RECT 13.165 44.580 212.020 46.080 ;
        RECT -0.440 43.390 212.020 44.580 ;
        RECT -0.440 41.890 -0.400 43.390 ;
        RECT 12.655 41.890 212.020 43.390 ;
        RECT -0.440 39.940 212.020 41.890 ;
        RECT -0.440 38.440 -0.400 39.940 ;
        RECT 13.165 38.440 212.020 39.940 ;
        RECT -0.440 37.250 212.020 38.440 ;
        RECT -0.440 35.750 -0.400 37.250 ;
        RECT 12.655 35.750 212.020 37.250 ;
        RECT -0.440 33.800 212.020 35.750 ;
        RECT -0.440 32.300 -0.400 33.800 ;
        RECT 13.165 32.300 212.020 33.800 ;
        RECT -0.440 31.110 212.020 32.300 ;
        RECT -0.440 29.610 -0.400 31.110 ;
        RECT 12.655 29.610 212.020 31.110 ;
        RECT -0.440 27.660 212.020 29.610 ;
        RECT -0.440 26.160 -0.400 27.660 ;
        RECT 13.165 26.160 212.020 27.660 ;
        RECT -0.440 24.970 212.020 26.160 ;
        RECT -0.440 23.470 -0.400 24.970 ;
        RECT 12.655 23.470 212.020 24.970 ;
        RECT -0.440 21.520 212.020 23.470 ;
        RECT -0.440 20.020 -0.400 21.520 ;
        RECT 13.165 20.020 212.020 21.520 ;
        RECT -0.440 18.830 212.020 20.020 ;
        RECT -0.440 17.330 -0.400 18.830 ;
        RECT 12.655 17.330 212.020 18.830 ;
        RECT -0.440 15.380 212.020 17.330 ;
        RECT -0.440 13.880 -0.400 15.380 ;
        RECT 13.165 13.880 212.020 15.380 ;
        RECT -0.440 12.690 212.020 13.880 ;
        RECT -0.440 11.190 -0.400 12.690 ;
        RECT 12.655 11.190 212.020 12.690 ;
        RECT -0.440 9.240 212.020 11.190 ;
        RECT -0.440 7.740 -0.400 9.240 ;
        RECT 13.165 7.740 212.020 9.240 ;
        RECT -0.440 6.550 212.020 7.740 ;
        RECT -0.440 5.050 -0.400 6.550 ;
        RECT 12.655 5.050 212.020 6.550 ;
        RECT -0.440 3.100 212.020 5.050 ;
        RECT -0.440 2.000 -0.400 3.100 ;
        RECT 13.165 2.000 212.020 3.100 ;
  END
END dac_top
END LIBRARY

