magic
tech sky130A
magscale 1 2
timestamp 1687027365
<< metal1 >>
rect 6968 20828 6974 20880
rect 7026 20828 7032 20880
rect 6838 20748 6844 20755
rect 6516 20709 6844 20748
rect 6838 20703 6844 20709
rect 6896 20703 6902 20755
rect 6985 20693 7015 20828
rect 5431 20218 5437 20270
rect 5489 20263 5495 20270
rect 5489 20224 5629 20263
rect 5489 20218 5495 20224
rect 7128 19823 7134 19835
rect 5429 19764 5435 19816
rect 5487 19809 5493 19816
rect 5487 19770 5572 19809
rect 6908 19795 7134 19823
rect 7128 19783 7134 19795
rect 7186 19783 7192 19835
rect 5487 19764 5493 19770
<< via1 >>
rect 6974 20828 7026 20880
rect 6844 20703 6896 20755
rect 5437 20218 5489 20270
rect 5435 19764 5487 19816
rect 7134 19783 7186 19835
<< metal2 >>
rect 274 39123 329 39296
rect 378 39147 433 39296
rect 3564 39184 3605 39296
rect 5122 39172 5163 39296
rect 5202 39160 5243 39296
rect 5282 39168 5323 39296
rect 5362 39174 5403 39296
rect 5442 39166 5483 39296
rect 7321 30411 7431 30450
rect 6974 20880 7026 20886
rect 42 19188 110 20768
rect 5122 20725 5164 20833
rect 5202 20733 5244 20832
rect 5282 20751 5324 20832
rect 5362 20757 5404 20832
rect 5442 20747 5484 20832
rect 5522 20745 5564 20832
rect 7392 20876 7431 30411
rect 7026 20837 7431 20876
rect 6974 20822 7026 20828
rect 6844 20755 6896 20761
rect 6896 20710 7470 20749
rect 6844 20697 6896 20703
rect 5437 20270 5489 20276
rect 144 18532 212 20118
rect 5122 20080 5163 20217
rect 5202 20028 5243 20222
rect 5282 20058 5323 20214
rect 5362 20034 5403 20237
rect 5437 20212 5489 20218
rect 5522 20068 5563 20214
rect 7134 19835 7186 19841
rect 5435 19816 5487 19822
rect 7186 19795 7427 19823
rect 7134 19777 7186 19783
rect 5435 19758 5487 19764
rect 5122 19513 5164 19655
rect 5202 19495 5244 19641
rect 5282 19489 5324 19637
rect 5362 19499 5404 19639
rect 5442 19509 5484 19651
rect 5522 19495 5564 19643
rect 7388 10802 7427 19795
rect 7321 10763 7427 10802
rect 5122 1141 5163 1274
rect 5202 1141 5243 1280
rect 5282 1141 5323 1278
rect 5362 1141 5403 1282
rect 5442 1141 5483 1286
rect 277 0 332 175
rect 378 0 433 193
rect 3564 0 3605 142
use 6_bit_dac  6_bit_dac_0
array 0 0 7360 0 1 19648
timestamp 1687027365
transform 1 0 0 0 1 0
box -2 0 7724 19648
use switch_n_3v3  switch_n_3v3_1
timestamp 1687027365
transform 1 0 12004 0 1 20553
box -6932 -990 -4922 236
<< labels >>
rlabel metal2 70 19650 70 19650 3 VCC
rlabel metal2 178 19646 178 19646 3 VSS
rlabel metal2 306 39236 306 39236 3 D0
rlabel metal2 390 39234 390 39234 3 VREFL
rlabel metal2 3572 39280 3572 39280 3 D1
rlabel metal2 5130 39288 5130 39288 3 D2
rlabel metal2 5212 39288 5212 39288 3 D3
rlabel metal2 5292 39286 5292 39286 3 D4
rlabel metal2 5374 39286 5374 39286 3 D5
rlabel metal2 5456 39280 5456 39280 3 D6
rlabel metal2 306 32 306 32 3 D0_BUF
rlabel metal2 396 40 396 40 3 VREFH
rlabel metal2 3580 30 3580 30 3 D1_BUF
rlabel metal2 5144 1164 5144 1164 3 D2_BUF
rlabel metal2 5210 1160 5210 1160 3 D3_BUF
rlabel metal2 5294 1156 5294 1156 3 D4_BUF
rlabel metal2 5370 1156 5370 1156 3 D5_BUF
rlabel metal2 5456 1154 5456 1154 3 D6_BUF
rlabel metal2 7434 20728 7434 20728 3 VOUT
<< end >>
