VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO dac_top
  CLASS BLOCK ;
  FOREIGN dac_top ;
  ORIGIN 5.000 5.000 ;
  SIZE 164.520 BY 436.055 ;
  PIN VDDA
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.615 154.520 425.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 401.915 154.520 402.415 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 5.155 154.520 5.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 11.295 154.520 11.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 17.435 154.520 18.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 23.575 154.520 24.275 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 29.715 154.520 30.415 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 35.855 154.520 36.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 41.995 154.520 42.695 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 48.135 154.520 48.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 54.275 154.520 54.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 60.415 154.520 61.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 66.555 154.520 67.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 72.695 154.520 73.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 78.835 154.520 79.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 84.975 154.520 85.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 91.115 154.520 91.815 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 97.255 154.520 97.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 103.395 154.520 104.095 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 109.535 154.520 110.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 115.675 154.520 116.375 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 121.815 154.520 122.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 127.955 154.520 128.655 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 134.095 154.520 134.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 140.235 154.520 140.935 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 146.375 154.520 147.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 152.515 154.520 153.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 158.655 154.520 159.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 164.795 154.520 165.495 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 170.935 154.520 171.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 177.075 154.520 177.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 183.215 154.520 183.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 189.355 154.520 190.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 195.495 154.520 196.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 201.635 154.520 202.335 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 207.775 154.520 208.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 213.915 154.520 214.615 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 220.055 154.520 220.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 226.195 154.520 226.895 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 232.335 154.520 233.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 238.475 154.520 239.175 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 244.615 154.520 245.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 250.755 154.520 251.455 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 256.895 154.520 257.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 263.035 154.520 263.735 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 269.175 154.520 269.875 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 275.315 154.520 276.015 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 281.455 154.520 282.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 287.595 154.520 288.295 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 293.735 154.520 294.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 299.875 154.520 300.575 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 306.015 154.520 306.715 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 312.155 154.520 312.855 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 318.295 154.520 318.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 324.435 154.520 325.135 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 330.575 154.520 331.275 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 336.715 154.520 337.415 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 342.855 154.520 343.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 348.995 154.520 349.695 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 355.135 154.520 355.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 361.275 154.520 361.975 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 367.415 154.520 368.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 373.555 154.520 374.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 379.695 154.520 380.395 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 385.835 154.520 386.535 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 391.975 154.520 392.675 ;
    END
  END VDDA
  PIN VSSA
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.000 407.565 154.520 409.065 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 1.705 154.520 2.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 7.845 154.520 8.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 13.985 154.520 14.685 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 20.125 154.520 20.825 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 26.265 154.520 26.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 32.405 154.520 33.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 38.545 154.520 39.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 44.685 154.520 45.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 50.825 154.520 51.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 56.965 154.520 57.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 63.105 154.520 63.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 69.245 154.520 69.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 75.385 154.520 76.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 81.525 154.520 82.225 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 87.665 154.520 88.365 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 93.805 154.520 94.505 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 99.945 154.520 100.645 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 106.085 154.520 106.785 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 112.225 154.520 112.925 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 118.365 154.520 119.065 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 124.505 154.520 125.205 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 130.645 154.520 131.345 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 136.785 154.520 137.485 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 142.925 154.520 143.625 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 149.065 154.520 149.765 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 155.205 154.520 155.905 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 161.345 154.520 162.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 167.485 154.520 168.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 173.625 154.520 174.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 179.765 154.520 180.465 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 185.905 154.520 186.605 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 192.045 154.520 192.745 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 198.185 154.520 198.885 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 204.325 154.520 205.025 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 210.465 154.520 211.165 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 216.605 154.520 217.305 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 222.745 154.520 223.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 228.885 154.520 229.585 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 235.025 154.520 235.725 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 241.165 154.520 241.865 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 247.305 154.520 248.005 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 253.445 154.520 254.145 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 259.585 154.520 260.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 265.725 154.520 266.425 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 271.865 154.520 272.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 278.005 154.520 278.705 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 284.145 154.520 284.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 290.285 154.520 290.985 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 296.425 154.520 297.125 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 302.565 154.520 303.265 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 308.705 154.520 309.405 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 314.845 154.520 315.545 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 320.985 154.520 321.685 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 327.125 154.520 327.825 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 333.265 154.520 333.965 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 339.405 154.520 340.105 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 345.545 154.520 346.245 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 351.685 154.520 352.385 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 357.825 154.520 358.525 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 363.965 154.520 364.665 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 370.105 154.520 370.805 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 376.245 154.520 376.945 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 382.385 154.520 383.085 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.000 388.525 154.520 389.225 ;
    END
  END VSSA
  PIN VCCD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.265 154.520 395.765 ;
    END
  END VCCD
  PIN VSSD
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.565 154.520 398.065 ;
    END
  END VSSD
  PIN VREFH
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -7.600 0.000 -1.500 0.500 ;
    END
  END VREFH
  PIN Din0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.210 403.645 3.410 434.300 ;
    END
  END Din0[0]
  PIN Din0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.900 404.095 4.100 434.300 ;
    END
  END Din0[1]
  PIN Din0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.580 404.545 4.780 434.300 ;
    END
  END Din0[2]
  PIN Din0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.250 404.995 5.450 434.300 ;
    END
  END Din0[3]
  PIN Din0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.910 405.455 6.110 434.300 ;
    END
  END Din0[4]
  PIN Din0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.570 405.955 6.770 434.300 ;
    END
  END Din0[5]
  PIN Din0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.230 406.445 7.430 434.300 ;
    END
  END Din0[6]
  PIN Din0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.900 406.985 8.100 434.300 ;
    END
  END Din0[7]
  PIN VOUT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.040 414.115 32.280 434.300 ;
    END
  END VOUT0
  PIN Din1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.840 403.645 42.040 434.300 ;
    END
  END Din1[0]
  PIN Din1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.530 404.095 42.730 434.300 ;
    END
  END Din1[1]
  PIN Din1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.210 404.545 43.410 434.300 ;
    END
  END Din1[2]
  PIN Din1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.880 404.995 44.080 434.300 ;
    END
  END Din1[3]
  PIN Din1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.540 405.455 44.740 434.300 ;
    END
  END Din1[4]
  PIN Din1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.200 405.955 45.400 434.300 ;
    END
  END Din1[5]
  PIN Din1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.860 406.445 46.060 434.300 ;
    END
  END Din1[6]
  PIN Din1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.530 406.985 46.730 434.300 ;
    END
  END Din1[7]
  PIN VOUT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.670 414.115 70.910 434.300 ;
    END
  END VOUT1
  PIN Din2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.470 403.645 80.670 434.300 ;
    END
  END Din2[0]
  PIN Din2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.160 404.095 81.360 434.300 ;
    END
  END Din2[1]
  PIN Din2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.840 404.545 82.040 434.300 ;
    END
  END Din2[2]
  PIN Din2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.510 404.995 82.710 434.300 ;
    END
  END Din2[3]
  PIN Din2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.170 405.455 83.370 434.300 ;
    END
  END Din2[4]
  PIN Din2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.830 405.955 84.030 434.300 ;
    END
  END Din2[5]
  PIN Din2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.490 406.445 84.690 434.300 ;
    END
  END Din2[6]
  PIN Din2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.160 406.985 85.360 434.300 ;
    END
  END Din2[7]
  PIN VOUT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.300 414.115 109.540 434.300 ;
    END
  END VOUT2
  PIN Din3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.100 403.645 119.300 434.300 ;
    END
  END Din3[0]
  PIN Din3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.790 404.095 119.990 434.300 ;
    END
  END Din3[1]
  PIN Din3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.470 404.545 120.670 434.300 ;
    END
  END Din3[2]
  PIN Din3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.140 404.995 121.340 434.300 ;
    END
  END Din3[3]
  PIN Din3[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.800 405.455 122.000 434.300 ;
    END
  END Din3[4]
  PIN Din3[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.460 405.955 122.660 434.300 ;
    END
  END Din3[5]
  PIN Din3[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.120 406.445 123.320 434.300 ;
    END
  END Din3[6]
  PIN Din3[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.790 406.985 123.990 434.300 ;
    END
  END Din3[7]
  PIN VOUT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.930 414.115 148.170 434.300 ;
    END
  END VOUT3
  OBS
      LAYER li1 ;
        RECT 2.710 1.210 150.200 425.115 ;
      LAYER met1 ;
        RECT -1.530 0.000 154.520 425.115 ;
      LAYER met2 ;
        RECT -1.500 403.365 2.930 425.115 ;
        RECT 8.380 413.835 31.760 425.115 ;
        RECT 32.560 413.835 41.560 425.115 ;
        RECT 8.380 406.705 41.560 413.835 ;
        RECT 47.010 413.835 70.390 425.115 ;
        RECT 71.190 413.835 80.190 425.115 ;
        RECT 47.010 406.705 80.190 413.835 ;
        RECT 85.640 413.835 109.020 425.115 ;
        RECT 109.820 413.835 118.820 425.115 ;
        RECT 85.640 406.705 118.820 413.835 ;
        RECT 124.270 413.835 147.650 425.115 ;
        RECT 148.450 413.835 154.180 425.115 ;
        RECT 124.270 406.705 154.180 413.835 ;
        RECT 7.710 406.165 41.560 406.705 ;
        RECT 46.340 406.165 80.190 406.705 ;
        RECT 84.970 406.165 118.820 406.705 ;
        RECT 123.600 406.165 154.180 406.705 ;
        RECT 7.050 405.675 41.560 406.165 ;
        RECT 45.680 405.675 80.190 406.165 ;
        RECT 84.310 405.675 118.820 406.165 ;
        RECT 122.940 405.675 154.180 406.165 ;
        RECT 6.390 405.175 41.560 405.675 ;
        RECT 45.020 405.175 80.190 405.675 ;
        RECT 83.650 405.175 118.820 405.675 ;
        RECT 122.280 405.175 154.180 405.675 ;
        RECT 5.730 404.715 41.560 405.175 ;
        RECT 44.360 404.715 80.190 405.175 ;
        RECT 82.990 404.715 118.820 405.175 ;
        RECT 121.620 404.715 154.180 405.175 ;
        RECT 5.060 404.265 41.560 404.715 ;
        RECT 43.690 404.265 80.190 404.715 ;
        RECT 82.320 404.265 118.820 404.715 ;
        RECT 120.950 404.265 154.180 404.715 ;
        RECT 4.380 403.815 41.560 404.265 ;
        RECT 43.010 403.815 80.190 404.265 ;
        RECT 81.640 403.815 118.820 404.265 ;
        RECT 120.270 403.815 154.180 404.265 ;
        RECT 3.690 403.365 41.560 403.815 ;
        RECT 42.320 403.365 80.190 403.815 ;
        RECT 80.950 403.365 118.820 403.815 ;
        RECT 119.580 403.365 154.180 403.815 ;
        RECT -1.500 0.780 154.180 403.365 ;
        RECT -1.220 -0.030 154.180 0.780 ;
      LAYER met3 ;
        RECT 9.635 389.625 151.310 390.970 ;
        RECT 9.635 386.935 151.310 388.125 ;
        RECT 9.635 383.485 151.310 385.435 ;
        RECT 9.635 380.795 151.310 381.985 ;
        RECT 9.635 377.345 151.310 379.295 ;
        RECT 9.635 374.655 151.310 375.845 ;
        RECT 9.635 371.205 151.310 373.155 ;
        RECT 9.635 368.515 151.310 369.705 ;
        RECT 9.635 365.065 151.310 367.015 ;
        RECT 9.635 362.375 151.310 363.565 ;
        RECT 9.635 358.925 151.310 360.875 ;
        RECT 9.635 356.235 151.310 357.425 ;
        RECT 9.635 352.785 151.310 354.735 ;
        RECT 9.635 350.095 151.310 351.285 ;
        RECT 9.635 346.645 151.310 348.595 ;
        RECT 9.635 343.955 151.310 345.145 ;
        RECT 9.635 340.505 151.310 342.455 ;
        RECT 9.635 337.815 151.310 339.005 ;
        RECT 9.635 334.365 151.310 336.315 ;
        RECT 9.635 331.675 151.310 332.865 ;
        RECT 9.635 328.225 151.310 330.175 ;
        RECT 9.635 325.535 151.310 326.725 ;
        RECT 9.635 322.085 151.310 324.035 ;
        RECT 9.635 319.395 151.310 320.585 ;
        RECT 9.635 315.945 151.310 317.895 ;
        RECT 9.635 313.255 151.310 314.445 ;
        RECT 9.635 309.805 151.310 311.755 ;
        RECT 9.635 307.115 151.310 308.305 ;
        RECT 9.635 303.665 151.310 305.615 ;
        RECT 9.635 300.975 151.310 302.165 ;
        RECT 9.635 297.525 151.310 299.475 ;
        RECT 9.635 294.835 151.310 296.025 ;
        RECT 9.635 291.385 151.310 293.335 ;
        RECT 9.635 288.695 151.310 289.885 ;
        RECT 9.635 285.245 151.310 287.195 ;
        RECT 9.635 282.555 151.310 283.745 ;
        RECT 9.635 279.105 151.310 281.055 ;
        RECT 9.635 276.415 151.310 277.605 ;
        RECT 9.635 272.965 151.310 274.915 ;
        RECT 9.635 270.275 151.310 271.465 ;
        RECT 9.635 266.825 151.310 268.775 ;
        RECT 9.635 264.135 151.310 265.325 ;
        RECT 9.635 260.685 151.310 262.635 ;
        RECT 9.635 257.995 151.310 259.185 ;
        RECT 9.635 254.545 151.310 256.495 ;
        RECT 9.635 251.855 151.310 253.045 ;
        RECT 9.635 248.405 151.310 250.355 ;
        RECT 9.635 245.715 151.310 246.905 ;
        RECT 9.635 242.265 151.310 244.215 ;
        RECT 9.635 239.575 151.310 240.765 ;
        RECT 9.635 236.125 151.310 238.075 ;
        RECT 9.635 233.435 151.310 234.625 ;
        RECT 9.635 229.985 151.310 231.935 ;
        RECT 9.635 227.295 151.310 228.485 ;
        RECT 9.635 223.845 151.310 225.795 ;
        RECT 9.635 221.155 151.310 222.345 ;
        RECT 9.635 217.705 151.310 219.655 ;
        RECT 9.635 215.015 151.310 216.205 ;
        RECT 9.635 211.565 151.310 213.515 ;
        RECT 9.635 208.875 151.310 210.065 ;
        RECT 9.635 205.425 151.310 207.375 ;
        RECT 9.635 202.735 151.310 203.925 ;
        RECT 9.635 199.285 151.310 201.235 ;
        RECT 9.635 196.595 151.310 197.785 ;
        RECT 9.635 193.145 151.310 195.095 ;
        RECT 9.635 190.455 151.310 191.645 ;
        RECT 9.635 187.005 151.310 188.955 ;
        RECT 9.635 184.315 151.310 185.505 ;
        RECT 9.635 180.865 151.310 182.815 ;
        RECT 9.635 178.175 151.310 179.365 ;
        RECT 9.635 174.725 151.310 176.675 ;
        RECT 9.635 172.035 151.310 173.225 ;
        RECT 9.635 168.585 151.310 170.535 ;
        RECT 9.635 165.895 151.310 167.085 ;
        RECT 9.635 162.445 151.310 164.395 ;
        RECT 9.635 159.755 151.310 160.945 ;
        RECT 9.635 156.305 151.310 158.255 ;
        RECT 9.635 153.615 151.310 154.805 ;
        RECT 9.635 150.165 151.310 152.115 ;
        RECT 9.635 147.475 151.310 148.665 ;
        RECT 9.635 144.025 151.310 145.975 ;
        RECT 9.635 141.335 151.310 142.525 ;
        RECT 9.635 137.885 151.310 139.835 ;
        RECT 9.635 135.195 151.310 136.385 ;
        RECT 9.635 131.745 151.310 133.695 ;
        RECT 9.635 129.055 151.310 130.245 ;
        RECT 9.635 125.605 151.310 127.555 ;
        RECT 9.635 122.915 151.310 124.105 ;
        RECT 9.635 119.465 151.310 121.415 ;
        RECT 9.635 116.775 151.310 117.965 ;
        RECT 9.635 113.325 151.310 115.275 ;
        RECT 9.635 110.635 151.310 111.825 ;
        RECT 9.635 107.185 151.310 109.135 ;
        RECT 9.635 104.495 151.310 105.685 ;
        RECT 9.635 101.045 151.310 102.995 ;
        RECT 9.635 98.355 151.310 99.545 ;
        RECT 9.635 94.905 151.310 96.855 ;
        RECT 9.635 92.215 151.310 93.405 ;
        RECT 9.635 88.765 151.310 90.715 ;
        RECT 9.635 86.075 151.310 87.265 ;
        RECT 9.635 82.625 151.310 84.575 ;
        RECT 9.635 79.935 151.310 81.125 ;
        RECT 9.635 76.485 151.310 78.435 ;
        RECT 9.635 73.795 151.310 74.985 ;
        RECT 9.635 70.345 151.310 72.295 ;
        RECT 9.635 67.655 151.310 68.845 ;
        RECT 9.635 64.205 151.310 66.155 ;
        RECT 9.635 61.515 151.310 62.705 ;
        RECT 9.635 58.065 151.310 60.015 ;
        RECT 9.635 55.375 151.310 56.565 ;
        RECT 9.635 51.925 151.310 53.875 ;
        RECT 9.635 49.235 151.310 50.425 ;
        RECT 9.635 45.785 151.310 47.735 ;
        RECT 9.635 43.095 151.310 44.285 ;
        RECT 9.635 39.645 151.310 41.595 ;
        RECT 9.635 36.955 151.310 38.145 ;
        RECT 9.635 33.505 151.310 35.455 ;
        RECT 9.635 30.815 151.310 32.005 ;
        RECT 9.635 27.365 151.310 29.315 ;
        RECT 9.635 24.675 151.310 25.865 ;
        RECT 9.635 21.225 151.310 23.175 ;
        RECT 9.635 18.535 151.310 19.725 ;
        RECT 9.635 15.085 151.310 17.035 ;
        RECT 9.635 12.395 151.310 13.585 ;
        RECT 9.635 8.945 151.310 10.895 ;
        RECT 9.635 6.255 151.310 7.445 ;
        RECT 9.635 2.805 151.310 4.755 ;
  END
END dac_top
END LIBRARY

