magic
tech sky130A
magscale 1 2
timestamp 1686240839
<< nwell >>
rect -1666 1758 -884 2034
rect -1580 1520 -920 1758
rect -1976 1034 -1498 1219
rect -1934 754 -1506 1034
<< pwell >>
rect -1454 650 -1028 1316
rect -1924 462 -1028 650
rect -1927 322 -1008 462
<< nmos >>
rect -1840 540 -1810 624
rect -1630 540 -1600 624
<< pmos >>
rect -1840 816 -1810 984
rect -1630 816 -1600 984
<< mvnmos >>
rect -1370 490 -1270 1290
rect -1212 490 -1112 1290
<< mvpmos >>
rect -1446 1590 -1346 1790
rect -1158 1590 -1058 1790
<< ndiff >>
rect -1898 599 -1840 624
rect -1898 565 -1886 599
rect -1852 565 -1840 599
rect -1898 540 -1840 565
rect -1810 599 -1752 624
rect -1810 565 -1798 599
rect -1764 565 -1752 599
rect -1810 540 -1752 565
rect -1688 599 -1630 624
rect -1688 565 -1676 599
rect -1642 565 -1630 599
rect -1688 540 -1630 565
rect -1600 599 -1542 624
rect -1600 565 -1588 599
rect -1554 565 -1542 599
rect -1600 540 -1542 565
<< pdiff >>
rect -1898 951 -1840 984
rect -1898 917 -1886 951
rect -1852 917 -1840 951
rect -1898 883 -1840 917
rect -1898 849 -1886 883
rect -1852 849 -1840 883
rect -1898 816 -1840 849
rect -1810 951 -1752 984
rect -1810 917 -1798 951
rect -1764 917 -1752 951
rect -1810 883 -1752 917
rect -1810 849 -1798 883
rect -1764 849 -1752 883
rect -1810 816 -1752 849
rect -1688 951 -1630 984
rect -1688 917 -1676 951
rect -1642 917 -1630 951
rect -1688 883 -1630 917
rect -1688 849 -1676 883
rect -1642 849 -1630 883
rect -1688 816 -1630 849
rect -1600 951 -1542 984
rect -1600 917 -1588 951
rect -1554 917 -1542 951
rect -1600 883 -1542 917
rect -1600 849 -1588 883
rect -1554 849 -1542 883
rect -1600 816 -1542 849
<< mvndiff >>
rect -1428 1247 -1370 1290
rect -1428 1213 -1416 1247
rect -1382 1213 -1370 1247
rect -1428 1179 -1370 1213
rect -1428 1145 -1416 1179
rect -1382 1145 -1370 1179
rect -1428 1111 -1370 1145
rect -1428 1077 -1416 1111
rect -1382 1077 -1370 1111
rect -1428 1043 -1370 1077
rect -1428 1009 -1416 1043
rect -1382 1009 -1370 1043
rect -1428 975 -1370 1009
rect -1428 941 -1416 975
rect -1382 941 -1370 975
rect -1428 907 -1370 941
rect -1428 873 -1416 907
rect -1382 873 -1370 907
rect -1428 839 -1370 873
rect -1428 805 -1416 839
rect -1382 805 -1370 839
rect -1428 771 -1370 805
rect -1428 737 -1416 771
rect -1382 737 -1370 771
rect -1428 703 -1370 737
rect -1428 669 -1416 703
rect -1382 669 -1370 703
rect -1428 635 -1370 669
rect -1428 601 -1416 635
rect -1382 601 -1370 635
rect -1428 567 -1370 601
rect -1428 533 -1416 567
rect -1382 533 -1370 567
rect -1428 490 -1370 533
rect -1270 1247 -1212 1290
rect -1270 1213 -1258 1247
rect -1224 1213 -1212 1247
rect -1270 1179 -1212 1213
rect -1270 1145 -1258 1179
rect -1224 1145 -1212 1179
rect -1270 1111 -1212 1145
rect -1270 1077 -1258 1111
rect -1224 1077 -1212 1111
rect -1270 1043 -1212 1077
rect -1270 1009 -1258 1043
rect -1224 1009 -1212 1043
rect -1270 975 -1212 1009
rect -1270 941 -1258 975
rect -1224 941 -1212 975
rect -1270 907 -1212 941
rect -1270 873 -1258 907
rect -1224 873 -1212 907
rect -1270 839 -1212 873
rect -1270 805 -1258 839
rect -1224 805 -1212 839
rect -1270 771 -1212 805
rect -1270 737 -1258 771
rect -1224 737 -1212 771
rect -1270 703 -1212 737
rect -1270 669 -1258 703
rect -1224 669 -1212 703
rect -1270 635 -1212 669
rect -1270 601 -1258 635
rect -1224 601 -1212 635
rect -1270 567 -1212 601
rect -1270 533 -1258 567
rect -1224 533 -1212 567
rect -1270 490 -1212 533
rect -1112 1247 -1054 1290
rect -1112 1213 -1100 1247
rect -1066 1213 -1054 1247
rect -1112 1179 -1054 1213
rect -1112 1145 -1100 1179
rect -1066 1145 -1054 1179
rect -1112 1111 -1054 1145
rect -1112 1077 -1100 1111
rect -1066 1077 -1054 1111
rect -1112 1043 -1054 1077
rect -1112 1009 -1100 1043
rect -1066 1009 -1054 1043
rect -1112 975 -1054 1009
rect -1112 941 -1100 975
rect -1066 941 -1054 975
rect -1112 907 -1054 941
rect -1112 873 -1100 907
rect -1066 873 -1054 907
rect -1112 839 -1054 873
rect -1112 805 -1100 839
rect -1066 805 -1054 839
rect -1112 771 -1054 805
rect -1112 737 -1100 771
rect -1066 737 -1054 771
rect -1112 703 -1054 737
rect -1112 669 -1100 703
rect -1066 669 -1054 703
rect -1112 635 -1054 669
rect -1112 601 -1100 635
rect -1066 601 -1054 635
rect -1112 567 -1054 601
rect -1112 533 -1100 567
rect -1066 533 -1054 567
rect -1112 490 -1054 533
<< mvpdiff >>
rect -1504 1775 -1446 1790
rect -1504 1741 -1492 1775
rect -1458 1741 -1446 1775
rect -1504 1707 -1446 1741
rect -1504 1673 -1492 1707
rect -1458 1673 -1446 1707
rect -1504 1639 -1446 1673
rect -1504 1605 -1492 1639
rect -1458 1605 -1446 1639
rect -1504 1590 -1446 1605
rect -1346 1775 -1288 1790
rect -1346 1741 -1334 1775
rect -1300 1741 -1288 1775
rect -1346 1707 -1288 1741
rect -1346 1673 -1334 1707
rect -1300 1673 -1288 1707
rect -1346 1639 -1288 1673
rect -1346 1605 -1334 1639
rect -1300 1605 -1288 1639
rect -1346 1590 -1288 1605
rect -1216 1775 -1158 1790
rect -1216 1741 -1204 1775
rect -1170 1741 -1158 1775
rect -1216 1707 -1158 1741
rect -1216 1673 -1204 1707
rect -1170 1673 -1158 1707
rect -1216 1639 -1158 1673
rect -1216 1605 -1204 1639
rect -1170 1605 -1158 1639
rect -1216 1590 -1158 1605
rect -1058 1775 -1000 1790
rect -1058 1741 -1046 1775
rect -1012 1741 -1000 1775
rect -1058 1707 -1000 1741
rect -1058 1673 -1046 1707
rect -1012 1673 -1000 1707
rect -1058 1639 -1000 1673
rect -1058 1605 -1046 1639
rect -1012 1605 -1000 1639
rect -1058 1590 -1000 1605
<< ndiffc >>
rect -1886 565 -1852 599
rect -1798 565 -1764 599
rect -1676 565 -1642 599
rect -1588 565 -1554 599
<< pdiffc >>
rect -1886 917 -1852 951
rect -1886 849 -1852 883
rect -1798 917 -1764 951
rect -1798 849 -1764 883
rect -1676 917 -1642 951
rect -1676 849 -1642 883
rect -1588 917 -1554 951
rect -1588 849 -1554 883
<< mvndiffc >>
rect -1416 1213 -1382 1247
rect -1416 1145 -1382 1179
rect -1416 1077 -1382 1111
rect -1416 1009 -1382 1043
rect -1416 941 -1382 975
rect -1416 873 -1382 907
rect -1416 805 -1382 839
rect -1416 737 -1382 771
rect -1416 669 -1382 703
rect -1416 601 -1382 635
rect -1416 533 -1382 567
rect -1258 1213 -1224 1247
rect -1258 1145 -1224 1179
rect -1258 1077 -1224 1111
rect -1258 1009 -1224 1043
rect -1258 941 -1224 975
rect -1258 873 -1224 907
rect -1258 805 -1224 839
rect -1258 737 -1224 771
rect -1258 669 -1224 703
rect -1258 601 -1224 635
rect -1258 533 -1224 567
rect -1100 1213 -1066 1247
rect -1100 1145 -1066 1179
rect -1100 1077 -1066 1111
rect -1100 1009 -1066 1043
rect -1100 941 -1066 975
rect -1100 873 -1066 907
rect -1100 805 -1066 839
rect -1100 737 -1066 771
rect -1100 669 -1066 703
rect -1100 601 -1066 635
rect -1100 533 -1066 567
<< mvpdiffc >>
rect -1492 1741 -1458 1775
rect -1492 1673 -1458 1707
rect -1492 1605 -1458 1639
rect -1334 1741 -1300 1775
rect -1334 1673 -1300 1707
rect -1334 1605 -1300 1639
rect -1204 1741 -1170 1775
rect -1204 1673 -1170 1707
rect -1204 1605 -1170 1639
rect -1046 1741 -1012 1775
rect -1046 1673 -1012 1707
rect -1046 1605 -1012 1639
<< psubdiff >>
rect -1901 405 -1034 436
rect -1901 371 -1859 405
rect -1825 371 -1791 405
rect -1757 371 -1723 405
rect -1689 371 -1655 405
rect -1621 371 -1587 405
rect -1553 371 -1519 405
rect -1485 371 -1451 405
rect -1417 371 -1383 405
rect -1349 371 -1315 405
rect -1281 371 -1247 405
rect -1213 371 -1179 405
rect -1145 371 -1111 405
rect -1077 371 -1034 405
rect -1901 348 -1034 371
<< nsubdiff >>
rect -1935 1143 -1538 1179
rect -1935 1109 -1889 1143
rect -1855 1109 -1821 1143
rect -1787 1109 -1753 1143
rect -1719 1109 -1685 1143
rect -1651 1109 -1617 1143
rect -1583 1109 -1538 1143
rect -1935 1081 -1538 1109
<< mvnsubdiff >>
rect -1568 1911 -957 1944
rect -1568 1877 -1522 1911
rect -1488 1877 -1454 1911
rect -1420 1877 -1386 1911
rect -1352 1877 -1318 1911
rect -1284 1877 -1250 1911
rect -1216 1877 -1182 1911
rect -1148 1877 -1114 1911
rect -1080 1877 -1046 1911
rect -1012 1877 -957 1911
rect -1568 1850 -957 1877
<< psubdiffcont >>
rect -1859 371 -1825 405
rect -1791 371 -1757 405
rect -1723 371 -1689 405
rect -1655 371 -1621 405
rect -1587 371 -1553 405
rect -1519 371 -1485 405
rect -1451 371 -1417 405
rect -1383 371 -1349 405
rect -1315 371 -1281 405
rect -1247 371 -1213 405
rect -1179 371 -1145 405
rect -1111 371 -1077 405
<< nsubdiffcont >>
rect -1889 1109 -1855 1143
rect -1821 1109 -1787 1143
rect -1753 1109 -1719 1143
rect -1685 1109 -1651 1143
rect -1617 1109 -1583 1143
<< mvnsubdiffcont >>
rect -1522 1877 -1488 1911
rect -1454 1877 -1420 1911
rect -1386 1877 -1352 1911
rect -1318 1877 -1284 1911
rect -1250 1877 -1216 1911
rect -1182 1877 -1148 1911
rect -1114 1877 -1080 1911
rect -1046 1877 -1012 1911
<< poly >>
rect -1446 1790 -1346 1816
rect -1158 1790 -1058 1816
rect -1446 1564 -1346 1590
rect -1158 1564 -1058 1590
rect -1424 1493 -1376 1564
rect -1433 1483 -1367 1493
rect -1126 1492 -1081 1564
rect -1433 1449 -1417 1483
rect -1383 1449 -1367 1483
rect -1433 1439 -1367 1449
rect -1136 1482 -1070 1492
rect -1136 1448 -1120 1482
rect -1086 1448 -1070 1482
rect -1136 1438 -1070 1448
rect -1533 1397 -1467 1407
rect -1533 1363 -1517 1397
rect -1483 1363 -1303 1397
rect -1533 1353 -1467 1363
rect -1337 1316 -1303 1363
rect -1212 1350 -1114 1351
rect -1013 1350 -947 1357
rect -1212 1347 -947 1350
rect -1370 1290 -1270 1316
rect -1212 1313 -997 1347
rect -963 1313 -947 1347
rect -1212 1310 -947 1313
rect -1212 1290 -1112 1310
rect -1013 1303 -947 1310
rect -1840 984 -1810 1010
rect -1630 984 -1600 1010
rect -2020 731 -1954 741
rect -2020 697 -2004 731
rect -1970 729 -1954 731
rect -1840 729 -1810 816
rect -1970 699 -1810 729
rect -1970 697 -1954 699
rect -2020 687 -1954 697
rect -1840 624 -1810 699
rect -1743 737 -1677 747
rect -1743 703 -1727 737
rect -1693 735 -1677 737
rect -1630 735 -1600 816
rect -1693 705 -1600 735
rect -1693 703 -1677 705
rect -1743 693 -1677 703
rect -1630 624 -1600 705
rect -1840 514 -1810 540
rect -1630 514 -1600 540
rect -1370 464 -1270 490
rect -1212 464 -1112 490
<< polycont >>
rect -1417 1449 -1383 1483
rect -1120 1448 -1086 1482
rect -1517 1363 -1483 1397
rect -997 1313 -963 1347
rect -2004 697 -1970 731
rect -1727 703 -1693 737
<< locali >>
rect -1568 1911 -957 1944
rect -1568 1877 -1536 1911
rect -1488 1877 -1464 1911
rect -1420 1877 -1392 1911
rect -1352 1877 -1320 1911
rect -1284 1877 -1250 1911
rect -1214 1877 -1182 1911
rect -1142 1877 -1114 1911
rect -1070 1877 -1046 1911
rect -998 1877 -957 1911
rect -1568 1850 -957 1877
rect -1492 1775 -1458 1794
rect -1492 1707 -1458 1709
rect -1492 1671 -1458 1673
rect -1334 1775 -1300 1794
rect -1334 1707 -1300 1709
rect -1334 1672 -1300 1673
rect -1204 1775 -1170 1794
rect -1204 1707 -1170 1709
rect -1492 1586 -1458 1605
rect -1336 1671 -1291 1672
rect -1336 1605 -1334 1671
rect -1300 1605 -1291 1671
rect -1417 1490 -1383 1499
rect -1424 1483 -1376 1490
rect -1424 1449 -1417 1483
rect -1383 1449 -1376 1483
rect -1424 1442 -1376 1449
rect -1336 1488 -1291 1605
rect -1204 1671 -1170 1673
rect -1204 1586 -1170 1605
rect -1046 1775 -1012 1794
rect -1046 1707 -1012 1709
rect -1046 1671 -1012 1673
rect -1046 1586 -1012 1605
rect -1120 1488 -1086 1498
rect -1336 1482 -1080 1488
rect -1336 1448 -1120 1482
rect -1086 1448 -1080 1482
rect -1336 1443 -1080 1448
rect -1417 1433 -1383 1442
rect -1517 1397 -1483 1413
rect -1336 1365 -1291 1443
rect -1120 1432 -1086 1443
rect -1517 1347 -1483 1363
rect -1426 1320 -1291 1365
rect -997 1350 -963 1363
rect -1000 1347 -960 1350
rect -1426 1267 -1381 1320
rect -1000 1313 -997 1347
rect -963 1313 -960 1347
rect -1000 1310 -960 1313
rect -997 1297 -963 1310
rect -1426 1213 -1416 1267
rect -1382 1213 -1381 1267
rect -1426 1195 -1381 1213
rect -1426 1182 -1416 1195
rect -1382 1182 -1381 1195
rect -1258 1267 -1224 1294
rect -1258 1195 -1224 1213
rect -1935 1143 -1538 1179
rect -1935 1109 -1897 1143
rect -1855 1109 -1825 1143
rect -1787 1109 -1753 1143
rect -1719 1109 -1685 1143
rect -1647 1109 -1617 1143
rect -1575 1109 -1538 1143
rect -1935 1081 -1538 1109
rect -1416 1123 -1382 1145
rect -1416 1051 -1382 1077
rect -1886 953 -1852 988
rect -1886 883 -1852 917
rect -1886 812 -1852 847
rect -1798 953 -1764 988
rect -1798 883 -1764 917
rect -1798 812 -1764 847
rect -1676 953 -1642 988
rect -1676 883 -1642 917
rect -1676 812 -1642 847
rect -1588 953 -1554 988
rect -1588 883 -1554 917
rect -1588 812 -1554 847
rect -1416 979 -1382 1009
rect -1416 907 -1382 941
rect -1416 839 -1382 873
rect -1416 771 -1382 801
rect -2004 731 -1970 747
rect -2004 681 -1970 697
rect -1727 737 -1693 753
rect -1727 687 -1693 703
rect -1416 703 -1382 729
rect -1416 635 -1382 657
rect -1886 599 -1852 628
rect -1886 536 -1852 565
rect -1798 599 -1764 628
rect -1798 536 -1764 565
rect -1676 599 -1642 628
rect -1676 536 -1642 565
rect -1588 599 -1554 628
rect -1588 536 -1554 565
rect -1416 567 -1382 585
rect -1416 486 -1382 513
rect -1258 1123 -1224 1145
rect -1258 1051 -1224 1077
rect -1258 979 -1224 1009
rect -1258 907 -1224 941
rect -1258 839 -1224 873
rect -1258 771 -1224 801
rect -1258 703 -1224 729
rect -1258 635 -1224 657
rect -1258 567 -1224 585
rect -1258 486 -1224 513
rect -1100 1267 -1066 1294
rect -1100 1195 -1066 1213
rect -1100 1123 -1066 1145
rect -1100 1051 -1066 1077
rect -1100 979 -1066 1009
rect -1100 907 -1066 941
rect -1100 839 -1066 873
rect -1100 771 -1066 801
rect -1100 703 -1066 729
rect -1100 635 -1066 657
rect -1100 567 -1066 585
rect -1100 486 -1066 513
rect -1901 405 -1033 448
rect -1901 371 -1859 405
rect -1811 371 -1791 405
rect -1739 371 -1723 405
rect -1667 371 -1655 405
rect -1595 371 -1587 405
rect -1523 371 -1519 405
rect -1417 371 -1413 405
rect -1349 371 -1341 405
rect -1281 371 -1269 405
rect -1213 371 -1197 405
rect -1145 371 -1125 405
rect -1077 371 -1033 405
rect -1901 348 -1033 371
<< viali >>
rect -1536 1877 -1522 1911
rect -1522 1877 -1502 1911
rect -1464 1877 -1454 1911
rect -1454 1877 -1430 1911
rect -1392 1877 -1386 1911
rect -1386 1877 -1358 1911
rect -1320 1877 -1318 1911
rect -1318 1877 -1286 1911
rect -1248 1877 -1216 1911
rect -1216 1877 -1214 1911
rect -1176 1877 -1148 1911
rect -1148 1877 -1142 1911
rect -1104 1877 -1080 1911
rect -1080 1877 -1070 1911
rect -1032 1877 -1012 1911
rect -1012 1877 -998 1911
rect -1492 1741 -1458 1743
rect -1492 1709 -1458 1741
rect -1334 1741 -1300 1743
rect -1334 1709 -1300 1741
rect -1204 1741 -1170 1743
rect -1204 1709 -1170 1741
rect -1492 1639 -1458 1671
rect -1492 1637 -1458 1639
rect -1334 1639 -1300 1671
rect -1334 1637 -1300 1639
rect -1417 1449 -1383 1483
rect -1204 1639 -1170 1671
rect -1204 1637 -1170 1639
rect -1046 1741 -1012 1743
rect -1046 1709 -1012 1741
rect -1046 1639 -1012 1671
rect -1046 1637 -1012 1639
rect -1517 1363 -1483 1397
rect -997 1313 -963 1347
rect -1416 1247 -1382 1267
rect -1416 1233 -1382 1247
rect -1416 1179 -1382 1195
rect -1258 1247 -1224 1267
rect -1258 1233 -1224 1247
rect -1897 1109 -1889 1143
rect -1889 1109 -1863 1143
rect -1825 1109 -1821 1143
rect -1821 1109 -1791 1143
rect -1753 1109 -1719 1143
rect -1681 1109 -1651 1143
rect -1651 1109 -1647 1143
rect -1609 1109 -1583 1143
rect -1583 1109 -1575 1143
rect -1416 1161 -1382 1179
rect -1416 1111 -1382 1123
rect -1416 1089 -1382 1111
rect -1416 1043 -1382 1051
rect -1416 1017 -1382 1043
rect -1886 951 -1852 953
rect -1886 919 -1852 951
rect -1886 849 -1852 881
rect -1886 847 -1852 849
rect -1798 951 -1764 953
rect -1798 919 -1764 951
rect -1798 849 -1764 881
rect -1798 847 -1764 849
rect -1676 951 -1642 953
rect -1676 919 -1642 951
rect -1676 849 -1642 881
rect -1676 847 -1642 849
rect -1588 951 -1554 953
rect -1588 919 -1554 951
rect -1588 849 -1554 881
rect -1588 847 -1554 849
rect -1416 975 -1382 979
rect -1416 945 -1382 975
rect -1416 873 -1382 907
rect -1416 805 -1382 835
rect -1416 801 -1382 805
rect -2004 697 -1970 731
rect -1727 703 -1693 737
rect -1416 737 -1382 763
rect -1416 729 -1382 737
rect -1416 669 -1382 691
rect -1416 657 -1382 669
rect -1886 565 -1852 599
rect -1798 565 -1764 599
rect -1676 565 -1642 599
rect -1588 565 -1554 599
rect -1416 601 -1382 619
rect -1416 585 -1382 601
rect -1416 533 -1382 547
rect -1416 513 -1382 533
rect -1258 1179 -1224 1195
rect -1258 1161 -1224 1179
rect -1258 1111 -1224 1123
rect -1258 1089 -1224 1111
rect -1258 1043 -1224 1051
rect -1258 1017 -1224 1043
rect -1258 975 -1224 979
rect -1258 945 -1224 975
rect -1258 873 -1224 907
rect -1258 805 -1224 835
rect -1258 801 -1224 805
rect -1258 737 -1224 763
rect -1258 729 -1224 737
rect -1258 669 -1224 691
rect -1258 657 -1224 669
rect -1258 601 -1224 619
rect -1258 585 -1224 601
rect -1258 533 -1224 547
rect -1258 513 -1224 533
rect -1100 1247 -1066 1267
rect -1100 1233 -1066 1247
rect -1100 1179 -1066 1195
rect -1100 1161 -1066 1179
rect -1100 1111 -1066 1123
rect -1100 1089 -1066 1111
rect -1100 1043 -1066 1051
rect -1100 1017 -1066 1043
rect -1100 975 -1066 979
rect -1100 945 -1066 975
rect -1100 873 -1066 907
rect -1100 805 -1066 835
rect -1100 801 -1066 805
rect -1100 737 -1066 763
rect -1100 729 -1066 737
rect -1100 669 -1066 691
rect -1100 657 -1066 669
rect -1100 601 -1066 619
rect -1100 585 -1066 601
rect -1100 533 -1066 547
rect -1100 513 -1066 533
rect -1845 371 -1825 405
rect -1825 371 -1811 405
rect -1773 371 -1757 405
rect -1757 371 -1739 405
rect -1701 371 -1689 405
rect -1689 371 -1667 405
rect -1629 371 -1621 405
rect -1621 371 -1595 405
rect -1557 371 -1553 405
rect -1553 371 -1523 405
rect -1485 371 -1451 405
rect -1413 371 -1383 405
rect -1383 371 -1379 405
rect -1341 371 -1315 405
rect -1315 371 -1307 405
rect -1269 371 -1247 405
rect -1247 371 -1235 405
rect -1197 371 -1179 405
rect -1179 371 -1163 405
rect -1125 371 -1111 405
rect -1111 371 -1091 405
<< metal1 >>
rect -1568 1923 -957 1944
rect -1568 1911 -1517 1923
rect -1465 1911 -1453 1923
rect -1401 1911 -1389 1923
rect -1568 1877 -1536 1911
rect -1465 1877 -1464 1911
rect -1401 1877 -1392 1911
rect -1568 1871 -1517 1877
rect -1465 1871 -1453 1877
rect -1401 1871 -1389 1877
rect -1337 1871 -1325 1923
rect -1273 1871 -1261 1923
rect -1209 1871 -1197 1923
rect -1145 1911 -1133 1923
rect -1081 1911 -1069 1923
rect -1017 1911 -957 1923
rect -1142 1877 -1133 1911
rect -1070 1877 -1069 1911
rect -998 1877 -957 1911
rect -1145 1871 -1133 1877
rect -1081 1871 -1069 1877
rect -1017 1871 -957 1877
rect -1568 1850 -957 1871
rect -1501 1783 -1450 1850
rect -1498 1743 -1452 1783
rect -1498 1709 -1492 1743
rect -1458 1709 -1452 1743
rect -1498 1671 -1452 1709
rect -1498 1637 -1492 1671
rect -1458 1637 -1452 1671
rect -1498 1590 -1452 1637
rect -1340 1743 -1294 1790
rect -1340 1709 -1334 1743
rect -1300 1709 -1294 1743
rect -1340 1671 -1294 1709
rect -1340 1637 -1334 1671
rect -1300 1637 -1294 1671
rect -1210 1743 -1164 1790
rect -1054 1780 -1003 1850
rect -1210 1709 -1204 1743
rect -1170 1709 -1164 1743
rect -1210 1671 -1164 1709
rect -1210 1658 -1204 1671
rect -1340 1590 -1294 1637
rect -1214 1637 -1204 1658
rect -1170 1637 -1164 1671
rect -1214 1590 -1164 1637
rect -1052 1743 -1006 1780
rect -1052 1709 -1046 1743
rect -1012 1709 -1006 1743
rect -1052 1671 -1006 1709
rect -1052 1637 -1046 1671
rect -1012 1637 -1006 1671
rect -1052 1590 -1006 1637
rect -1430 1490 -1370 1502
rect -1214 1490 -1166 1590
rect -1430 1483 -1166 1490
rect -1430 1449 -1417 1483
rect -1383 1449 -1166 1483
rect -1430 1442 -1166 1449
rect -1430 1430 -1370 1442
rect -1523 1397 -1464 1409
rect -1537 1363 -1517 1397
rect -1483 1363 -1464 1397
rect -1523 1351 -1464 1363
rect -2013 1312 -1961 1318
rect -2013 1254 -1961 1260
rect -2004 743 -1970 1254
rect -1935 1157 -1538 1178
rect -1935 1143 -1890 1157
rect -1935 1109 -1897 1143
rect -1935 1105 -1890 1109
rect -1838 1105 -1826 1157
rect -1774 1105 -1762 1157
rect -1710 1105 -1698 1157
rect -1646 1105 -1634 1157
rect -1582 1143 -1538 1157
rect -1575 1109 -1538 1143
rect -1582 1105 -1538 1109
rect -1935 1081 -1538 1105
rect -1889 984 -1849 1081
rect -1797 984 -1763 988
rect -1679 984 -1639 1081
rect -1892 953 -1846 984
rect -1892 919 -1886 953
rect -1852 919 -1846 953
rect -1892 881 -1846 919
rect -1892 847 -1886 881
rect -1852 847 -1846 881
rect -1892 816 -1846 847
rect -1804 953 -1758 984
rect -1804 919 -1798 953
rect -1764 919 -1758 953
rect -1804 881 -1758 919
rect -1804 847 -1798 881
rect -1764 847 -1758 881
rect -1804 816 -1758 847
rect -1682 953 -1636 984
rect -1682 919 -1676 953
rect -1642 919 -1636 953
rect -1682 881 -1636 919
rect -1682 847 -1676 881
rect -1642 847 -1636 881
rect -1682 816 -1636 847
rect -1594 963 -1548 984
rect -1498 963 -1464 1351
rect -1214 1368 -1166 1442
rect -1214 1320 -1062 1368
rect -1006 1356 -954 1362
rect -1110 1290 -1062 1320
rect -1012 1304 -1006 1356
rect -954 1304 -948 1356
rect -1006 1298 -954 1304
rect -1594 953 -1464 963
rect -1594 919 -1588 953
rect -1554 927 -1464 953
rect -1422 1267 -1376 1290
rect -1422 1233 -1416 1267
rect -1382 1233 -1376 1267
rect -1422 1195 -1376 1233
rect -1422 1161 -1416 1195
rect -1382 1161 -1376 1195
rect -1422 1123 -1376 1161
rect -1422 1089 -1416 1123
rect -1382 1089 -1376 1123
rect -1422 1051 -1376 1089
rect -1422 1017 -1416 1051
rect -1382 1017 -1376 1051
rect -1422 979 -1376 1017
rect -1422 945 -1416 979
rect -1382 945 -1376 979
rect -1554 919 -1548 927
rect -1594 881 -1548 919
rect -1594 847 -1588 881
rect -1554 847 -1548 881
rect -1594 816 -1548 847
rect -1422 907 -1376 945
rect -1422 873 -1416 907
rect -1382 873 -1376 907
rect -1422 835 -1376 873
rect -2010 731 -1964 743
rect -2010 697 -2004 731
rect -1970 697 -1964 731
rect -2010 685 -1964 697
rect -1797 737 -1763 816
rect -1733 746 -1687 749
rect -1733 737 -1715 746
rect -1797 703 -1727 737
rect -1797 624 -1763 703
rect -1733 694 -1715 703
rect -1663 694 -1657 746
rect -1733 691 -1687 694
rect -1587 624 -1553 816
rect -1422 801 -1416 835
rect -1382 801 -1376 835
rect -1422 763 -1376 801
rect -1422 729 -1416 763
rect -1382 729 -1376 763
rect -1422 691 -1376 729
rect -1422 657 -1416 691
rect -1382 657 -1376 691
rect -1892 599 -1846 624
rect -1892 565 -1886 599
rect -1852 565 -1846 599
rect -1892 540 -1846 565
rect -1804 599 -1758 624
rect -1804 565 -1798 599
rect -1764 565 -1758 599
rect -1804 540 -1758 565
rect -1682 599 -1636 624
rect -1682 565 -1676 599
rect -1642 565 -1636 599
rect -1682 540 -1636 565
rect -1594 599 -1548 624
rect -1594 565 -1588 599
rect -1554 565 -1548 599
rect -1594 540 -1548 565
rect -1422 619 -1376 657
rect -1422 585 -1416 619
rect -1382 585 -1376 619
rect -1422 547 -1376 585
rect -1887 448 -1854 540
rect -1674 448 -1641 540
rect -1422 513 -1416 547
rect -1382 513 -1376 547
rect -1422 490 -1376 513
rect -1264 1267 -1218 1290
rect -1264 1233 -1258 1267
rect -1224 1233 -1218 1267
rect -1264 1195 -1218 1233
rect -1264 1161 -1258 1195
rect -1224 1161 -1218 1195
rect -1264 1123 -1218 1161
rect -1264 1089 -1258 1123
rect -1224 1089 -1218 1123
rect -1264 1051 -1218 1089
rect -1264 1017 -1258 1051
rect -1224 1017 -1218 1051
rect -1264 979 -1218 1017
rect -1264 945 -1258 979
rect -1224 945 -1218 979
rect -1264 907 -1218 945
rect -1264 873 -1258 907
rect -1224 873 -1218 907
rect -1264 835 -1218 873
rect -1264 801 -1258 835
rect -1224 801 -1218 835
rect -1264 763 -1218 801
rect -1264 729 -1258 763
rect -1224 729 -1218 763
rect -1264 691 -1218 729
rect -1264 657 -1258 691
rect -1224 657 -1218 691
rect -1264 619 -1218 657
rect -1264 585 -1258 619
rect -1224 585 -1218 619
rect -1264 547 -1218 585
rect -1110 1267 -1060 1290
rect -1110 1233 -1100 1267
rect -1066 1233 -1060 1267
rect -1110 1195 -1060 1233
rect -1110 1161 -1100 1195
rect -1066 1161 -1060 1195
rect -1110 1123 -1060 1161
rect -1110 1089 -1100 1123
rect -1066 1089 -1060 1123
rect -1110 1051 -1060 1089
rect -1110 1017 -1100 1051
rect -1066 1017 -1060 1051
rect -1110 979 -1060 1017
rect -1110 945 -1100 979
rect -1066 945 -1060 979
rect -1110 907 -1060 945
rect -1110 873 -1100 907
rect -1066 873 -1060 907
rect -1110 835 -1060 873
rect -1110 801 -1100 835
rect -1066 801 -1060 835
rect -1110 763 -1060 801
rect -1110 729 -1100 763
rect -1066 729 -1060 763
rect -1110 691 -1060 729
rect -1110 657 -1100 691
rect -1066 657 -1060 691
rect -1110 619 -1060 657
rect -1110 585 -1100 619
rect -1066 585 -1060 619
rect -1110 577 -1060 585
rect -1264 513 -1258 547
rect -1224 513 -1218 547
rect -1115 574 -936 577
rect -1115 547 -997 574
rect -1115 519 -1100 547
rect -1264 490 -1218 513
rect -1106 513 -1100 519
rect -1066 522 -997 547
rect -945 522 -936 574
rect -1066 519 -936 522
rect -1066 513 -1060 519
rect -1106 490 -1060 513
rect -1258 448 -1219 490
rect -1901 414 -1033 448
rect -1901 362 -1846 414
rect -1794 362 -1782 414
rect -1730 362 -1718 414
rect -1666 362 -1654 414
rect -1602 405 -1590 414
rect -1538 405 -1526 414
rect -1474 405 -1462 414
rect -1410 405 -1398 414
rect -1346 405 -1334 414
rect -1595 371 -1590 405
rect -1346 371 -1341 405
rect -1602 362 -1590 371
rect -1538 362 -1526 371
rect -1474 362 -1462 371
rect -1410 362 -1398 371
rect -1346 362 -1334 371
rect -1282 362 -1270 414
rect -1218 362 -1206 414
rect -1154 362 -1142 414
rect -1090 362 -1033 414
rect -1901 348 -1033 362
<< via1 >>
rect -1517 1911 -1465 1923
rect -1453 1911 -1401 1923
rect -1389 1911 -1337 1923
rect -1517 1877 -1502 1911
rect -1502 1877 -1465 1911
rect -1453 1877 -1430 1911
rect -1430 1877 -1401 1911
rect -1389 1877 -1358 1911
rect -1358 1877 -1337 1911
rect -1517 1871 -1465 1877
rect -1453 1871 -1401 1877
rect -1389 1871 -1337 1877
rect -1325 1911 -1273 1923
rect -1325 1877 -1320 1911
rect -1320 1877 -1286 1911
rect -1286 1877 -1273 1911
rect -1325 1871 -1273 1877
rect -1261 1911 -1209 1923
rect -1261 1877 -1248 1911
rect -1248 1877 -1214 1911
rect -1214 1877 -1209 1911
rect -1261 1871 -1209 1877
rect -1197 1911 -1145 1923
rect -1133 1911 -1081 1923
rect -1069 1911 -1017 1923
rect -1197 1877 -1176 1911
rect -1176 1877 -1145 1911
rect -1133 1877 -1104 1911
rect -1104 1877 -1081 1911
rect -1069 1877 -1032 1911
rect -1032 1877 -1017 1911
rect -1197 1871 -1145 1877
rect -1133 1871 -1081 1877
rect -1069 1871 -1017 1877
rect -2013 1260 -1961 1312
rect -1890 1143 -1838 1157
rect -1890 1109 -1863 1143
rect -1863 1109 -1838 1143
rect -1890 1105 -1838 1109
rect -1826 1143 -1774 1157
rect -1826 1109 -1825 1143
rect -1825 1109 -1791 1143
rect -1791 1109 -1774 1143
rect -1826 1105 -1774 1109
rect -1762 1143 -1710 1157
rect -1762 1109 -1753 1143
rect -1753 1109 -1719 1143
rect -1719 1109 -1710 1143
rect -1762 1105 -1710 1109
rect -1698 1143 -1646 1157
rect -1698 1109 -1681 1143
rect -1681 1109 -1647 1143
rect -1647 1109 -1646 1143
rect -1698 1105 -1646 1109
rect -1634 1143 -1582 1157
rect -1634 1109 -1609 1143
rect -1609 1109 -1582 1143
rect -1634 1105 -1582 1109
rect -1006 1347 -954 1356
rect -1006 1313 -997 1347
rect -997 1313 -963 1347
rect -963 1313 -954 1347
rect -1006 1304 -954 1313
rect -1715 737 -1663 746
rect -1715 703 -1693 737
rect -1693 703 -1663 737
rect -1715 694 -1663 703
rect -997 522 -945 574
rect -1846 405 -1794 414
rect -1846 371 -1845 405
rect -1845 371 -1811 405
rect -1811 371 -1794 405
rect -1846 362 -1794 371
rect -1782 405 -1730 414
rect -1782 371 -1773 405
rect -1773 371 -1739 405
rect -1739 371 -1730 405
rect -1782 362 -1730 371
rect -1718 405 -1666 414
rect -1718 371 -1701 405
rect -1701 371 -1667 405
rect -1667 371 -1666 405
rect -1718 362 -1666 371
rect -1654 405 -1602 414
rect -1590 405 -1538 414
rect -1526 405 -1474 414
rect -1462 405 -1410 414
rect -1398 405 -1346 414
rect -1334 405 -1282 414
rect -1654 371 -1629 405
rect -1629 371 -1602 405
rect -1590 371 -1557 405
rect -1557 371 -1538 405
rect -1526 371 -1523 405
rect -1523 371 -1485 405
rect -1485 371 -1474 405
rect -1462 371 -1451 405
rect -1451 371 -1413 405
rect -1413 371 -1410 405
rect -1398 371 -1379 405
rect -1379 371 -1346 405
rect -1334 371 -1307 405
rect -1307 371 -1282 405
rect -1654 362 -1602 371
rect -1590 362 -1538 371
rect -1526 362 -1474 371
rect -1462 362 -1410 371
rect -1398 362 -1346 371
rect -1334 362 -1282 371
rect -1270 405 -1218 414
rect -1270 371 -1269 405
rect -1269 371 -1235 405
rect -1235 371 -1218 405
rect -1270 362 -1218 371
rect -1206 405 -1154 414
rect -1206 371 -1197 405
rect -1197 371 -1163 405
rect -1163 371 -1154 405
rect -1206 362 -1154 371
rect -1142 405 -1090 414
rect -1142 371 -1125 405
rect -1125 371 -1091 405
rect -1091 371 -1090 405
rect -1142 362 -1090 371
<< metal2 >>
rect -2004 1312 -1970 2036
rect -1568 1925 -957 1944
rect -1568 1869 -1535 1925
rect -1479 1923 -1455 1925
rect -1399 1923 -1375 1925
rect -1319 1923 -1295 1925
rect -1239 1923 -1215 1925
rect -1159 1923 -1135 1925
rect -1079 1923 -1055 1925
rect -1465 1871 -1455 1923
rect -1399 1871 -1389 1923
rect -1145 1871 -1135 1923
rect -1079 1871 -1069 1923
rect -1479 1869 -1455 1871
rect -1399 1869 -1375 1871
rect -1319 1869 -1295 1871
rect -1239 1869 -1215 1871
rect -1159 1869 -1135 1871
rect -1079 1869 -1055 1871
rect -999 1869 -957 1925
rect -1568 1850 -957 1869
rect -1006 1356 -954 1362
rect -1507 1316 -1006 1350
rect -2019 1260 -2013 1312
rect -1961 1260 -1955 1312
rect -1935 1159 -1538 1178
rect -1935 1157 -1884 1159
rect -1828 1157 -1804 1159
rect -1748 1157 -1724 1159
rect -1668 1157 -1644 1159
rect -1588 1157 -1538 1159
rect -1935 1105 -1890 1157
rect -1828 1105 -1826 1157
rect -1646 1105 -1644 1157
rect -1582 1105 -1538 1157
rect -1935 1103 -1884 1105
rect -1828 1103 -1804 1105
rect -1748 1103 -1724 1105
rect -1668 1103 -1644 1105
rect -1588 1103 -1538 1105
rect -1935 1081 -1538 1103
rect -1715 746 -1663 752
rect -1507 737 -1473 1316
rect -1006 1298 -954 1304
rect -1663 703 -1473 737
rect -1715 688 -1663 694
rect -1000 574 -942 583
rect -1000 522 -997 574
rect -945 522 -942 574
rect -1000 513 -942 522
rect -1901 419 -1033 448
rect -1901 363 -1855 419
rect -1799 414 -1775 419
rect -1719 414 -1695 419
rect -1639 414 -1615 419
rect -1559 414 -1535 419
rect -1479 414 -1455 419
rect -1399 414 -1375 419
rect -1319 414 -1295 419
rect -1239 414 -1215 419
rect -1159 414 -1135 419
rect -1901 362 -1846 363
rect -1794 362 -1782 414
rect -1719 363 -1718 414
rect -1538 363 -1535 414
rect -1730 362 -1718 363
rect -1666 362 -1654 363
rect -1602 362 -1590 363
rect -1538 362 -1526 363
rect -1474 362 -1462 414
rect -1399 363 -1398 414
rect -1218 363 -1215 414
rect -1410 362 -1398 363
rect -1346 362 -1334 363
rect -1282 362 -1270 363
rect -1218 362 -1206 363
rect -1154 362 -1142 414
rect -1079 363 -1033 419
rect -1090 362 -1033 363
rect -1901 348 -1033 362
rect -992 243 -949 513
<< via2 >>
rect -1535 1923 -1479 1925
rect -1455 1923 -1399 1925
rect -1375 1923 -1319 1925
rect -1295 1923 -1239 1925
rect -1215 1923 -1159 1925
rect -1135 1923 -1079 1925
rect -1055 1923 -999 1925
rect -1535 1871 -1517 1923
rect -1517 1871 -1479 1923
rect -1455 1871 -1453 1923
rect -1453 1871 -1401 1923
rect -1401 1871 -1399 1923
rect -1375 1871 -1337 1923
rect -1337 1871 -1325 1923
rect -1325 1871 -1319 1923
rect -1295 1871 -1273 1923
rect -1273 1871 -1261 1923
rect -1261 1871 -1239 1923
rect -1215 1871 -1209 1923
rect -1209 1871 -1197 1923
rect -1197 1871 -1159 1923
rect -1135 1871 -1133 1923
rect -1133 1871 -1081 1923
rect -1081 1871 -1079 1923
rect -1055 1871 -1017 1923
rect -1017 1871 -999 1923
rect -1535 1869 -1479 1871
rect -1455 1869 -1399 1871
rect -1375 1869 -1319 1871
rect -1295 1869 -1239 1871
rect -1215 1869 -1159 1871
rect -1135 1869 -1079 1871
rect -1055 1869 -999 1871
rect -1884 1157 -1828 1159
rect -1804 1157 -1748 1159
rect -1724 1157 -1668 1159
rect -1644 1157 -1588 1159
rect -1884 1105 -1838 1157
rect -1838 1105 -1828 1157
rect -1804 1105 -1774 1157
rect -1774 1105 -1762 1157
rect -1762 1105 -1748 1157
rect -1724 1105 -1710 1157
rect -1710 1105 -1698 1157
rect -1698 1105 -1668 1157
rect -1644 1105 -1634 1157
rect -1634 1105 -1588 1157
rect -1884 1103 -1828 1105
rect -1804 1103 -1748 1105
rect -1724 1103 -1668 1105
rect -1644 1103 -1588 1105
rect -1855 414 -1799 419
rect -1775 414 -1719 419
rect -1695 414 -1639 419
rect -1615 414 -1559 419
rect -1535 414 -1479 419
rect -1455 414 -1399 419
rect -1375 414 -1319 419
rect -1295 414 -1239 419
rect -1215 414 -1159 419
rect -1135 414 -1079 419
rect -1855 363 -1846 414
rect -1846 363 -1799 414
rect -1775 363 -1730 414
rect -1730 363 -1719 414
rect -1695 363 -1666 414
rect -1666 363 -1654 414
rect -1654 363 -1639 414
rect -1615 363 -1602 414
rect -1602 363 -1590 414
rect -1590 363 -1559 414
rect -1535 363 -1526 414
rect -1526 363 -1479 414
rect -1455 363 -1410 414
rect -1410 363 -1399 414
rect -1375 363 -1346 414
rect -1346 363 -1334 414
rect -1334 363 -1319 414
rect -1295 363 -1282 414
rect -1282 363 -1270 414
rect -1270 363 -1239 414
rect -1215 363 -1206 414
rect -1206 363 -1159 414
rect -1135 363 -1090 414
rect -1090 363 -1079 414
<< metal3 >>
rect -2042 1944 -1568 1947
rect -957 1944 -883 1947
rect -2042 1925 -883 1944
rect -2042 1869 -1535 1925
rect -1479 1869 -1455 1925
rect -1399 1869 -1375 1925
rect -1319 1869 -1295 1925
rect -1239 1869 -1215 1925
rect -1159 1869 -1135 1925
rect -1079 1869 -1055 1925
rect -999 1869 -883 1925
rect -2042 1847 -883 1869
rect -2042 1159 -883 1180
rect -2042 1103 -1884 1159
rect -1828 1103 -1804 1159
rect -1748 1103 -1724 1159
rect -1668 1103 -1644 1159
rect -1588 1103 -883 1159
rect -2042 1080 -883 1103
rect -2042 419 -883 448
rect -2042 363 -1855 419
rect -1799 363 -1775 419
rect -1719 363 -1695 419
rect -1639 363 -1615 419
rect -1559 363 -1535 419
rect -1479 363 -1455 419
rect -1399 363 -1375 419
rect -1319 363 -1295 419
rect -1239 363 -1215 419
rect -1159 363 -1135 419
rect -1079 363 -883 419
rect -2042 348 -883 363
<< labels >>
rlabel metal3 s -2003 400 -2003 400 4 DVSS
rlabel metal3 s -2030 1133 -2030 1133 4 VCCL
rlabel metal3 s -2025 1905 -2025 1905 4 VCC
rlabel metal2 s -1987 2024 -1987 2024 4 VIN
rlabel metal2 s -969 259 -969 259 4 VOUT
<< end >>
