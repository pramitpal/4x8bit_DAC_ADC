* SPICE3 file created from sample_hold.ext - technology: sky130A

.lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice.tt.red tt
.include /foss/pdks/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

**.subckt sample_hold_tb
x1 CLK VIN VOUT VCC VSS sample_hold
V1 VSS 0 0
.save i(v1)
V2 VCC VSS VCC
.save i(v2)
VMINUS VIN VSS sin(1.65 1.65 freq)
.save i(vminus)
E5 TEMPERAT VSS VOL=' temper '
V4 CLK VSS pulse(0 3.3 0 1p 1p {t/10} {t})
.save i(v4)
**** begin user architecture code



.param freq = 4e4
.param t = {1/(10*freq)}
.param VCC = 3.3

.save all
.tran 50n 100u
**** interactive sim
.control
run
plot vout vin clk/3
.endc

.subckt sample_hold CLK VIN VOUT VCC VSS
X0 m1_900_n309# a_804_n134# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1 m1_1467_624# a_1250_n133# VSS VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.87 ps=7.74 w=1 l=0.5
X2 m1_1068_n250# CLK m1_900_n309# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=5.16 as=0.87 ps=7.74 w=1 l=0.5
X3 VSS a_804_n134# sky130_fd_pr__nfet_g5v0d10v5_SACDK5_5/a_50_n100# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.59 w=1 l=0.5
X4 sky130_fd_pr__nfet_g5v0d10v5_SACDK5_5/a_50_n100# VCC a_1250_n133# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X5 m1_900_n309# a_1250_n133# m1_1068_n250# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0 ps=0 w=1 l=0.5
X6 VSS CLK a_804_n134# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=0.5
X7 VIN a_1250_n133# m1_900_n309# VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=5.16 as=0 ps=0 w=1 l=0.5
X8 m1_1467_624# a_1250_n133# VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X9 a_804_n134# CLK VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=1.16 ps=10.3 w=1 l=0.5
X10 m1_1068_n250# CLK VCC VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X11 VOUT a_1250_n133# VIN VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X12 VIN a_1250_n133# VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X13 VOUT m1_1467_624# VIN VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X14 VIN m1_1467_624# VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X15 VCC a_1250_n133# m1_1059_437# VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X16 m1_1059_437# m1_1068_n250# a_1250_n133# VCC sky130_fd_pr__pfet_g5v0d10v5 ad=0.58 pd=5.16 as=0.29 ps=2.58 w=1 l=0.5
X17 m1_1059_437# m1_900_n309# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X18 m1_1059_437# m1_900_n309# sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X19 VOUT VSS sky130_fd_pr__cap_mim_m3_1 l=10 w=10
X20 VOUT VSS sky130_fd_pr__cap_mim_m3_1 l=10 w=10
C0 m1_1059_437# m1_900_n309# 19.8f
C1 VIN VOUT 1.24f
C2 m1_900_n309# a_1250_n133# 1.04f
C3 m1_1059_437# VCC 1.26f
C4 m1_900_n309# a_804_n134# 1.04f
C5 m1_900_n309# VCC 1.14f
C6 VOUT VSS 22.9f
C7 m1_1059_437# VSS 1.7f 
C8 a_1250_n133# VSS 2.08f 
C9 VCC VSS 7.2f
C10 m1_900_n309# VSS 7.46f 
.ends
