magic
tech sky130A
timestamp 1687456746
<< nwell >>
rect -3191 98 -2877 102
rect -3191 -158 -2531 98
<< pwell >>
rect -2841 -181 -2553 -180
rect -3171 -256 -2553 -181
rect -3171 -257 -2883 -256
rect -3171 -259 -2888 -257
rect -3184 -355 -2888 -259
<< mvnmos >>
rect -3129 -244 -3079 -194
rect -2975 -244 -2925 -194
rect -2799 -243 -2749 -193
rect -2645 -243 -2595 -193
<< mvpmos >>
rect -3129 -125 -3079 -25
rect -2975 -125 -2925 -25
rect -2799 -125 -2749 -25
rect -2645 -125 -2595 -25
<< mvndiff >>
rect -3158 -210 -3129 -194
rect -3158 -227 -3152 -210
rect -3135 -227 -3129 -210
rect -3158 -244 -3129 -227
rect -3079 -210 -3050 -194
rect -3079 -227 -3073 -210
rect -3056 -227 -3050 -210
rect -3079 -244 -3050 -227
rect -3004 -210 -2975 -194
rect -3004 -227 -2998 -210
rect -2981 -227 -2975 -210
rect -3004 -244 -2975 -227
rect -2925 -210 -2896 -194
rect -2925 -227 -2919 -210
rect -2902 -227 -2896 -210
rect -2925 -244 -2896 -227
rect -2828 -209 -2799 -193
rect -2828 -226 -2822 -209
rect -2805 -226 -2799 -209
rect -2828 -243 -2799 -226
rect -2749 -209 -2720 -193
rect -2749 -226 -2743 -209
rect -2726 -226 -2720 -209
rect -2749 -243 -2720 -226
rect -2674 -209 -2645 -193
rect -2674 -226 -2668 -209
rect -2651 -226 -2645 -209
rect -2674 -243 -2645 -226
rect -2595 -209 -2566 -193
rect -2595 -226 -2589 -209
rect -2572 -226 -2566 -209
rect -2595 -243 -2566 -226
<< mvpdiff >>
rect -3158 -32 -3129 -25
rect -3158 -49 -3152 -32
rect -3135 -49 -3129 -32
rect -3158 -66 -3129 -49
rect -3158 -83 -3152 -66
rect -3135 -83 -3129 -66
rect -3158 -100 -3129 -83
rect -3158 -117 -3152 -100
rect -3135 -117 -3129 -100
rect -3158 -125 -3129 -117
rect -3079 -32 -3050 -25
rect -3079 -49 -3073 -32
rect -3056 -49 -3050 -32
rect -3079 -66 -3050 -49
rect -3079 -83 -3073 -66
rect -3056 -83 -3050 -66
rect -3079 -100 -3050 -83
rect -3079 -117 -3073 -100
rect -3056 -117 -3050 -100
rect -3079 -125 -3050 -117
rect -3004 -32 -2975 -25
rect -3004 -49 -2998 -32
rect -2981 -49 -2975 -32
rect -3004 -66 -2975 -49
rect -3004 -83 -2998 -66
rect -2981 -83 -2975 -66
rect -3004 -100 -2975 -83
rect -3004 -117 -2998 -100
rect -2981 -117 -2975 -100
rect -3004 -125 -2975 -117
rect -2925 -32 -2896 -25
rect -2925 -49 -2919 -32
rect -2902 -49 -2896 -32
rect -2925 -66 -2896 -49
rect -2925 -83 -2919 -66
rect -2902 -83 -2896 -66
rect -2925 -100 -2896 -83
rect -2925 -117 -2919 -100
rect -2902 -117 -2896 -100
rect -2925 -125 -2896 -117
rect -2828 -32 -2799 -25
rect -2828 -49 -2822 -32
rect -2805 -49 -2799 -32
rect -2828 -66 -2799 -49
rect -2828 -83 -2822 -66
rect -2805 -83 -2799 -66
rect -2828 -100 -2799 -83
rect -2828 -117 -2822 -100
rect -2805 -117 -2799 -100
rect -2828 -125 -2799 -117
rect -2749 -32 -2720 -25
rect -2749 -49 -2743 -32
rect -2726 -49 -2720 -32
rect -2749 -66 -2720 -49
rect -2749 -83 -2743 -66
rect -2726 -83 -2720 -66
rect -2749 -100 -2720 -83
rect -2749 -117 -2743 -100
rect -2726 -117 -2720 -100
rect -2749 -125 -2720 -117
rect -2674 -32 -2645 -25
rect -2674 -49 -2668 -32
rect -2651 -49 -2645 -32
rect -2674 -66 -2645 -49
rect -2674 -83 -2668 -66
rect -2651 -83 -2645 -66
rect -2674 -100 -2645 -83
rect -2674 -117 -2668 -100
rect -2651 -117 -2645 -100
rect -2674 -125 -2645 -117
rect -2595 -32 -2566 -25
rect -2595 -49 -2589 -32
rect -2572 -49 -2566 -32
rect -2595 -66 -2566 -49
rect -2595 -83 -2589 -66
rect -2572 -83 -2566 -66
rect -2595 -100 -2566 -83
rect -2595 -117 -2589 -100
rect -2572 -117 -2566 -100
rect -2595 -125 -2566 -117
<< mvndiffc >>
rect -3152 -227 -3135 -210
rect -3073 -227 -3056 -210
rect -2998 -227 -2981 -210
rect -2919 -227 -2902 -210
rect -2822 -226 -2805 -209
rect -2743 -226 -2726 -209
rect -2668 -226 -2651 -209
rect -2589 -226 -2572 -209
<< mvpdiffc >>
rect -3152 -49 -3135 -32
rect -3152 -83 -3135 -66
rect -3152 -117 -3135 -100
rect -3073 -49 -3056 -32
rect -3073 -83 -3056 -66
rect -3073 -117 -3056 -100
rect -2998 -49 -2981 -32
rect -2998 -83 -2981 -66
rect -2998 -117 -2981 -100
rect -2919 -49 -2902 -32
rect -2919 -83 -2902 -66
rect -2919 -117 -2902 -100
rect -2822 -49 -2805 -32
rect -2822 -83 -2805 -66
rect -2822 -117 -2805 -100
rect -2743 -49 -2726 -32
rect -2743 -83 -2726 -66
rect -2743 -117 -2726 -100
rect -2668 -49 -2651 -32
rect -2668 -83 -2651 -66
rect -2668 -117 -2651 -100
rect -2589 -49 -2572 -32
rect -2589 -83 -2572 -66
rect -2589 -117 -2572 -100
<< psubdiff >>
rect -3171 -298 -2901 -272
rect -3171 -315 -3146 -298
rect -3129 -315 -3112 -298
rect -3095 -315 -3078 -298
rect -3061 -315 -3044 -298
rect -3027 -315 -3010 -298
rect -2993 -315 -2976 -298
rect -2959 -315 -2942 -298
rect -2925 -315 -2901 -298
rect -3171 -342 -2901 -315
<< mvnsubdiff >>
rect -3156 46 -2896 68
rect -3156 29 -3136 46
rect -3119 29 -3102 46
rect -3085 29 -3068 46
rect -3051 29 -3034 46
rect -3017 29 -3000 46
rect -2983 29 -2966 46
rect -2949 29 -2932 46
rect -2915 29 -2896 46
rect -3156 8 -2896 29
<< psubdiffcont >>
rect -3146 -315 -3129 -298
rect -3112 -315 -3095 -298
rect -3078 -315 -3061 -298
rect -3044 -315 -3027 -298
rect -3010 -315 -2993 -298
rect -2976 -315 -2959 -298
rect -2942 -315 -2925 -298
<< mvnsubdiffcont >>
rect -3136 29 -3119 46
rect -3102 29 -3085 46
rect -3068 29 -3051 46
rect -3034 29 -3017 46
rect -3000 29 -2983 46
rect -2966 29 -2949 46
rect -2932 29 -2915 46
<< poly >>
rect -3129 -25 -3079 -12
rect -2975 -25 -2925 -12
rect -2799 -25 -2749 -12
rect -2645 -25 -2595 -12
rect -3196 -145 -3163 -141
rect -3129 -145 -3079 -125
rect -3196 -146 -3079 -145
rect -3196 -163 -3188 -146
rect -3171 -163 -3079 -146
rect -3196 -165 -3079 -163
rect -3196 -168 -3163 -165
rect -3129 -194 -3079 -165
rect -3039 -150 -3006 -146
rect -2975 -150 -2925 -125
rect -3039 -151 -2925 -150
rect -3039 -168 -3031 -151
rect -3014 -168 -2925 -151
rect -3039 -169 -2925 -168
rect -3039 -173 -3006 -169
rect -2975 -194 -2925 -169
rect -2878 -154 -2845 -149
rect -2799 -154 -2749 -125
rect -2878 -171 -2870 -154
rect -2853 -171 -2749 -154
rect -2709 -145 -2682 -137
rect -2709 -162 -2704 -145
rect -2687 -146 -2682 -145
rect -2645 -146 -2595 -125
rect -2687 -161 -2595 -146
rect -2687 -162 -2682 -161
rect -2709 -170 -2682 -162
rect -2878 -176 -2845 -171
rect -2799 -193 -2749 -171
rect -2645 -193 -2595 -161
rect -3129 -257 -3079 -244
rect -2975 -257 -2925 -244
rect -2799 -256 -2749 -243
rect -2645 -256 -2595 -243
<< polycont >>
rect -3188 -163 -3171 -146
rect -3031 -168 -3014 -151
rect -2870 -171 -2853 -154
rect -2704 -162 -2687 -145
<< locali >>
rect -3161 46 -2891 73
rect -3161 29 -3136 46
rect -3107 29 -3102 46
rect -3071 29 -3068 46
rect -3035 29 -3034 46
rect -3017 29 -3016 46
rect -2983 29 -2980 46
rect -2949 29 -2944 46
rect -2915 29 -2891 46
rect -3161 3 -2891 29
rect -3152 -32 -3135 -23
rect -3152 -66 -3135 -65
rect -3152 -84 -3135 -83
rect -3152 -127 -3135 -117
rect -3073 -32 -3056 -23
rect -3073 -66 -3056 -65
rect -3073 -84 -3056 -83
rect -3073 -127 -3056 -117
rect -2998 -32 -2981 -23
rect -2998 -66 -2981 -65
rect -2998 -84 -2981 -83
rect -2998 -127 -2981 -117
rect -2919 -32 -2902 -23
rect -2919 -66 -2902 -65
rect -2919 -84 -2902 -83
rect -2919 -127 -2902 -117
rect -2822 -32 -2805 -23
rect -2822 -66 -2805 -65
rect -2822 -84 -2805 -83
rect -2822 -127 -2805 -117
rect -2743 -32 -2726 -23
rect -2743 -66 -2726 -65
rect -2743 -84 -2726 -83
rect -2743 -127 -2726 -117
rect -2668 -32 -2651 -23
rect -2668 -66 -2651 -65
rect -2668 -84 -2651 -83
rect -2668 -127 -2651 -117
rect -2589 -32 -2572 -23
rect -2589 -66 -2572 -65
rect -2589 -84 -2572 -83
rect -2589 -127 -2572 -117
rect -3188 -145 -3171 -138
rect -3189 -146 -3169 -145
rect -3189 -163 -3188 -146
rect -3171 -163 -3169 -146
rect -3031 -149 -3014 -143
rect -3189 -164 -3169 -163
rect -3032 -151 -3012 -149
rect -3188 -171 -3171 -164
rect -3032 -168 -3031 -151
rect -3014 -168 -3012 -151
rect -3032 -169 -3012 -168
rect -2870 -153 -2853 -146
rect -2870 -154 -2852 -153
rect -3031 -176 -3014 -169
rect -2853 -171 -2852 -154
rect -2712 -162 -2704 -145
rect -2687 -162 -2679 -145
rect -2870 -179 -2853 -171
rect -3152 -210 -3135 -192
rect -3152 -246 -3135 -227
rect -3073 -210 -3056 -192
rect -3073 -246 -3056 -227
rect -2998 -210 -2981 -192
rect -2998 -246 -2981 -227
rect -2919 -210 -2902 -192
rect -2919 -246 -2902 -227
rect -2822 -209 -2805 -191
rect -2822 -245 -2805 -226
rect -2743 -209 -2726 -191
rect -2743 -245 -2726 -226
rect -2668 -209 -2651 -191
rect -2668 -245 -2651 -226
rect -2589 -209 -2572 -191
rect -2589 -245 -2572 -226
rect -3171 -298 -2901 -272
rect -3171 -315 -3152 -298
rect -3129 -315 -3116 -298
rect -3095 -315 -3080 -298
rect -3061 -315 -3044 -298
rect -3027 -315 -3010 -298
rect -2991 -315 -2976 -298
rect -2955 -315 -2942 -298
rect -2919 -315 -2901 -298
rect -3171 -342 -2901 -315
<< viali >>
rect -3124 29 -3119 46
rect -3119 29 -3107 46
rect -3088 29 -3085 46
rect -3085 29 -3071 46
rect -3052 29 -3051 46
rect -3051 29 -3035 46
rect -3016 29 -3000 46
rect -3000 29 -2999 46
rect -2980 29 -2966 46
rect -2966 29 -2963 46
rect -2944 29 -2932 46
rect -2932 29 -2927 46
rect -3152 -49 -3135 -48
rect -3152 -65 -3135 -49
rect -3152 -100 -3135 -84
rect -3152 -101 -3135 -100
rect -3073 -49 -3056 -48
rect -3073 -65 -3056 -49
rect -3073 -100 -3056 -84
rect -3073 -101 -3056 -100
rect -2998 -49 -2981 -48
rect -2998 -65 -2981 -49
rect -2998 -100 -2981 -84
rect -2998 -101 -2981 -100
rect -2919 -49 -2902 -48
rect -2919 -65 -2902 -49
rect -2919 -100 -2902 -84
rect -2919 -101 -2902 -100
rect -2822 -49 -2805 -48
rect -2822 -65 -2805 -49
rect -2822 -100 -2805 -84
rect -2822 -101 -2805 -100
rect -2743 -49 -2726 -48
rect -2743 -65 -2726 -49
rect -2743 -100 -2726 -84
rect -2743 -101 -2726 -100
rect -2668 -49 -2651 -48
rect -2668 -65 -2651 -49
rect -2668 -100 -2651 -84
rect -2668 -101 -2651 -100
rect -2589 -49 -2572 -48
rect -2589 -65 -2572 -49
rect -2589 -100 -2572 -84
rect -2589 -101 -2572 -100
rect -3188 -163 -3171 -146
rect -3031 -168 -3014 -151
rect -2870 -171 -2853 -154
rect -2704 -162 -2687 -145
rect -3152 -227 -3135 -210
rect -3073 -227 -3056 -210
rect -2998 -227 -2981 -210
rect -2919 -227 -2902 -210
rect -2822 -226 -2805 -209
rect -2743 -226 -2726 -209
rect -2668 -226 -2651 -209
rect -2589 -226 -2572 -209
rect -3152 -315 -3146 -298
rect -3146 -315 -3135 -298
rect -3116 -315 -3112 -298
rect -3112 -315 -3099 -298
rect -3080 -315 -3078 -298
rect -3078 -315 -3063 -298
rect -3044 -315 -3027 -298
rect -3008 -315 -2993 -298
rect -2993 -315 -2991 -298
rect -2972 -315 -2959 -298
rect -2959 -315 -2955 -298
rect -2936 -315 -2925 -298
rect -2925 -315 -2919 -298
<< metal1 >>
rect -3161 51 -2891 73
rect -3161 25 -3135 51
rect -3109 46 -3103 51
rect -3077 46 -3071 51
rect -3045 46 -3039 51
rect -3013 46 -3007 51
rect -2981 46 -2975 51
rect -2949 46 -2943 51
rect -3107 29 -3103 46
rect -2981 29 -2980 46
rect -2949 29 -2944 46
rect -3109 25 -3103 29
rect -3077 25 -3071 29
rect -3045 25 -3039 29
rect -3013 25 -3007 29
rect -2981 25 -2975 29
rect -2949 25 -2943 29
rect -2917 25 -2891 51
rect -3161 3 -2891 25
rect -3152 -25 -3129 3
rect -3155 -48 -3132 -25
rect -3155 -65 -3152 -48
rect -3135 -65 -3132 -48
rect -3155 -84 -3132 -65
rect -3155 -101 -3152 -84
rect -3135 -101 -3132 -84
rect -3155 -125 -3132 -101
rect -3076 -48 -3053 -25
rect -3076 -65 -3073 -48
rect -3056 -65 -3053 -48
rect -3076 -84 -3053 -65
rect -3076 -101 -3073 -84
rect -3056 -101 -3053 -84
rect -3076 -125 -3053 -101
rect -3001 -48 -2978 3
rect -2744 -25 -2724 97
rect -3001 -65 -2998 -48
rect -2981 -65 -2978 -48
rect -3001 -84 -2978 -65
rect -3001 -101 -2998 -84
rect -2981 -101 -2978 -84
rect -3001 -125 -2978 -101
rect -2922 -48 -2899 -25
rect -2922 -65 -2919 -48
rect -2902 -65 -2899 -48
rect -2825 -48 -2802 -25
rect -2825 -61 -2822 -48
rect -2922 -84 -2899 -65
rect -2922 -101 -2919 -84
rect -2902 -101 -2899 -84
rect -2880 -62 -2822 -61
rect -2880 -88 -2877 -62
rect -2851 -65 -2822 -62
rect -2805 -65 -2802 -48
rect -2851 -84 -2802 -65
rect -2851 -88 -2822 -84
rect -2880 -89 -2822 -88
rect -2922 -125 -2899 -101
rect -2825 -101 -2822 -89
rect -2805 -101 -2802 -84
rect -2825 -125 -2802 -101
rect -2746 -48 -2723 -25
rect -2746 -65 -2743 -48
rect -2726 -65 -2723 -48
rect -2671 -48 -2648 -25
rect -2671 -65 -2668 -48
rect -2651 -65 -2648 -48
rect -2746 -84 -2648 -65
rect -2746 -101 -2743 -84
rect -2726 -98 -2668 -84
rect -2726 -101 -2723 -98
rect -2746 -125 -2723 -101
rect -2671 -101 -2668 -98
rect -2651 -101 -2648 -84
rect -2671 -125 -2648 -101
rect -2592 -48 -2569 -25
rect -2592 -65 -2589 -48
rect -2572 -65 -2569 -48
rect -2509 -63 -2494 95
rect -2592 -84 -2569 -65
rect -2592 -101 -2589 -84
rect -2572 -101 -2569 -84
rect -2518 -89 -2515 -63
rect -2489 -89 -2486 -63
rect -2592 -125 -2569 -101
rect -2510 -109 -2494 -89
rect -3192 -145 -3166 -139
rect -3221 -146 -3166 -145
rect -3221 -163 -3188 -146
rect -3171 -163 -3166 -146
rect -3221 -164 -3166 -163
rect -3192 -170 -3166 -164
rect -3074 -149 -3055 -125
rect -3035 -146 -3009 -143
rect -3038 -149 -3035 -146
rect -3074 -169 -3035 -149
rect -3074 -194 -3055 -169
rect -3038 -172 -3035 -169
rect -3009 -172 -3006 -146
rect -2920 -153 -2900 -125
rect -2873 -153 -2849 -147
rect -2920 -154 -2849 -153
rect -2920 -170 -2870 -154
rect -3035 -175 -3009 -172
rect -2920 -194 -2900 -170
rect -2873 -171 -2870 -170
rect -2853 -171 -2849 -154
rect -2873 -177 -2849 -171
rect -3155 -210 -3132 -194
rect -3155 -227 -3152 -210
rect -3135 -227 -3132 -210
rect -3155 -244 -3132 -227
rect -3076 -210 -3053 -194
rect -3076 -227 -3073 -210
rect -3056 -227 -3053 -210
rect -3001 -210 -2978 -194
rect -3001 -225 -2998 -210
rect -3076 -244 -3053 -227
rect -3002 -227 -2998 -225
rect -2981 -227 -2978 -210
rect -3155 -272 -3133 -244
rect -3002 -272 -2978 -227
rect -2922 -210 -2899 -194
rect -2922 -227 -2919 -210
rect -2902 -227 -2899 -210
rect -2922 -244 -2899 -227
rect -3171 -294 -2901 -272
rect -3171 -298 -3145 -294
rect -3119 -298 -3113 -294
rect -3171 -315 -3152 -298
rect -3119 -315 -3116 -298
rect -3171 -320 -3145 -315
rect -3119 -320 -3113 -315
rect -3087 -320 -3081 -294
rect -3055 -320 -3049 -294
rect -3023 -320 -3017 -294
rect -2991 -320 -2985 -294
rect -2959 -298 -2953 -294
rect -2927 -298 -2901 -294
rect -2955 -315 -2953 -298
rect -2919 -315 -2901 -298
rect -2959 -320 -2953 -315
rect -2927 -320 -2901 -315
rect -3171 -342 -2901 -320
rect -2870 -372 -2850 -177
rect -2744 -193 -2724 -125
rect -2709 -140 -2683 -137
rect -2710 -165 -2709 -142
rect -2683 -165 -2681 -142
rect -2585 -163 -2571 -125
rect -2709 -169 -2683 -166
rect -2585 -177 -2534 -163
rect -2825 -209 -2802 -193
rect -2825 -226 -2822 -209
rect -2805 -226 -2802 -209
rect -2825 -243 -2802 -226
rect -2746 -203 -2723 -193
rect -2671 -203 -2648 -193
rect -2592 -203 -2569 -193
rect -2746 -209 -2648 -203
rect -2746 -226 -2743 -209
rect -2726 -226 -2668 -209
rect -2651 -226 -2648 -209
rect -2746 -236 -2648 -226
rect -2595 -229 -2592 -203
rect -2566 -229 -2563 -203
rect -2746 -243 -2723 -236
rect -2671 -243 -2648 -236
rect -2592 -243 -2569 -229
rect -2822 -318 -2808 -243
rect -2744 -265 -2724 -243
rect -2747 -268 -2721 -265
rect -2747 -297 -2721 -294
rect -2548 -318 -2534 -177
rect -2510 -202 -2495 -109
rect -2518 -228 -2515 -202
rect -2489 -228 -2486 -202
rect -2822 -332 -2534 -318
rect -3235 -391 -2850 -372
rect -2548 -379 -2534 -332
<< via1 >>
rect -3135 46 -3109 51
rect -3103 46 -3077 51
rect -3071 46 -3045 51
rect -3039 46 -3013 51
rect -3007 46 -2981 51
rect -2975 46 -2949 51
rect -2943 46 -2917 51
rect -3135 29 -3124 46
rect -3124 29 -3109 46
rect -3103 29 -3088 46
rect -3088 29 -3077 46
rect -3071 29 -3052 46
rect -3052 29 -3045 46
rect -3039 29 -3035 46
rect -3035 29 -3016 46
rect -3016 29 -3013 46
rect -3007 29 -2999 46
rect -2999 29 -2981 46
rect -2975 29 -2963 46
rect -2963 29 -2949 46
rect -2943 29 -2927 46
rect -2927 29 -2917 46
rect -3135 25 -3109 29
rect -3103 25 -3077 29
rect -3071 25 -3045 29
rect -3039 25 -3013 29
rect -3007 25 -2981 29
rect -2975 25 -2949 29
rect -2943 25 -2917 29
rect -2877 -88 -2851 -62
rect -2515 -89 -2489 -63
rect -3035 -151 -3009 -146
rect -3035 -168 -3031 -151
rect -3031 -168 -3014 -151
rect -3014 -168 -3009 -151
rect -3035 -172 -3009 -168
rect -3145 -298 -3119 -294
rect -3113 -298 -3087 -294
rect -3145 -315 -3135 -298
rect -3135 -315 -3119 -298
rect -3113 -315 -3099 -298
rect -3099 -315 -3087 -298
rect -3145 -320 -3119 -315
rect -3113 -320 -3087 -315
rect -3081 -298 -3055 -294
rect -3081 -315 -3080 -298
rect -3080 -315 -3063 -298
rect -3063 -315 -3055 -298
rect -3081 -320 -3055 -315
rect -3049 -298 -3023 -294
rect -3049 -315 -3044 -298
rect -3044 -315 -3027 -298
rect -3027 -315 -3023 -298
rect -3049 -320 -3023 -315
rect -3017 -298 -2991 -294
rect -3017 -315 -3008 -298
rect -3008 -315 -2991 -298
rect -3017 -320 -2991 -315
rect -2985 -298 -2959 -294
rect -2953 -298 -2927 -294
rect -2985 -315 -2972 -298
rect -2972 -315 -2959 -298
rect -2953 -315 -2936 -298
rect -2936 -315 -2927 -298
rect -2985 -320 -2959 -315
rect -2953 -320 -2927 -315
rect -2709 -145 -2683 -140
rect -2709 -162 -2704 -145
rect -2704 -162 -2687 -145
rect -2687 -162 -2683 -145
rect -2709 -166 -2683 -162
rect -2592 -209 -2566 -203
rect -2592 -226 -2589 -209
rect -2589 -226 -2572 -209
rect -2572 -226 -2566 -209
rect -2592 -229 -2566 -226
rect -2747 -294 -2721 -268
rect -2515 -228 -2489 -202
<< metal2 >>
rect -3441 -190 -3420 118
rect -3401 -190 -3380 118
rect -3361 -190 -3340 118
rect -3321 -190 -3300 118
rect -3281 -190 -3260 118
rect -3241 -190 -3220 118
rect -3161 52 -2891 73
rect -3161 24 -3140 52
rect -3112 51 -3100 52
rect -3072 51 -3060 52
rect -3032 51 -3020 52
rect -2992 51 -2980 52
rect -2952 51 -2940 52
rect -3109 25 -3103 51
rect -3072 25 -3071 51
rect -2981 25 -2980 51
rect -2949 25 -2943 51
rect -3112 24 -3100 25
rect -3072 24 -3060 25
rect -3032 24 -3020 25
rect -2992 24 -2980 25
rect -2952 24 -2940 25
rect -2912 24 -2891 52
rect -3161 3 -2891 24
rect -2877 -61 -2850 -58
rect -2515 -61 -2489 -60
rect -2877 -62 -2481 -61
rect -2851 -63 -2481 -62
rect -2851 -88 -2515 -63
rect -2877 -89 -2515 -88
rect -2489 -89 -2481 -63
rect -2877 -92 -2850 -89
rect -2515 -92 -2489 -89
rect -3035 -146 -3009 -143
rect -2712 -166 -2709 -140
rect -2683 -166 -2680 -140
rect -3035 -175 -3009 -172
rect -3033 -198 -3014 -175
rect -2704 -198 -2687 -166
rect -3033 -218 -2686 -198
rect -2592 -203 -2566 -200
rect -2515 -202 -2489 -199
rect -2566 -223 -2515 -208
rect -3441 -495 -3420 -230
rect -3401 -495 -3380 -230
rect -3361 -495 -3340 -230
rect -3321 -495 -3300 -230
rect -3281 -495 -3260 -230
rect -3241 -495 -3220 -230
rect -2592 -232 -2566 -229
rect -2515 -231 -2489 -228
rect -3171 -293 -2901 -272
rect -3171 -321 -3150 -293
rect -3122 -294 -3110 -293
rect -3082 -294 -3070 -293
rect -3042 -294 -3030 -293
rect -3002 -294 -2990 -293
rect -2962 -294 -2950 -293
rect -3119 -320 -3113 -294
rect -3082 -320 -3081 -294
rect -2991 -320 -2990 -294
rect -2959 -320 -2953 -294
rect -3122 -321 -3110 -320
rect -3082 -321 -3070 -320
rect -3042 -321 -3030 -320
rect -3002 -321 -2990 -320
rect -2962 -321 -2950 -320
rect -2922 -321 -2901 -293
rect -2750 -294 -2747 -268
rect -2721 -294 -2718 -268
rect -3171 -342 -2901 -321
rect -2743 -376 -2724 -294
<< via2 >>
rect -3140 51 -3112 52
rect -3100 51 -3072 52
rect -3060 51 -3032 52
rect -3020 51 -2992 52
rect -2980 51 -2952 52
rect -2940 51 -2912 52
rect -3140 25 -3135 51
rect -3135 25 -3112 51
rect -3100 25 -3077 51
rect -3077 25 -3072 51
rect -3060 25 -3045 51
rect -3045 25 -3039 51
rect -3039 25 -3032 51
rect -3020 25 -3013 51
rect -3013 25 -3007 51
rect -3007 25 -2992 51
rect -2980 25 -2975 51
rect -2975 25 -2952 51
rect -2940 25 -2917 51
rect -2917 25 -2912 51
rect -3140 24 -3112 25
rect -3100 24 -3072 25
rect -3060 24 -3032 25
rect -3020 24 -2992 25
rect -2980 24 -2952 25
rect -2940 24 -2912 25
rect -3150 -294 -3122 -293
rect -3110 -294 -3082 -293
rect -3070 -294 -3042 -293
rect -3030 -294 -3002 -293
rect -2990 -294 -2962 -293
rect -2950 -294 -2922 -293
rect -3150 -320 -3145 -294
rect -3145 -320 -3122 -294
rect -3110 -320 -3087 -294
rect -3087 -320 -3082 -294
rect -3070 -320 -3055 -294
rect -3055 -320 -3049 -294
rect -3049 -320 -3042 -294
rect -3030 -320 -3023 -294
rect -3023 -320 -3017 -294
rect -3017 -320 -3002 -294
rect -2990 -320 -2985 -294
rect -2985 -320 -2962 -294
rect -2950 -320 -2927 -294
rect -2927 -320 -2922 -294
rect -3150 -321 -3122 -320
rect -3110 -321 -3082 -320
rect -3070 -321 -3042 -320
rect -3030 -321 -3002 -320
rect -2990 -321 -2962 -320
rect -2950 -321 -2922 -320
<< metal3 >>
rect -3466 52 -2461 73
rect -3466 24 -3140 52
rect -3112 24 -3100 52
rect -3072 24 -3060 52
rect -3032 24 -3020 52
rect -2992 24 -2980 52
rect -2952 24 -2940 52
rect -2912 24 -2461 52
rect -3466 3 -2461 24
rect -3466 -293 -2461 -272
rect -3466 -321 -3150 -293
rect -3122 -321 -3110 -293
rect -3082 -321 -3070 -293
rect -3042 -321 -3030 -293
rect -3002 -321 -2990 -293
rect -2962 -321 -2950 -293
rect -2922 -321 -2461 -293
rect -3466 -342 -2461 -321
<< labels >>
flabel metal1 s -3221 -164 -3211 -145 7 FreeSans 300 0 0 0 DX
port 1 w
flabel metal1 s -3235 -391 -3221 -372 7 FreeSans 300 0 0 0 DX_BUF
port 2 w
flabel metal3 s -2476 3 -2461 73 3 FreeSans 300 0 0 0 VCC
port 3 e
flabel metal3 s -2476 -342 -2461 -272 3 FreeSans 300 0 0 0 VSS
port 4 e
flabel metal3 s -3466 -342 -3451 -272 7 FreeSans 300 0 0 0 VSS
port 4 w
flabel metal3 s -3466 3 -3451 73 7 FreeSans 300 0 0 0 VCC
port 3 w
flabel metal2 s -3431 111 -3431 111 1 FreeSans 200 0 0 0 D2
port 5 n
flabel metal2 s -3391 113 -3391 113 1 FreeSans 200 0 0 0 D3
port 6 n
flabel metal2 s -3350 113 -3350 113 1 FreeSans 200 0 0 0 D4
port 7 n
flabel metal2 s -3310 114 -3310 114 1 FreeSans 200 0 0 0 D5
port 8 n
flabel metal2 s -3271 114 -3271 114 1 FreeSans 200 0 0 0 D6
port 9 n
flabel metal2 s -3231 113 -3231 113 1 FreeSans 200 0 0 0 D7
port 10 n
flabel metal1 s -2744 85 -2724 97 3 FreeSans 300 0 0 0 VOUT
port 11 e
flabel metal2 s -2743 -376 -2724 -364 7 FreeSans 300 0 0 0 VOUT
port 11 w
flabel metal1 s -2548 -379 -2534 -367 3 FreeSans 300 0 0 0 VREFH
port 12 e
flabel metal1 s -2509 83 -2494 93 3 FreeSans 300 0 0 0 VREFL
port 13 e
<< end >>
