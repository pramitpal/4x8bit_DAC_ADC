** sch_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/All_schematic/8_bit_dac.sch
.subckt 8_bit_dac D0 D1 D2 D7 VREFH VREFL D0_BUF D1_BUF D2_BUF D7_BUF VOUT VCC VSS D3 D3_BUF D4
+ D4_BUF D5 D5_BUF D6_BUF D6
*.PININFO D0:I D1:I D2:I D7:I VREFH:I VREFL:I D0_BUF:O D1_BUF:O D2_BUF:O D7_BUF:O VOUT:O VCC:B VSS:B
*+ D3:I D3_BUF:O D4:I D4_BUF:O D5:I D5_BUF:O D6_BUF:O D6:I
x1 VCC VREFH VSS D0_BUF D1_BUF D2_BUF D3_BUF D4_BUF D5_BUF BUF6 D6_BUF VINH BUF0 BUF1 BUF2 BUF3 BUF4
+ BUF5 VINT 7_bit_dac
x2 VCC VINT VSS BUF0 BUF1 BUF2 BUF3 BUF4 BUF5 D6 BUF6 VINL D0 D1 D2 D3 D4 D5 VREFL 7_bit_dac
x3 VCC D7 D7_BUF VSS VINH VOUT VINL switch_n_3v3
.ends

* expanding   symbol:  /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/All_schematic/7_bit_dac.sym
*+ # of pins=19
** sym_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/All_schematic/7_bit_dac.sym
** sch_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/All_schematic/7_bit_dac.sch
.subckt 7_bit_dac VCC VREFH VSS D0_BUF D1_BUF D2_BUF D3_BUF D4_BUF D5_BUF D6 D6_BUF VOUT D0 D1 D2 D3
+ D4 D5 VREFL
*.PININFO D0:I D1:I D2:I D6:I VREFH:I VREFL:I D0_BUF:O D1_BUF:O D2_BUF:O D6_BUF:O VOUT:O VCC:B VSS:B
*+ D3:I D3_BUF:O D4:I D4_BUF:O D5:I D5_BUF:O
x1 VCC VREFH VSS D0_BUF D1_BUF D2_BUF D3_BUF D4_BUF BUF5 D5_BUF VINH BUF0 BUF1 BUF2 BUF3 BUF4 VINT
+ 6_bit_dac
x2 VCC VINT VSS BUF0 BUF1 BUF2 BUF3 BUF4 D5 BUF5 VINL D0 D1 D2 D3 D4 VREFL 6_bit_dac
x3 VCC D6 D6_BUF VSS VINH VOUT VINL switch_n_3v3
.ends


* expanding   symbol:
*+  /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/All_schematic/switch_n_3v3.sym # of pins=7
** sym_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/All_schematic/switch_n_3v3.sym
** sch_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/All_schematic/switch_n_3v3.sch
.subckt switch_n_3v3 VCC DX DX_BUF VSS VREFH VOUT VREFL
*.PININFO VCC:B VSS:B DX_BUF:O VOUT:O DX:I VREFH:I VREFL:I
XM1 net1 DX VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM2 net1 DX VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM3 DX_BUF net1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM4 DX_BUF net1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM5 VOUT net1 VREFL VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM6 VOUT net1 VREFH VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM7 VREFL DX_BUF VOUT VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM8 VREFH DX_BUF VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
.ends


* expanding   symbol:  /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/All_schematic/6_bit_dac.sym
*+ # of pins=17
** sym_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/All_schematic/6_bit_dac.sym
** sch_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/All_schematic/6_bit_dac.sch
.subckt 6_bit_dac VCC VREFH VSS D0_BUF D1_BUF D2_BUF D3_BUF D4_BUF D5 D5_BUF VOUT D0 D1 D2 D3 D4
+ VREFL
*.PININFO D0:I D1:I D2:I D5:I VREFH:I VREFL:I D0_BUF:O D1_BUF:O D2_BUF:O D5_BUF:O VOUT:O VCC:B VSS:B
*+ D3:I D3_BUF:O D4:I D4_BUF:O
X1 VCC VREFH VSS D0_BUF D1_BUF D2_BUF D3_BUF BUF4 D4_BUF VINH BUF0 BUF1 BUF2 BUF3 VINT 5_bit_dac
X2 VCC VINT VSS BUF0 BUF1 BUF2 BUF3 D4 BUF4 VINL D0 D1 D2 D3 VREFL 5_bit_dac
x3 VCC D5 D5_BUF VSS VINH VOUT VINL switch_n_3v3
.ends


* expanding   symbol:  /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/All_schematic/5_bit_dac.sym
*+ # of pins=15
** sym_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/All_schematic/5_bit_dac.sym
** sch_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/All_schematic/5_bit_dac.sch
.subckt 5_bit_dac VCC VREFH VSS D0_BUF D1_BUF D2_BUF D3_BUF D4 D4_BUF VOUT D0 D1 D2 D3 VREFL
*.PININFO D0:I D1:I D2:I D4:I VREFH:I VREFL:I D0_BUF:O D1_BUF:O D2_BUF:O D4_BUF:O VOUT:O VCC:B VSS:B
*+ D3:I D3_BUF:O
X1 VCC VREFH VSS D0_BUF D1_BUF D2_BUF BUF3 D3_BUF VINH BUF0 BUF1 BUF2 VINT 4_bit_dac
X2 VCC VINT VSS BUF0 BUF1 BUF2 D3 BUF3 VINL D0 D1 D2 VREFL 4_bit_dac
x3 VCC D4 D4_BUF VSS VINH VOUT VINL switch_n_3v3
.ends


* expanding   symbol:  /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/All_schematic/4_bit_dac.sym
*+ # of pins=13
** sym_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/All_schematic/4_bit_dac.sym
** sch_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/All_schematic/4_bit_dac.sch
.subckt 4_bit_dac VCC VREFH VSS D0_BUF D1_BUF D2_BUF D3 D3_BUF VOUT D0 D1 D2 VREFL
*.PININFO D0:I D1:I D2:I D3:I VREFH:I VREFL:I D0_BUF:O D1_BUF:O D2_BUF:O D3_BUF:O VOUT:O VCC:B VSS:B
X1 VCC VSS VREFH D0_BUF D1_BUF BUF2 D2_BUF VINH BUF0 BUF1 VINT 3_bit_dac
X2 VCC VSS VINT BUF0 BUF1 D2 BUF2 VINL D0 D1 VREFL 3_bit_dac
x3 VCC D3 D3_BUF VSS VINH VOUT VINL switch_n_3v3
.ends


* expanding   symbol:  /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/All_schematic/3_bit_dac.sym
*+ # of pins=11
** sym_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/All_schematic/3_bit_dac.sym
** sch_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/All_schematic/3_bit_dac.sch
.subckt 3_bit_dac VCC VSS VREFH D0_BUF D1_BUF D2 D2_BUF VOUT D0 D1 VREFL
*.PININFO D2:I D0_BUF:O D2_BUF:O VOUT:O VREFH:I VCC:B VSS:B D1_BUF:O D1:I VREFL:I D0:I
x2 VCC D2 D2_BUF VSS VINH VOUT VINL switch_n_3v3
X1 VCC VSS BUF0 BUF1 VREFH D0_BUF D1_BUF VINT VINH 2_bit_dac
X3 VCC VSS D0 D1 VINT BUF0 BUF1 VREFL VINL 2_bit_dac
.ends


* expanding   symbol:  /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/All_schematic/2_bit_dac.sym
*+ # of pins=9
** sym_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/All_schematic/2_bit_dac.sym
** sch_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/All_schematic/2_bit_dac.sch
.subckt 2_bit_dac VCC VSS D0 D1 VREFH D0_BUF D1_BUF VREFL VOUT
*.PININFO D1:I D0:I D0_BUF:O D1_BUF:O VOUT:O VREFL:I VREFH:I VCC:B VSS:B
x1 VCC D0_BUF D0 VREFH VSS VINL VINH VREFL switch2n_3v3
x2 VCC D1 D1_BUF VSS VINH VOUT VINL switch_n_3v3
.ends


* expanding   symbol:
*+  /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/All_schematic/switch2n_3v3.sym # of pins=8
** sym_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/All_schematic/switch2n_3v3.sym
** sch_path: /foss/designs/8_bit_dac/All_layouts/Layout_v2/lvs/All_schematic/switch2n_3v3.sch
.subckt switch2n_3v3 VCC DX_BUF DX VREFH VSS VOUTL VOUTH VREFL
*.PININFO VCC:B VSS:B VOUTL:O DX:I VOUTH:O DX_BUF:O VREFH:I VREFL:I
XM1 net1 DX VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM2 net1 DX VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM3 DX_BUF net1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM4 DX_BUF net1 VCC VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM5 VOUTL net1 VREFL VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM6 VOUTL net1 net2 VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM7 VREFL DX_BUF VOUTL VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM8 net2 DX_BUF VOUTL VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM9 VOUTH net1 net3 VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM10 VOUTH net1 net4 VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM11 net3 DX_BUF VOUTH VCC sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM12 net4 DX_BUF VOUTH VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XR1 net3 net4 VSS sky130_fd_pr__res_generic_nd__hv W=1 L=1 mult=1 m=1
XR2 net2 net3 VSS sky130_fd_pr__res_generic_nd__hv W=1 L=1 mult=1 m=1
XR3 VREFL net2 VSS sky130_fd_pr__res_generic_nd__hv W=1 L=1 mult=1 m=1
XR4 net4 VREFH VSS sky130_fd_pr__res_generic_nd__hv W=1 L=1 mult=1 m=1
.ends

.end
