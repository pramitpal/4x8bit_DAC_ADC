magic
tech sky130A
magscale 1 2
timestamp 1686569624
<< locali >>
rect 3 78948 476 79088
<< viali >>
rect -137 78948 3 79088
rect 0 0 140 140
<< metal1 >>
rect -153 79094 22 79108
rect -153 78942 -143 79094
rect 9 78942 22 79094
rect -153 78932 22 78942
rect -6 146 146 152
rect -12 -6 -6 146
rect 134 140 146 146
rect 140 0 146 140
rect 134 -6 146 0
rect -6 -12 146 -6
<< via1 >>
rect -143 79088 9 79094
rect -143 78948 -137 79088
rect -137 78948 3 79088
rect 3 78948 9 79088
rect -143 78942 9 78948
rect -6 140 134 146
rect -6 0 0 140
rect 0 0 134 140
rect -6 -6 134 0
<< metal2 >>
rect 745 85774 779 86800
rect 848 85794 882 86800
rect 946 85794 980 86800
rect 1050 85794 1084 86800
rect 1158 85793 1192 86800
rect 1258 85785 1292 86800
rect 1366 85794 1400 86800
rect 1478 85782 1512 86800
rect 9265 85699 9373 86800
rect 11346 85794 11380 86800
rect 11449 85794 11483 86800
rect 11547 85794 11581 86800
rect 11651 85794 11685 86800
rect 11759 85786 11793 86800
rect 11859 85794 11893 86800
rect 11967 85794 12001 86800
rect 12079 85794 12113 86800
rect 19866 85716 19974 86800
rect 21947 85794 21981 86800
rect 22050 85788 22084 86800
rect 22148 85794 22182 86800
rect 22252 85788 22286 86800
rect 22360 85794 22394 86800
rect 22460 85794 22494 86800
rect 22568 85786 22602 86800
rect 22680 85794 22714 86800
rect 30467 85720 30575 86800
rect 32548 85794 32582 86800
rect 32651 85794 32685 86800
rect 32749 85794 32783 86800
rect 32853 85794 32887 86800
rect 32961 85794 32995 86800
rect 33061 85782 33095 86800
rect 33169 85794 33203 86800
rect 33281 85794 33315 86800
rect 41068 85720 41176 86800
rect -153 79094 22 79108
rect -153 79088 -143 79094
rect -800 78948 -143 79088
rect -153 78942 -143 78948
rect 9 78942 22 79094
rect -153 78932 22 78942
rect -6 146 134 152
rect -800 0 -6 140
rect -6 -12 134 -6
use 4x8bit_tx_buffer  4x8bit_tx_buffer_0
timestamp 1686560844
transform 1 0 0 0 1 0
box 0 0 42404 85828
<< labels >>
rlabel metal2 745 86000 779 86800 1 D00
port 1 n signal input
rlabel metal2 848 86000 882 86800 1 D01
port 2 n signal input
rlabel metal2 946 86000 980 86800 1 D02
port 3 n signal input
rlabel metal2 1050 86000 1084 86800 1 D03
port 4 n signal input
rlabel metal2 1158 86000 1192 86800 1 D04
port 5 n signal input
rlabel metal2 1258 86000 1292 86800 1 D05
port 6 n signal input
rlabel metal2 1366 86000 1400 86800 1 D06
port 7 n signal input
rlabel metal2 1478 86000 1512 86800 1 D07
port 8 n signal input
rlabel metal2 11346 86000 11380 86800 1 D10
port 9 n signal input
rlabel metal2 11449 86000 11483 86800 1 D11
port 10 n signal input
rlabel metal2 11547 86000 11581 86800 1 D12
port 11 n signal input
rlabel metal2 11651 86000 11685 86800 1 D13
port 12 n signal input
rlabel metal2 11759 86000 11793 86800 1 D14
port 13 n signal input
rlabel metal2 11859 86000 11893 86800 1 D15
port 14 n signal input
rlabel metal2 11967 86000 12001 86800 1 D16
port 15 n signal input
rlabel metal2 12079 86000 12113 86800 1 D17
port 16 n signal input
rlabel metal2 21947 86000 21981 86800 1 D20
port 17 n signal input
rlabel metal2 22050 86000 22084 86800 1 D21
port 18 n signal input
rlabel metal2 22148 86000 22182 86800 1 D22
port 19 n signal input
rlabel metal2 22252 86000 22286 86800 1 D23
port 20 n signal input
rlabel metal2 22360 86000 22394 86800 1 D24
port 21 n signal input
rlabel metal2 22460 86000 22494 86800 1 D25
port 22 n signal input
rlabel metal2 22568 86000 22602 86800 1 D26
port 23 n signal input
rlabel metal2 22680 86000 22714 86800 1 D27
port 24 n signal input
rlabel metal2 32548 86000 32582 86800 1 D30
port 25 n signal input
rlabel metal2 32651 86000 32685 86800 1 D31
port 26 n signal input
rlabel metal2 32749 86000 32783 86800 1 D32
port 27 n signal input
rlabel metal2 32853 86000 32887 86800 1 D33
port 28 n signal input
rlabel metal2 32961 86000 32995 86800 1 D34
port 29 n signal input
rlabel metal2 33061 86000 33095 86800 1 D35
port 30 n signal input
rlabel metal2 33169 86000 33203 86800 1 D36
port 31 n signal input
rlabel metal2 33281 86000 33315 86800 1 D37
port 32 n signal input
rlabel metal2 9265 86000 9373 86800 1 VOUT0
port 33 n signal output
rlabel metal2 19866 86000 19974 86800 1 VOUT1
port 34 n signal output
rlabel metal2 30467 86000 30575 86800 1 VOUT2
port 35 n signal output
rlabel metal2 41068 86000 41176 86800 1 VOUT3
port 36 n signal output
rlabel metal2 -800 78948 -200 79088 7 VREFL
port 37 w signal input
rlabel metal2 -800 0 -200 140 7 VREFH
port 38 w signal input
<< properties >>
string FIXED_BBOX -500 -500 43000 86390
<< end >>
