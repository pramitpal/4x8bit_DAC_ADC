magic
tech sky130A
magscale 1 2
timestamp 1686021299
<< metal1 >>
rect 6968 6086 6974 6138
rect 7026 6086 7032 6138
rect 6985 5977 7015 6086
rect 5273 5481 5279 5533
rect 5331 5526 5337 5533
rect 5331 5487 5601 5526
rect 5331 5481 5337 5487
rect 5273 5027 5279 5079
rect 5331 5072 5337 5079
rect 5331 5033 5584 5072
rect 5331 5027 5337 5033
rect 6908 4964 6936 5094
rect 6908 4936 7234 4964
rect 7206 4678 7234 4936
rect 7194 4672 7246 4678
rect 7194 4614 7246 4620
<< via1 >>
rect 6974 6086 7026 6138
rect 5279 5481 5331 5533
rect 5279 5027 5331 5079
rect 7194 4620 7246 4672
<< metal2 >>
rect 274 9499 329 9822
rect 378 9521 433 9824
rect 3564 9684 3605 9824
rect 5122 9706 5163 9824
rect 5202 9694 5243 9824
rect 5282 9698 5323 9824
rect 7111 8429 7241 8468
rect 6974 6138 7026 6144
rect 7202 6127 7241 8429
rect 7026 6097 7241 6127
rect 6974 6080 7026 6086
rect 42 4542 110 6042
rect 5279 5533 5331 5539
rect 144 3836 212 5382
rect 5122 5322 5163 5477
rect 5202 5332 5243 5477
rect 5279 5475 5331 5481
rect 5362 5316 5403 5477
rect 5442 5328 5483 5477
rect 5522 5296 5563 5477
rect 5279 5079 5331 5085
rect 6517 5063 7193 5102
rect 5279 5021 5331 5027
rect 7188 4620 7194 4672
rect 7246 4620 7252 4672
rect 7196 3556 7235 4620
rect 7103 3517 7235 3556
rect 5122 1272 5163 1450
rect 5202 1272 5243 1418
rect 5282 1272 5323 1410
rect 277 0 332 213
rect 378 0 433 373
rect 3564 0 3605 104
use 4_bit_dac  4_bit_dac_0
array 0 0 7165 0 1 4912
timestamp 1686021299
transform 1 0 0 0 1 0
box 0 0 7329 4912
use switch_n_3v3  switch_n_3v3_0
timestamp 1686019770
transform 1 0 12004 0 1 5816
box -6932 -991 -4922 237
<< labels >>
rlabel metal2 72 4824 72 4824 7 VCC
rlabel metal2 170 4830 170 4830 7 VSS
rlabel metal2 308 9780 308 9780 7 D0
rlabel metal2 416 9768 416 9768 7 VREFL
rlabel metal2 312 44 312 44 7 D0_BUF
rlabel metal2 402 34 402 34 7 VREFH
rlabel metal2 3574 22 3574 22 7 D1_BUF
rlabel metal2 3586 9790 3586 9790 7 D1
rlabel metal2 5150 9800 5150 9800 7 D2
rlabel metal2 5222 9798 5222 9798 7 D3
rlabel metal2 5302 9806 5302 9806 7 D4
rlabel metal2 5152 1296 5152 1296 3 D2_BUF
rlabel metal2 5220 1306 5220 1306 3 D3_BUF
rlabel metal2 5294 1284 5294 1284 3 D4_BUF
rlabel metal2 7176 5084 7176 5084 3 VOUT
<< end >>
