* SPICE3 file created from 6_bit_dac.ext - technology: sky130A

.subckt x6_bit_dac D0 VREFL D1 D2 D3 D4 D5 D0_BUF VREFH D1_BUF D2_BUF D3_BUF D4_BUF
+ D5_BUF VOUT VCC VSS
X0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H D0_BUF.t2 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VCC.t129 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t29 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X2 5_bit_dac_0[1].4_bit_dac_0[0].VOUT 5_bit_dac_0[1].switch_n_3v3_0.DX_ 5_bit_dac_0[1].VOUT VCC.t210 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X3 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 a_1556_7774# VSS.t231 VSS.t230 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X4 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X5 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X6 5_bit_dac_0[0].4_bit_dac_0[0].D0 a_1556_5318# VCC.t170 VCC.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X7 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_2862# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L VCC.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X8 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X9 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X10 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_6546# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X11 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_1634# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH VCC.t220 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X12 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_4090# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH VCC.t110 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X13 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VSS.t223 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X14 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VREFH VSS.t29 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X15 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 VSS.t126 VSS.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X16 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].VREFH VSS.t29 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X17 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 VCC.t243 VCC.t242 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X18 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VCC.t101 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X19 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X20 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X21 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t174 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X22 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 a_1556_9002# VCC.t114 VCC.t113 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X23 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VCC.t136 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X24 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X25 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].VOUT VSS.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X26 a_1556_11458# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 VCC.t275 VCC.t274 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X27 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X28 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 VSS.t266 VSS.t265 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X29 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS.t123 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X30 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 VCC.t207 VCC.t206 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X31 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_4090# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X32 a_1556_17598# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 VCC.t285 VCC.t284 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X33 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[0].switch_n_3v3_0.D2 VCC.t83 VCC.t82 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X34 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].VOUT D2_BUF.t2 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X35 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X36 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_7774# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH VCC.t225 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X37 5_bit_dac_0[1].VOUT switch_n_3v3_0.D4.t2 5_bit_dac_0[1].4_bit_dac_0[0].VOUT VSS.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X38 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VCC.t106 VCC.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X39 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t93 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X40 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t275 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X41 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 VCC.t64 VCC.t63 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X42 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_11458# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t279 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X43 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VCC.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X44 switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ VSS.t296 VSS.t295 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X45 a_1556_10230# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 VSS.t107 VSS.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X46 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t2 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X47 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS.t240 VSS.t239 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X48 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_12686# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH VCC.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X49 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.DX_ VSS.t310 VSS.t309 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X50 VOUT.t0 D5_BUF.t2 5_bit_dac_0[1].VOUT VCC.t204 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X51 switch_n_3v3_0.D3.t1 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.DX_ VCC.t186 VCC.t185 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X52 a_1556_15142# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 VCC.t3 VCC.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X53 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VREFH VSS.t2 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X54 5_bit_dac_0[0].4_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VCC.t16 VCC.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X55 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 VCC.t213 VCC.t212 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X56 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 5_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VCC.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X57 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.DX_ switch_n_3v3_0.D3.t2 VCC.t126 VCC.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X58 5_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS.t210 VSS.t209 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X59 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 a_1556_11458# VSS.t278 VSS.t277 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X60 5_bit_dac_0[0].VOUT D4_BUF.t2 5_bit_dac_0[0].4_bit_dac_0[0].VOUT VSS.t242 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X61 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t132 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X62 5_bit_dac_0[1].4_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VCC.t51 VCC.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X63 D3_BUF.t0 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.DX_ VSS.t20 VSS.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X64 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 VSS.t317 VSS.t316 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X65 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VREFH VSS.t2 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X66 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 a_1556_12686# VCC.t96 VCC.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X67 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t211 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X68 D4_BUF.t0 5_bit_dac_0[0].switch_n_3v3_0.DX_ VSS.t69 VSS.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X69 5_bit_dac_0[0].4_bit_dac_0[0].VOUT 5_bit_dac_0[0].switch_n_3v3_0.DX_ 5_bit_dac_0[0].VOUT VCC.t61 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X70 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X71 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.DX_ D3.t0 VSS.t271 VSS.t270 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X72 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].VREFH VSS.t2 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X73 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.DX_ 5_bit_dac_0[1].switch_n_3v3_0.D3 VCC.t148 VCC.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X74 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_15142# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X75 switch_n_3v3_0.D4.t0 5_bit_dac_0[1].switch_n_3v3_0.DX_ VSS.t217 VSS.t216 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X76 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 VSS.t97 VSS.t96 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X77 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X78 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].VREFH VSS.t2 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X79 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X80 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t29 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X81 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_12686# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X82 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 VCC.t19 VCC.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X83 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS.t165 VSS.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X84 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS.t207 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X85 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VCC.t313 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X86 a_1556_1634# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 VCC.t40 VCC.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X87 a_1556_6546# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 VSS.t16 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X88 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[1].VREFH VSS.t29 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X89 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X90 5_bit_dac_0[1].4_bit_dac_0[1].VOUT 5_bit_dac_0[1].switch_n_3v3_0.DX_ 5_bit_dac_0[1].VOUT VSS.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X91 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X92 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VCC.t87 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X93 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VCC.t160 VCC.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X94 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_10230# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L VCC.t303 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X95 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_18826# VREFL.t1 VSS.t260 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X96 a_1556_4090# 5_bit_dac_0[0].4_bit_dac_0[0].D0 VCC.t86 VCC.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X97 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X98 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VCC.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X99 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_16370# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L VCC.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X100 5_bit_dac_0[1].4_bit_dac_0[0].D0 a_1556_15142# VSS.t32 VSS.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X101 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X102 5_bit_dac_0[1].switch_n_3v3_0.DX_ D4.t0 VSS.t46 VSS.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X103 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ VSS.t66 VSS.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X104 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VOUT VCC.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X105 5_bit_dac_0[0].VOUT switch_n_3v3_0.DX_ VOUT.t3 VCC.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X106 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_7774# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t229 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X107 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t2 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X108 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].VOUT VCC.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X109 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_5318# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L VCC.t168 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X110 a_1556_4090# 5_bit_dac_0[0].4_bit_dac_0[0].D0 VSS.t93 VSS.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X111 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_16370# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VREFH VSS.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X112 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X113 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 VSS.t286 VSS.t285 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X114 VREFL.t2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t283 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X115 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VCC.t250 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X116 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VCC.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X117 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_13914# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L VCC.t190 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X118 a_1556_7774# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 VCC.t117 VCC.t116 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X119 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X120 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VOUT VCC.t228 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X121 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 a_1556_1634# VCC.t219 VCC.t218 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X122 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 a_1556_6546# VSS.t252 VSS.t251 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X123 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X124 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS.t303 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X125 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 a_1556_4090# VCC.t109 VCC.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X126 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t190 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X127 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_9002# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L VCC.t112 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X128 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t240 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X129 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t220 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X130 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_406# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L VCC.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X131 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_2862# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X132 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_5318# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X133 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VSS.t238 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X134 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t29 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X135 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 VSS.t171 VSS.t170 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X136 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 a_1556_4090# VSS.t114 VSS.t113 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X137 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VSS.t315 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X138 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X139 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X140 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 VCC.t166 VCC.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X141 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X142 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VCC.t267 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X143 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t293 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X144 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X145 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].VOUT VSS.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X146 a_1556_12686# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 VSS.t206 VSS.t205 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X147 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X148 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 a_1556_7774# VCC.t224 VCC.t223 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X149 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VCC.t1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X150 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.DX_ 5_bit_dac_0[0].switch_n_3v3_0.D3 VSS.t181 VSS.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X151 a_1556_10230# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 VCC.t100 VCC.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X152 a_1556_18826# D0.t0 VSS.t103 VSS.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X153 5_bit_dac_0[0].switch_n_3v3_0.DX_ switch_n_3v3_0.D4.t3 VSS.t137 VSS.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X154 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X155 a_1556_406# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 VSS.t302 VSS.t301 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X156 D0_BUF.t1 a_1556_406# VSS.t76 VSS.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X157 a_1556_16370# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 VCC.t135 VCC.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X158 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS.t299 VSS.t298 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X159 5_bit_dac_0[0].4_bit_dac_0[1].VOUT 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].VOUT VSS.t179 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X160 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_9002# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X161 5_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VCC.t203 VCC.t202 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X162 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VOUT switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS.t184 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X163 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS.t256 VSS.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X164 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VSS.t163 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X165 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VSS.t297 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X166 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].D1 VSS.t140 VSS.t139 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X167 5_bit_dac_0[1].4_bit_dac_0[1].VOUT 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].VOUT VSS.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X168 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t257 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X169 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VCC.t139 VCC.t138 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X170 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X171 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VSS.t254 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X172 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_17598# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X173 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].D1 VCC.t124 VCC.t123 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X174 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t29 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X175 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 VSS.t237 VSS.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X176 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_13914# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t197 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X177 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VCC.t200 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X178 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t169 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X179 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ VSS.t234 VSS.t233 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X180 a_1556_16370# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 VSS.t143 VSS.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X181 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VCC.t216 VCC.t215 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X182 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS.t200 VSS.t199 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X183 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VCC.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X184 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 VCC.t92 VCC.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X185 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t2 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X186 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ D1.t0 VSS.t28 VSS.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X187 switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ VCC.t288 VCC.t287 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X188 5_bit_dac_0[1].4_bit_dac_0[0].VOUT switch_n_3v3_0.D3.t3 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VOUT VCC.t127 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X189 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VOUT VSS.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X190 a_1556_13914# 5_bit_dac_0[1].4_bit_dac_0[0].D0 VCC.t46 VCC.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X191 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VCC.t157 VCC.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X192 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ switch_n_3v3_0.D2 VSS.t183 VSS.t182 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X193 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VOUT VSS.t232 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X194 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 VCC.t256 VCC.t255 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X195 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t278 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X196 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 a_1556_17598# VSS.t40 VSS.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X197 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS.t147 VSS.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X198 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VSS.t214 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X199 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t62 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X200 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 a_1556_13914# VSS.t196 VSS.t195 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X201 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].VOUT VCC.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X202 D2_BUF.t0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ VSS.t87 VSS.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X203 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VCC.t196 VCC.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X204 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t145 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X205 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[1].switch_n_3v3_0.D2 VSS.t44 VSS.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X206 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t2 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X207 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VSS.t145 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X208 5_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ VCC.t54 VCC.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X209 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VOUT VCC.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X210 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 VCC.t312 VCC.t311 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X211 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT D1_BUF.t2 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t55 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X212 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 5_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VCC.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X213 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 VSS.t263 VSS.t262 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X214 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_18826# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH VCC.t254 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X215 a_1556_2862# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 VSS.t314 VSS.t313 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X216 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VREFH VSS.t29 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X217 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X218 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ VCC.t263 VCC.t262 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X219 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VCC.t297 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X220 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t246 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X221 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VOUT VSS.t294 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X222 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_11458# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VREFH VSS.t276 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X223 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X224 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VCC.t281 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X225 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].D1 VCC.t144 VCC.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X226 a_1556_5318# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 VSS.t245 VSS.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X227 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t29 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X228 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X229 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VCC.t310 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X230 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VCC.t234 VCC.t233 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X231 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X232 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t133 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X233 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].VOUT VSS.t308 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X234 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VCC.t104 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X235 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_12686# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L VCC.t94 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X236 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X237 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t241 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X238 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_406# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH VCC.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X239 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 a_1556_18826# VCC.t253 VCC.t252 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X240 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ D2.t0 VCC.t290 VCC.t289 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X241 D3_BUF.t1 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.DX_ VCC.t13 VCC.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X242 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].VOUT VCC.t142 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X243 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_6546# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VREFH VSS.t250 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X244 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_1634# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L VCC.t217 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X245 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].VOUT VCC.t184 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X246 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t312 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X247 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L D0_BUF.t3 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS.t134 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X248 D1_BUF.t0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS.t161 VSS.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X249 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_4090# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L VCC.t107 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X250 5_bit_dac_0[0].4_bit_dac_0[0].VOUT D3_BUF.t2 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VOUT VCC.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X251 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS.t274 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X252 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t44 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X253 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_15142# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X254 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VCC.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X255 a_1556_9002# 5_bit_dac_0[0].D0 VSS.t273 VSS.t272 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X256 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH D0_BUF.t4 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X257 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VCC.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X258 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X259 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_4090# 5_bit_dac_0[0].4_bit_dac_0[1].VREFH VSS.t112 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X260 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 a_1556_2862# VSS.t79 VSS.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X261 5_bit_dac_0[0].4_bit_dac_0[0].D0 a_1556_5318# VSS.t177 VSS.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X262 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X263 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_7774# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L VCC.t222 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X264 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t84 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X265 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_1634# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t227 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X266 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH VREFH.t0 VSS.t2 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X267 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_6546# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH VCC.t247 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X268 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VREFH VSS.t29 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X269 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VSS.t198 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X270 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].VREFH VSS.t29 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X271 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 VCC.t121 VCC.t120 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X272 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 VSS.t249 VSS.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X273 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X274 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t105 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X275 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].D1 VCC.t131 VCC.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X276 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t284 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X277 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X278 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 a_1556_9002# VSS.t118 VSS.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X279 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VCC.t273 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X280 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].VOUT VSS.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X281 a_1556_11458# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 VSS.t282 VSS.t281 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X282 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t153 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X283 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 VSS.t213 VSS.t212 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X284 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 VCC.t260 VCC.t259 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X285 5_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t115 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X286 a_1556_12686# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 VCC.t199 VCC.t198 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X287 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT D1_BUF.t3 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X288 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS.t187 VSS.t186 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X289 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 5_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X290 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_2862# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH VCC.t71 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X291 VOUT.t1 D5_BUF.t3 5_bit_dac_0[0].VOUT VSS.t211 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X292 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS.t111 VSS.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X293 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X294 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VCC.t293 VCC.t292 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X295 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X296 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X297 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 VCC.t162 VCC.t161 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X298 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X299 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_11458# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH VCC.t271 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X300 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS.t289 VSS.t288 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X301 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 VSS.t189 VSS.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X302 a_1556_15142# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 VSS.t5 VSS.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X303 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_17598# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH VCC.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X304 5_bit_dac_0[0].4_bit_dac_0[1].VOUT 5_bit_dac_0[0].switch_n_3v3_0.DX_ 5_bit_dac_0[0].VOUT VSS.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X305 5_bit_dac_0[0].4_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS.t22 VSS.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X306 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VCC.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X307 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.DX_ VCC.t306 VCC.t305 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X308 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 VSS.t219 VSS.t218 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X309 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 VCC.t231 VCC.t230 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X310 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VOUT switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VCC.t177 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X311 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.DX_ 5_bit_dac_0[0].switch_n_3v3_0.D3 VCC.t173 VCC.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X312 5_bit_dac_0[1].4_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS.t60 VSS.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X313 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 a_1556_11458# VCC.t270 VCC.t269 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X314 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.DX_ VSS.t150 VSS.t149 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X315 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VREFH VSS.t2 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X316 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t229 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X317 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 a_1556_17598# VCC.t30 VCC.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X318 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS.t58 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X319 D4_BUF.t1 5_bit_dac_0[0].switch_n_3v3_0.DX_ VCC.t60 VCC.t59 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X320 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.DX_ D3.t1 VCC.t236 VCC.t235 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X321 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_10230# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t307 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X322 D5_BUF.t0 switch_n_3v3_0.DX_ VSS.t83 VSS.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X323 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_15142# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH VCC.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X324 5_bit_dac_0[0].VOUT D4_BUF.t3 5_bit_dac_0[0].4_bit_dac_0[1].VOUT VCC.t221 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X325 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS.t280 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X326 switch_n_3v3_0.D4.t1 5_bit_dac_0[1].switch_n_3v3_0.DX_ VCC.t209 VCC.t208 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X327 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X328 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].VREFH VSS.t2 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X329 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 VSS.t25 VSS.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X330 a_1556_1634# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 VSS.t48 VSS.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X331 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_17598# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X332 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t29 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X333 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X334 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VCC.t151 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X335 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X336 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS.t168 VSS.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X337 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VCC.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X338 5_bit_dac_0[1].VOUT switch_n_3v3_0.DX_ VOUT.t2 VSS.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X339 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t266 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X340 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L VREFL.t0 VSS.t29 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X341 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS.t292 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X342 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VCC.t201 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X343 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_13914# 5_bit_dac_0[1].4_bit_dac_0[1].VREFH VSS.t194 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X344 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X345 a_1556_6546# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 VCC.t9 VCC.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X346 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X347 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X348 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VCC.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X349 5_bit_dac_0[0].D0 a_1556_10230# VSS.t306 VSS.t305 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X350 switch_n_3v3_0.DX_ D5.t0 VSS.t11 VSS.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X351 5_bit_dac_0[1].4_bit_dac_0[0].D0 a_1556_15142# VCC.t22 VCC.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X352 5_bit_dac_0[1].switch_n_3v3_0.DX_ D4.t1 VCC.t77 VCC.t76 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X353 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ VSS.t53 VSS.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X354 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_2862# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X355 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t2 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X356 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ VCC.t57 VCC.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X357 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_5318# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X358 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VOUT VCC.t286 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X359 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VCC.t258 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X360 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X361 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X362 5_bit_dac_0[1].4_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t197 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X363 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VCC.t194 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X364 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 VCC.t277 VCC.t276 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X365 a_1556_2862# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 VCC.t309 VCC.t308 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X366 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_18826# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L VCC.t251 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X367 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X368 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 a_1556_1634# VSS.t226 VSS.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X369 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X370 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VOUT VCC.t261 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X371 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 a_1556_6546# VCC.t246 VCC.t245 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X372 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_9002# 5_bit_dac_0[1].VREFH VSS.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X373 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X374 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS.t243 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X375 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t296 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X376 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_406# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X377 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X378 5_bit_dac_0[0].4_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t307 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X379 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_7774# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t228 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X380 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_5318# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH VCC.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X381 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VSS.t287 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X382 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t29 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X383 5_bit_dac_0[1].4_bit_dac_0[0].VOUT switch_n_3v3_0.D3.t4 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VOUT VSS.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X384 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 VSS.t72 VSS.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X385 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VSS.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X386 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 VSS.t173 VSS.t172 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X387 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X388 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X389 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X390 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t204 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X391 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t247 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X392 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS.t311 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X393 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X394 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X395 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 a_1556_2862# VCC.t70 VCC.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X396 a_1556_17598# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 VSS.t291 VSS.t290 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X397 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].VOUT VSS.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X398 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.DX_ switch_n_3v3_0.D3.t5 VSS.t13 VSS.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X399 a_1556_13914# 5_bit_dac_0[1].4_bit_dac_0[0].D0 VSS.t56 VSS.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X400 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X401 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X402 5_bit_dac_0[0].switch_n_3v3_0.DX_ switch_n_3v3_0.D4.t4 VCC.t89 VCC.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X403 5_bit_dac_0[0].4_bit_dac_0[0].VOUT D3_BUF.t3 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].VOUT VSS.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X404 a_1556_406# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 VCC.t295 VCC.t294 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X405 D0_BUF.t0 a_1556_406# VCC.t66 VCC.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X406 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_9002# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH VCC.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X407 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS.t203 VSS.t202 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X408 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 5_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X409 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VCC.t179 VCC.t178 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X410 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X411 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VSS.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X412 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].D1 VSS.t128 VSS.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X413 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_12686# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X414 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VSS.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X415 switch_n_3v3_0.D3.t0 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.DX_ VSS.t193 VSS.t192 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X416 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_10230# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH VCC.t302 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X417 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VCC.t282 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X418 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_18826# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X419 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t70 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X420 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VREFH VSS.t2 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X421 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VCC.t214 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X422 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS.t222 VSS.t221 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X423 D5_BUF.t1 switch_n_3v3_0.DX_ VCC.t74 VCC.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X424 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ VSS.t269 VSS.t268 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X425 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].D1 VSS.t152 VSS.t151 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X426 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].VOUT VSS.t191 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X427 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t2 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X428 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_16370# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH VCC.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X429 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VOUT VSS.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X430 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VCC.t155 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X431 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VCC.t192 VCC.t191 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X432 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[0].switch_n_3v3_0.D2 VSS.t89 VSS.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X433 5_bit_dac_0[1].4_bit_dac_0[1].VOUT 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VOUT VCC.t146 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X434 5_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ VCC.t5 VCC.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X435 a_1556_18826# D0.t1 VCC.t36 VCC.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X436 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 VCC.t182 VCC.t181 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X437 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VOUT VSS.t267 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X438 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ switch_n_3v3_0.D2 VCC.t176 VCC.t175 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X439 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 a_1556_12686# VSS.t99 VSS.t98 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X440 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VCC.t164 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X441 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.DX_ 5_bit_dac_0[1].switch_n_3v3_0.D3 VSS.t155 VSS.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X442 5_bit_dac_0[0].D0 a_1556_10230# VCC.t301 VCC.t300 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X443 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 a_1556_18826# VSS.t258 VSS.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X444 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VSS.t264 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X445 5_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ VSS.t62 VSS.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X446 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].VOUT VCC.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X447 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VCC.t249 VCC.t248 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X448 D2_BUF.t1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ VCC.t79 VCC.t78 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X449 switch_n_3v3_0.DX_ D5.t1 VCC.t299 VCC.t298 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X450 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VSS.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X451 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ D2.t1 VSS.t132 VSS.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X452 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VCC.t154 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X453 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t2 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X454 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 a_1556_16370# VCC.t25 VCC.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X455 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ VCC.t42 VCC.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X456 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VSS.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X457 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 VCC.t150 VCC.t149 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X458 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_16370# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X459 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].VOUT D2_BUF.t3 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VCC.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X460 5_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ VSS.t9 VSS.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X461 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH a_1556_13914# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH VCC.t189 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X462 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t2 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X463 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VCC.t205 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X464 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X465 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS.t104 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X466 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VREFH VSS.t29 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X467 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ VCC.t227 VCC.t226 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X468 5_bit_dac_0[1].VOUT switch_n_3v3_0.D4.t5 5_bit_dac_0[1].4_bit_dac_0[1].VOUT VCC.t90 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X469 a_1556_7774# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 VSS.t121 VSS.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X470 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X471 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].VOUT VSS.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X472 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ D1.t1 VCC.t103 VCC.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X473 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VCC.t239 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X474 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VCC.t232 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X475 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_11458# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L VCC.t268 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X476 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS.t29 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X477 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VCC.t280 VCC.t279 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X478 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS.t1 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X479 a_1556_5318# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 VCC.t238 VCC.t237 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X480 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
X481 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t272 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X482 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VCC.t291 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X483 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_17598# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L VCC.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X484 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 a_1556_16370# VSS.t35 VSS.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X485 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 VSS.t158 VSS.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X486 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t119 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X487 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH a_1556_406# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X488 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 a_1556_13914# VCC.t188 VCC.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X489 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].VOUT VCC.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X490 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[1].switch_n_3v3_0.D2 VCC.t33 VCC.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X491 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_1634# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VREFH VSS.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X492 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.DX_ VCC.t141 VCC.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X493 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].VOUT VCC.t304 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X494 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_6546# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L VCC.t244 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X495 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH D0_BUF.t5 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VCC.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X496 D1_BUF.t1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VCC.t153 VCC.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X497 5_bit_dac_0[0].4_bit_dac_0[1].VOUT 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VOUT VCC.t171 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X498 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X499 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_10230# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS.t304 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=0.5
X500 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_15142# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L VCC.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X501 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VCC.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X502 a_1556_9002# 5_bit_dac_0[0].D0 VCC.t265 VCC.t264 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.5
X503 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS.t0 sky130_fd_pr__res_generic_nd__hv w=0.42 l=2.1
C0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.229f
C1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D6 1.72e-19
C2 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT switch_n_3v3_0.D6 0.0199f
C3 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.00349f
C4 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 0.339f
C5 5_bit_dac_0[0].4_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 0.546f
C6 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.635f
C7 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.00143f
C8 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.00577f
C9 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 D5 2.05e-20
C10 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2.38e-19
C11 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 2.78e-22
C12 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL switch_n_3v3_0.D7 0.00143f
C13 5_bit_dac_0[0].4_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.037f
C14 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00306f
C15 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH a_1556_13914# 0.175f
C16 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.0923f
C17 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.0579f
C18 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5.59e-19
C19 5_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 0.0694f
C20 5_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 3.68e-19
C21 a_1556_11458# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 1.21e-20
C22 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 2.51e-20
C23 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 0.797f
C24 5_bit_dac_0[1].switch_n_3v3_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 9.82e-21
C25 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.579f
C26 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT D3 0.0607f
C27 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.00183f
C28 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.472f
C29 D4 switch_n_3v3_0.D4 0.0541f
C30 a_1556_406# D0_BUF 0.325f
C31 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].VOUT 0.0157f
C32 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L a_1556_9002# 0.403f
C33 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH VREFH 0.0124f
C34 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VREFL 0.404f
C35 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT switch_n_3v3_0.D7 0.0397f
C36 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.765f
C37 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.0107f
C38 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.138f
C39 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.00105f
C40 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.482f
C41 switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.177f
C42 5_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.036f
C43 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.48e-19
C44 5_bit_dac_0[0].4_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 0.0988f
C45 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL switch_n_3v3_0.D7 0.00143f
C46 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.0579f
C47 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.0923f
C48 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.00183f
C49 5_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.177f
C50 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 3.74e-19
C51 5_bit_dac_0[0].4_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3.53e-19
C52 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ switch_n_3v3_0.D7 0.0268f
C53 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.322f
C54 VCC a_1556_5318# 0.713f
C55 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.347f
C56 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3.53e-19
C57 5_bit_dac_0[1].VOUT switch_n_3v3_0.DX_ 0.124f
C58 D2_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.177f
C59 switch_n_3v3_0.D4 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 2.38e-20
C60 5_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 5.68e-19
C61 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.349f
C62 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 1.9e-19
C63 VCC 5_bit_dac_0[0].D0 1.18f
C64 5_bit_dac_0[0].switch_n_3v3_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00394f
C65 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.DX_ 3.53e-19
C66 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 2.38e-19
C67 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.00105f
C68 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.24f
C69 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.504f
C70 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0102f
C71 VCC 5_bit_dac_0[1].VOUT 0.751f
C72 D3_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 3.74e-19
C73 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 8.92e-19
C74 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ D5 2.07e-19
C75 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H a_1556_17598# 0.397f
C76 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 0.0988f
C77 5_bit_dac_0[1].VOUT 5_bit_dac_0[0].VOUT 0.344f
C78 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 0.236f
C79 switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00189f
C80 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL switch_n_3v3_0.D7 0.00143f
C81 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3.36e-19
C82 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00306f
C83 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.132f
C84 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VOUT D5 3.23e-20
C85 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 1.9e-19
C86 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 0.315f
C87 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.303f
C88 D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 8.97e-20
C89 D5 switch_n_3v3_0.DX_ 0.0905f
C90 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.0057f
C91 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 6.14e-19
C92 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0824f
C93 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.00117f
C94 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 1.46e-19
C95 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 D5 0.0663f
C96 D4 5_bit_dac_0[1].switch_n_3v3_0.DX_ 0.0904f
C97 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00163f
C98 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.68e-19
C99 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.511f
C100 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00163f
C101 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT switch_n_3v3_0.D7 0.0397f
C102 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL D1_BUF 4.15e-19
C103 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.511f
C104 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.265f
C105 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].D0 1.9e-19
C106 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].D1 3.54e-19
C107 5_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.177f
C108 VCC D5 0.648f
C109 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.0104f
C110 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH D0_BUF 0.538f
C111 5_bit_dac_0[0].D1 a_1556_9002# 0.003f
C112 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[1].VREFH 0.0104f
C113 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 3.62e-20
C114 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 0.00132f
C115 D5 5_bit_dac_0[0].VOUT 1.26e-20
C116 5_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0701f
C117 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.00577f
C118 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].VREFH 0.0104f
C119 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VREFH D0_BUF 4.97e-19
C120 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.0107f
C121 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.291f
C122 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.189f
C123 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.00819f
C124 VCC a_1556_2862# 0.713f
C125 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 0.00132f
C126 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 0.712f
C127 a_1556_15142# 5_bit_dac_0[1].4_bit_dac_0[0].D0 0.325f
C128 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.00164f
C129 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.805f
C130 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.265f
C131 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH a_1556_15142# 0.175f
C132 5_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 4.62e-19
C133 5_bit_dac_0[1].switch_n_3v3_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 4.09e-19
C134 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00394f
C135 switch_n_3v3_0.D3 D5_BUF 0.0337f
C136 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.00577f
C137 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.836f
C138 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.714f
C139 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.379f
C140 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VOUT switch_n_3v3_0.D6 4.36e-20
C141 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 0.14f
C142 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.00349f
C143 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL switch_n_3v3_0.D6 0.00202f
C144 switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00189f
C145 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.229f
C146 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00143f
C147 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.115f
C148 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].D0 0.00164f
C149 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L a_1556_10230# 0.403f
C150 5_bit_dac_0[1].switch_n_3v3_0.D3 switch_n_3v3_0.D6 0.0625f
C151 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.315f
C152 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 a_1556_5318# 0.003f
C153 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH a_1556_9002# 0.175f
C154 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 3.54e-19
C155 5_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 1.9e-19
C156 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 8.97e-19
C157 a_1556_18826# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 4.09e-19
C158 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT D3_BUF 0.00505f
C159 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 0.0988f
C160 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.229f
C161 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.229f
C162 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 1.81e-20
C163 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.579f
C164 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.DX_ switch_n_3v3_0.D6 2.54e-19
C165 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.00143f
C166 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.635f
C167 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.00319f
C168 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 2.29e-20
C169 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].D0 0.00105f
C170 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 3.82e-19
C171 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.482f
C172 5_bit_dac_0[0].4_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].D1 0.00262f
C173 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 2.29e-20
C174 5_bit_dac_0[1].4_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.00491f
C175 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 0.0124f
C176 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 3.82e-19
C177 D0_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.38f
C178 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5.59e-19
C179 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 2.78e-22
C180 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT switch_n_3v3_0.D7 0.0397f
C181 a_1556_13914# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 4.09e-19
C182 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H a_1556_12686# 4.83e-19
C183 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 switch_n_3v3_0.D2 1.48e-19
C184 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.176f
C185 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D6 1.72e-19
C186 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.39f
C187 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00805f
C188 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 a_1556_406# 0.003f
C189 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.00819f
C190 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 1.46e-19
C191 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.404f
C192 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 2.29e-20
C193 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.DX_ 1.34e-20
C194 5_bit_dac_0[1].4_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0551f
C195 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT switch_n_3v3_0.D3 0.00505f
C196 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.229f
C197 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH VREFL 0.201f
C198 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.394f
C199 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.088f
C200 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.138f
C201 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 2.78e-19
C202 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 0.0155f
C203 a_1556_6546# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 2.93e-19
C204 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5.89e-20
C205 a_1556_4090# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 6.04e-19
C206 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.229f
C207 VCC a_1556_15142# 0.713f
C208 5_bit_dac_0[1].4_bit_dac_0[0].VOUT switch_n_3v3_0.D6 4.7e-20
C209 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.347f
C210 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00473f
C211 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.394f
C212 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_9002# 0.00538f
C213 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.303f
C214 a_1556_11458# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 4.09e-19
C215 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H a_1556_10230# 4.83e-19
C216 5_bit_dac_0[1].4_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2.38e-19
C217 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 1.9e-19
C218 5_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.265f
C219 D1 D2 0.00881f
C220 switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 1.75e-20
C221 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 0.00426f
C222 switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.DX_ 0.0904f
C223 switch_n_3v3_0.D4 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 0.0888f
C224 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 6.14e-19
C225 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 0.0124f
C226 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[0].VOUT 4.14e-20
C227 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ switch_n_3v3_0.D7 0.0268f
C228 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ D3_BUF 8.04e-20
C229 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].D1 0.0757f
C230 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 a_1556_16370# 0.003f
C231 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].D0 0.00105f
C232 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5.59e-19
C233 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 2.29e-20
C234 5_bit_dac_0[1].4_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 4.97e-19
C235 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH switch_n_3v3_0.D6 6.1e-19
C236 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 1.34e-20
C237 D4_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00116f
C238 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 9.68e-20
C239 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 0.0124f
C240 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.836f
C241 a_1556_9002# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 2.93e-19
C242 5_bit_dac_0[0].4_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 0.302f
C243 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.00319f
C244 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 1.46e-19
C245 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 1.9e-19
C246 D3 D4 1.02f
C247 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5.89e-20
C248 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH D0 0.0572f
C249 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 3.54e-19
C250 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL D5 0.00306f
C251 switch_n_3v3_0.D4 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00517f
C252 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.322f
C253 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D7 1.45e-19
C254 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.14f
C255 5_bit_dac_0[0].4_bit_dac_0[0].D1 switch_n_3v3_0.D6 1.79e-20
C256 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.00213f
C257 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].switch_n_3v3_0.DX_ 3.68e-19
C258 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5.84e-19
C259 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].VREFH 0.0124f
C260 a_1556_7774# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 6.04e-19
C261 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 0.14f
C262 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ D3_BUF 6.07e-19
C263 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ D5 1.8e-19
C264 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.312f
C265 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 1.7e-19
C266 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 5_bit_dac_0[1].switch_n_3v3_0.D3 0.15f
C267 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 1.06f
C268 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 7.75e-19
C269 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0668f
C270 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 3.54e-19
C271 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.DX_ D5 1.8e-19
C272 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 2.34e-21
C273 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH D0_BUF 0.00164f
C274 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.472f
C275 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 0.628f
C276 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 0.525f
C277 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT switch_n_3v3_0.D7 0.0324f
C278 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.312f
C279 switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.613f
C280 5_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 0.0477f
C281 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].switch_n_3v3_0.D2 0.0694f
C282 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH a_1556_11458# 1.97e-19
C283 5_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.613f
C284 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH D4 0.00127f
C285 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D6 1.72e-19
C286 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00189f
C287 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.00114f
C288 VCC 5_bit_dac_0[1].switch_n_3v3_0.D3 0.773f
C289 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.DX_ 3.53e-19
C290 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00143f
C291 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.635f
C292 5_bit_dac_0[0].D0 5_bit_dac_0[0].D1 0.00262f
C293 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5.59e-19
C294 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.00819f
C295 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.0757f
C296 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.0179f
C297 VCC 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.DX_ 0.712f
C298 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH switch_n_3v3_0.D6 6.1e-19
C299 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.302f
C300 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 1.7e-19
C301 D2_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.546f
C302 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[0].D1 3.54e-20
C303 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 switch_n_3v3_0.D7 1.57e-20
C304 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH switch_n_3v3_0.D7 4.71e-19
C305 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0927f
C306 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT switch_n_3v3_0.D7 0.0324f
C307 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.68e-19
C308 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.115f
C309 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 0.219f
C310 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.236f
C311 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.714f
C312 a_1556_15142# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.00365f
C313 5_bit_dac_0[1].4_bit_dac_0[0].D0 a_1556_13914# 0.0981f
C314 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.00368f
C315 switch_n_3v3_0.D4 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00517f
C316 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.115f
C317 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH a_1556_13914# 9.57e-20
C318 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 0.00262f
C319 5_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.0211f
C320 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 0.14f
C321 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 D3 3.11e-20
C322 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00805f
C323 a_1556_6546# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 4.09e-19
C324 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H a_1556_5318# 4.83e-19
C325 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.291f
C326 5_bit_dac_0[1].4_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 0.00231f
C327 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 8.92e-19
C328 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0701f
C329 D2 switch_n_3v3_0.D7 0.0518f
C330 5_bit_dac_0[0].switch_n_3v3_0.DX_ D4_BUF 0.219f
C331 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.051f
C332 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 2.34e-21
C333 5_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.0824f
C334 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0927f
C335 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3.53e-19
C336 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 3.62e-20
C337 VCC 5_bit_dac_0[1].4_bit_dac_0[0].VOUT 0.441f
C338 5_bit_dac_0[0].D1 D5 4.65e-19
C339 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.504f
C340 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VOUT switch_n_3v3_0.D7 0.0191f
C341 switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 3.11e-20
C342 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.0259f
C343 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 1.9e-19
C344 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.005f
C345 5_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.613f
C346 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 0.0104f
C347 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H a_1556_406# 4.83e-19
C348 a_1556_1634# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 4.09e-19
C349 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ D4 1.33e-19
C350 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.39f
C351 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 1.46e-19
C352 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 6.14e-19
C353 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.347f
C354 D5_BUF switch_n_3v3_0.D6 4.68f
C355 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0801f
C356 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L a_1556_5318# 0.403f
C357 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D6 1.72e-19
C358 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0801f
C359 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 0.0104f
C360 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.622f
C361 D3_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.0204f
C362 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH switch_n_3v3_0.D6 6.1e-19
C363 switch_n_3v3_0.D4 switch_n_3v3_0.D3 2.53f
C364 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.128f
C365 switch_n_3v3_0.D4 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 2.51e-19
C366 D4_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00116f
C367 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H a_1556_4090# 0.397f
C368 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.0104f
C369 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 4.15e-19
C370 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 0.00262f
C371 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.0102f
C372 D3_BUF switch_n_3v3_0.D7 0.0405f
C373 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].VOUT switch_n_3v3_0.D6 4.32e-20
C374 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D7 1.45e-19
C375 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.68e-19
C376 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 switch_n_3v3_0.D6 1.79e-20
C377 5_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 2.96e-19
C378 5_bit_dac_0[0].4_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.0745f
C379 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.835f
C380 VCC a_1556_13914# 0.713f
C381 switch_n_3v3_0.D4 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00517f
C382 5_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.38f
C383 VCC 5_bit_dac_0[0].4_bit_dac_0[0].D1 0.797f
C384 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.177f
C385 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 9.82e-21
C386 a_1556_7774# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.00365f
C387 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 a_1556_6546# 0.0981f
C388 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.24f
C389 switch_n_3v3_0.D2 switch_n_3v3_0.D7 0.0916f
C390 D3 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 2.69e-19
C391 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.38f
C392 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ D5 2.07e-19
C393 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D7 1.45e-19
C394 D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00872f
C395 5_bit_dac_0[1].4_bit_dac_0[0].D1 switch_n_3v3_0.D6 1.79e-20
C396 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5.89e-20
C397 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.176f
C398 a_1556_16370# a_1556_15142# 0.00981f
C399 5_bit_dac_0[1].VREFH a_1556_9002# 0.337f
C400 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.176f
C401 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ switch_n_3v3_0.D7 0.0268f
C402 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT switch_n_3v3_0.D6 0.0258f
C403 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.00368f
C404 D5_BUF 5_bit_dac_0[0].switch_n_3v3_0.D3 0.0849f
C405 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 2.07e-19
C406 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.205f
C407 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT switch_n_3v3_0.D7 0.0324f
C408 a_1556_2862# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.00365f
C409 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 a_1556_1634# 0.0981f
C410 VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.00583f
C411 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.00213f
C412 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 3.47e-20
C413 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 8.92e-19
C414 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.138f
C415 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 3.82e-19
C416 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT switch_n_3v3_0.D4 0.00505f
C417 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].VOUT D4_BUF 1.79e-20
C418 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.00114f
C419 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.714f
C420 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.DX_ 7.51e-19
C421 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.0204f
C422 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 1.85e-19
C423 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.176f
C424 5_bit_dac_0[0].4_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 3.54e-19
C425 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 1.26e-20
C426 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 2.51e-20
C427 a_1556_6546# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 1.21e-20
C428 a_1556_10230# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 4.09e-19
C429 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].VOUT D4 2.45e-20
C430 D5 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00894f
C431 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5.89e-20
C432 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 4.81e-19
C433 switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.0222f
C434 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.0579f
C435 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.0923f
C436 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.622f
C437 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.0107f
C438 a_1556_2862# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2.93e-19
C439 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 2.78e-22
C440 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.DX_ switch_n_3v3_0.D6 2.54e-19
C441 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.00114f
C442 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[1].switch_n_3v3_0.D3 6.07e-19
C443 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5.89e-20
C444 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3.36e-19
C445 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH a_1556_16370# 0.175f
C446 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.138f
C447 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L a_1556_11458# 1.29e-19
C448 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 4.5e-19
C449 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 1.81e-20
C450 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.0261f
C451 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].VOUT 0.0157f
C452 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.051f
C453 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.836f
C454 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.DX_ 5_bit_dac_0[1].switch_n_3v3_0.D3 0.219f
C455 D4_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 2.38e-20
C456 switch_n_3v3_0.D4 5_bit_dac_0[0].4_bit_dac_0[0].VOUT 1.26e-20
C457 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 1.06e-19
C458 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.005f
C459 5_bit_dac_0[1].switch_n_3v3_0.D2 switch_n_3v3_0.D6 0.0618f
C460 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 0.00237f
C461 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH D5 8.21e-19
C462 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5.55e-20
C463 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.00319f
C464 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH a_1556_4090# 1.97e-19
C465 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.115f
C466 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.482f
C467 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 0.00105f
C468 5_bit_dac_0[1].4_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].D1 0.00262f
C469 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.00819f
C470 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.00183f
C471 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].D1 0.00375f
C472 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.176f
C473 D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0778f
C474 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.00577f
C475 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5.84e-19
C476 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ D2_BUF 0.00132f
C477 switch_n_3v3_0.DX_ D5_BUF 0.219f
C478 5_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 0.0904f
C479 a_1556_9002# a_1556_7774# 0.00981f
C480 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.303f
C481 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VOUT 0.0113f
C482 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2.38e-19
C483 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT D4 0.0259f
C484 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 2.96e-19
C485 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].D1 0.044f
C486 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.DX_ 5_bit_dac_0[0].switch_n_3v3_0.D3 0.219f
C487 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0927f
C488 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.24f
C489 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.DX_ 1.79e-20
C490 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].switch_n_3v3_0.DX_ 0.00373f
C491 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 5_bit_dac_0[0].switch_n_3v3_0.DX_ 1.05e-19
C492 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3.38e-20
C493 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 D0_BUF 0.0179f
C494 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00872f
C495 VCC D5_BUF 0.714f
C496 a_1556_13914# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.325f
C497 a_1556_5318# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2.93e-19
C498 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.805f
C499 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.00319f
C500 D4 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 2.69e-19
C501 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].D1 6.11e-19
C502 D5_BUF 5_bit_dac_0[0].VOUT 0.176f
C503 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.111f
C504 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.714f
C505 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].D0 0.00105f
C506 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.482f
C507 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.125f
C508 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL switch_n_3v3_0.D6 0.00202f
C509 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.125f
C510 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.622f
C511 D4_BUF 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.DX_ 1.33e-19
C512 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 2.29e-20
C513 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 0.338f
C514 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 0.797f
C515 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 2.34e-21
C516 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL switch_n_3v3_0.D7 0.00143f
C517 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0018f
C518 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 1.9e-19
C519 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L a_1556_2862# 0.403f
C520 5_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 0.00179f
C521 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.125f
C522 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL D5 0.00306f
C523 5_bit_dac_0[0].4_bit_dac_0[0].D0 a_1556_4090# 0.0981f
C524 a_1556_5318# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.00365f
C525 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.DX_ 0.0104f
C526 5_bit_dac_0[1].4_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 1.48e-19
C527 a_1556_18826# D1 0.003f
C528 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 2.51e-20
C529 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.0018f
C530 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 0.552f
C531 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.613f
C532 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.0102f
C533 VCC 5_bit_dac_0[1].4_bit_dac_0[0].D1 0.797f
C534 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.0261f
C535 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3.82e-19
C536 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 2.34e-21
C537 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.322f
C538 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 8.92e-19
C539 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.529f
C540 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 0.00375f
C541 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.0172f
C542 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 0.00237f
C543 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.00692f
C544 VCC a_1556_1634# 0.713f
C545 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].switch_n_3v3_0.D2 0.00132f
C546 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.0579f
C547 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 2.29e-20
C548 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.0923f
C549 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ D5 1.8e-19
C550 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.0172f
C551 VREFH a_1556_406# 2.68e-20
C552 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 8.92e-19
C553 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.0261f
C554 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5.59e-19
C555 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D7 1.45e-19
C556 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3.82e-19
C557 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.125f
C558 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 switch_n_3v3_0.D6 1.79e-20
C559 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.00692f
C560 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].D0 0.00349f
C561 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH a_1556_17598# 0.337f
C562 D3_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 1.15e-19
C563 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.0018f
C564 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.138f
C565 VCC 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.DX_ 0.712f
C566 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 1.79e-20
C567 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0102f
C568 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_2862# 0.00538f
C569 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].switch_n_3v3_0.D3 8.04e-20
C570 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 2.66e-20
C571 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VREFH a_1556_12686# 2.68e-20
C572 5_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.0129f
C573 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.39f
C574 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.236f
C575 5_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.DX_ 3.14e-19
C576 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.651f
C577 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.037f
C578 switch_n_3v3_0.D4 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.0259f
C579 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 switch_n_3v3_0.D7 1.57e-20
C580 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.651f
C581 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0018f
C582 5_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 0.0694f
C583 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH switch_n_3v3_0.D7 5.14e-19
C584 switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.00213f
C585 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.0104f
C586 5_bit_dac_0[1].VREFH 5_bit_dac_0[0].D0 1.06f
C587 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 1.79e-20
C588 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL D5 0.00306f
C589 switch_n_3v3_0.D4 switch_n_3v3_0.D6 0.0852f
C590 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 0.0124f
C591 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH switch_n_3v3_0.D7 4.71e-19
C592 VCC 5_bit_dac_0[1].switch_n_3v3_0.D2 0.779f
C593 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 3.7e-20
C594 5_bit_dac_0[0].switch_n_3v3_0.D2 switch_n_3v3_0.D7 0.0916f
C595 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.291f
C596 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 2.05e-20
C597 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.394f
C598 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.128f
C599 5_bit_dac_0[0].4_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.138f
C600 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.805f
C601 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5.84e-19
C602 a_1556_4090# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 0.00365f
C603 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 a_1556_2862# 0.0981f
C604 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_12686# 0.00538f
C605 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.128f
C606 5_bit_dac_0[1].4_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 3.54e-19
C607 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.315f
C608 5_bit_dac_0[1].4_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 0.0988f
C609 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.00805f
C610 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.115f
C611 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3.53e-19
C612 D5 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 2.71e-19
C613 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 1.9e-19
C614 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.265f
C615 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 7.75e-19
C616 5_bit_dac_0[0].4_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.0295f
C617 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 3.7e-20
C618 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.128f
C619 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 0.24f
C620 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 6.11e-19
C621 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.111f
C622 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 switch_n_3v3_0.D7 1.57e-20
C623 switch_n_3v3_0.D4 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 2.52e-20
C624 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2.38e-19
C625 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 0.0744f
C626 D4 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.00147f
C627 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.00577f
C628 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.579f
C629 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 D3 0.628f
C630 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.404f
C631 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 1.7e-19
C632 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.0222f
C633 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00189f
C634 D4_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 2.52e-20
C635 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.312f
C636 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3.53e-19
C637 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 0.315f
C638 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.00805f
C639 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].VOUT 3.47e-20
C640 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.394f
C641 switch_n_3v3_0.D4 5_bit_dac_0[0].switch_n_3v3_0.D3 1.25f
C642 5_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.046f
C643 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VREFH 0.0988f
C644 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0824f
C645 switch_n_3v3_0.D4 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 2.51e-19
C646 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].D0 0.132f
C647 5_bit_dac_0[1].4_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.0179f
C648 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0824f
C649 5_bit_dac_0[0].4_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.00107f
C650 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[0].switch_n_3v3_0.D2 1.48e-19
C651 5_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0145f
C652 5_bit_dac_0[1].4_bit_dac_0[1].VOUT switch_n_3v3_0.D7 0.0151f
C653 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.312f
C654 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH a_1556_18826# 2.68e-20
C655 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 1.34e-20
C656 VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 0.00549f
C657 D5_BUF D2_BUF 0.0293f
C658 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.68e-19
C659 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L a_1556_15142# 0.403f
C660 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.0222f
C661 5_bit_dac_0[1].switch_n_3v3_0.DX_ switch_n_3v3_0.D6 2.54e-19
C662 5_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0801f
C663 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.128f
C664 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H D0_BUF 0.00379f
C665 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3.38e-20
C666 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0824f
C667 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.00832f
C668 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.0261f
C669 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.404f
C670 D3_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.249f
C671 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].VOUT D2_BUF 0.0719f
C672 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.0035f
C673 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 D2_BUF 1.48e-19
C674 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0145f
C675 switch_n_3v3_0.D4 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 1.33e-19
C676 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT D3 0.0236f
C677 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5.84e-19
C678 a_1556_15142# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.296f
C679 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H a_1556_10230# 0.397f
C680 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT D5 0.027f
C681 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.0035f
C682 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0102f
C683 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].VOUT 0.546f
C684 a_1556_18826# a_1556_17598# 0.00981f
C685 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.205f
C686 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].VREFH 0.0988f
C687 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0145f
C688 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 0.00349f
C689 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.0107f
C690 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.037f
C691 5_bit_dac_0[0].4_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.38f
C692 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.138f
C693 a_1556_5318# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 1.21e-20
C694 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].D1 2.51e-20
C695 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.017f
C696 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 9.68e-20
C697 a_1556_13914# a_1556_12686# 0.00981f
C698 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 0.797f
C699 switch_n_3v3_0.D2 VOUT 1.25e-20
C700 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H a_1556_406# 0.397f
C701 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.236f
C702 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.0104f
C703 switch_n_3v3_0.D4 switch_n_3v3_0.DX_ 1.33e-19
C704 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00394f
C705 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0824f
C706 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.0109f
C707 D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0701f
C708 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 1.18f
C709 5_bit_dac_0[1].4_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 1.9e-19
C710 switch_n_3v3_0.D4 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 0.0895f
C711 a_1556_18826# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0892f
C712 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00163f
C713 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.511f
C714 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ switch_n_3v3_0.D2 0.219f
C715 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH switch_n_3v3_0.D7 2.94e-20
C716 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 0.132f
C717 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3.82e-19
C718 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.39f
C719 5_bit_dac_0[0].D1 D5_BUF 1.13e-21
C720 a_1556_10230# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0892f
C721 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 6.14e-19
C722 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VOUT 0.0533f
C723 VCC switch_n_3v3_0.D4 0.981f
C724 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.805f
C725 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 1.7e-19
C726 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00394f
C727 switch_n_3v3_0.D4 5_bit_dac_0[0].VOUT 5.58e-19
C728 a_1556_13914# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0892f
C729 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].D1 1.85e-19
C730 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0801f
C731 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0018f
C732 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 0.0104f
C733 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5.55e-20
C734 5_bit_dac_0[0].4_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 1.48e-19
C735 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 1.03e-19
C736 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VREFH a_1556_7774# 2.68e-20
C737 a_1556_11458# a_1556_10230# 0.00981f
C738 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.088f
C739 VCC a_1556_4090# 0.713f
C740 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.00379f
C741 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 0.0904f
C742 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.349f
C743 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.088f
C744 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.DX_ 0.0104f
C745 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.0261f
C746 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.176f
C747 5_bit_dac_0[0].4_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].D0 1.06f
C748 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 3.82e-19
C749 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00163f
C750 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.511f
C751 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.DX_ 5_bit_dac_0[1].switch_n_3v3_0.D2 6.07e-19
C752 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.138f
C753 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.088f
C754 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0102f
C755 5_bit_dac_0[1].4_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.005f
C756 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.48e-19
C757 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.0119f
C758 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.0179f
C759 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3.36e-19
C760 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0102f
C761 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL switch_n_3v3_0.D6 0.00202f
C762 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 3.7e-20
C763 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 6.14e-19
C764 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.394f
C765 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.00164f
C766 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 8.92e-19
C767 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 D4 2.52e-20
C768 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 4.25e-19
C769 5_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 3.7e-20
C770 5_bit_dac_0[1].4_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 0.0174f
C771 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.511f
C772 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.836f
C773 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00163f
C774 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.138f
C775 5_bit_dac_0[1].switch_n_3v3_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 6.07e-19
C776 D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.007f
C777 a_1556_13914# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 2.93e-19
C778 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 3.7e-20
C779 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.00491f
C780 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 9.68e-20
C781 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VOUT switch_n_3v3_0.D2 0.0719f
C782 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.0102f
C783 VCC 5_bit_dac_0[1].switch_n_3v3_0.DX_ 0.71f
C784 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.00183f
C785 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 0.472f
C786 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.0179f
C787 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00306f
C788 D3 switch_n_3v3_0.D6 0.0326f
C789 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.514f
C790 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D6 1.72e-19
C791 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.0923f
C792 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.0579f
C793 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.088f
C794 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.00491f
C795 switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.00193f
C796 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 1.06e-19
C797 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3.36e-19
C798 D5_BUF 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.0104f
C799 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 D5 2.05e-20
C800 5_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 0.0137f
C801 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].VOUT 3.47e-20
C802 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00123f
C803 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.045f
C804 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 0.00237f
C805 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH D5 8.21e-19
C806 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.314f
C807 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00805f
C808 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].D0 0.24f
C809 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 1.85e-20
C810 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.314f
C811 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT switch_n_3v3_0.D7 0.0397f
C812 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].D1 1.81e-20
C813 a_1556_10230# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 1.21e-20
C814 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.511f
C815 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].D1 2.51e-20
C816 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00163f
C817 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 0.0104f
C818 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].D0 4.97e-19
C819 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.00319f
C820 5_bit_dac_0[0].4_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 4.97e-19
C821 switch_n_3v3_0.D4 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 2.52e-20
C822 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 1.18f
C823 5_bit_dac_0[0].4_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00805f
C824 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 2.34e-21
C825 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0551f
C826 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.0119f
C827 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 1.85e-20
C828 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 0.00375f
C829 VOUT switch_n_3v3_0.D7 0.00688f
C830 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 0.0124f
C831 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 2.34e-21
C832 switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.00213f
C833 D2 D5 0.0322f
C834 a_1556_1634# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.325f
C835 a_1556_11458# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.296f
C836 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 1.06e-19
C837 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 0.219f
C838 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 0.0616f
C839 D4_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.00127f
C840 5_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 0.0988f
C841 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00306f
C842 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L a_1556_13914# 1.29e-19
C843 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.111f
C844 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 6.11e-19
C845 a_1556_16370# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.296f
C846 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.125f
C847 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.0261f
C848 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.115f
C849 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 0.00132f
C850 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH switch_n_3v3_0.D6 6.67e-19
C851 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 2.51e-20
C852 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ switch_n_3v3_0.D7 0.0268f
C853 a_1556_9002# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 1.21e-20
C854 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 0.0104f
C855 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 0.0179f
C856 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.00349f
C857 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT D4 0.0271f
C858 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0172f
C859 5_bit_dac_0[0].4_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.0179f
C860 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H a_1556_7774# 0.397f
C861 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 1.06f
C862 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 1.85e-20
C863 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 2.69e-19
C864 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2.66e-20
C865 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_13914# 0.00538f
C866 a_1556_1634# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.296f
C867 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 0.0189f
C868 5_bit_dac_0[1].VOUT switch_n_3v3_0.D2 0.00297f
C869 5_bit_dac_0[0].4_bit_dac_0[1].VOUT switch_n_3v3_0.D7 0.0151f
C870 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 0.00112f
C871 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.00577f
C872 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.0199f
C873 VREFH D0_BUF 0.281f
C874 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 3.68e-19
C875 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.312f
C876 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].D0 2.29e-20
C877 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.613f
C878 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 3.7e-20
C879 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0824f
C880 5_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.0241f
C881 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 2.34e-21
C882 5_bit_dac_0[1].4_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0801f
C883 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0018f
C884 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.0109f
C885 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5.55e-20
C886 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 1.81e-20
C887 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.00114f
C888 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 0.14f
C889 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0824f
C890 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 3.68e-19
C891 5_bit_dac_0[0].4_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.48e-19
C892 switch_n_3v3_0.D2 D5 0.0353f
C893 switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 2.09e-21
C894 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 2.51e-20
C895 a_1556_2862# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 1.21e-20
C896 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0927f
C897 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ D5 2.07e-19
C898 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL switch_n_3v3_0.D7 0.00143f
C899 a_1556_6546# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.296f
C900 D4_BUF 5_bit_dac_0[0].4_bit_dac_0[0].VOUT 0.177f
C901 VCC a_1556_406# 0.706f
C902 5_bit_dac_0[1].4_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.00583f
C903 switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 4.58e-19
C904 D3_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.0201f
C905 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 3.38e-20
C906 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.312f
C907 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ switch_n_3v3_0.D6 2.54e-19
C908 D1_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.176f
C909 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.189f
C910 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH a_1556_7774# 0.337f
C911 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.511f
C912 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00163f
C913 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VOUT D3 2.78e-19
C914 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 1.9e-19
C915 a_1556_16370# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.325f
C916 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L a_1556_6546# 1.29e-19
C917 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.394f
C918 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.805f
C919 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT D5 0.0492f
C920 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00394f
C921 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.349f
C922 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0172f
C923 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 7.75e-19
C924 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.189f
C925 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 0.132f
C926 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VOUT switch_n_3v3_0.D7 0.0133f
C927 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.027f
C928 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.0222f
C929 5_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 0.044f
C930 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 1.79e-20
C931 5_bit_dac_0[0].4_bit_dac_0[1].VOUT 5_bit_dac_0[0].switch_n_3v3_0.D2 0.0034f
C932 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.0104f
C933 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 0.00262f
C934 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH a_1556_9002# 9.57e-20
C935 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00306f
C936 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.236f
C937 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.514f
C938 VCC D3 0.331f
C939 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.714f
C940 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.236f
C941 5_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00872f
C942 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH D1 0.00491f
C943 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.128f
C944 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 0.132f
C945 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L a_1556_1634# 1.29e-19
C946 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_17598# 0.00538f
C947 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 1.46e-19
C948 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 switch_n_3v3_0.D7 1.57e-20
C949 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.68e-19
C950 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 3.54e-19
C951 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00473f
C952 switch_n_3v3_0.D4 5_bit_dac_0[0].D1 2.91e-20
C953 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.00123f
C954 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 2.29e-20
C955 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 4.15e-19
C956 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.302f
C957 5_bit_dac_0[0].4_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 0.0104f
C958 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 1.7e-19
C959 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT switch_n_3v3_0.D7 0.0397f
C960 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0018f
C961 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.00832f
C962 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L D1_BUF 2.51e-20
C963 a_1556_406# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 1.21e-20
C964 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH a_1556_5318# 0.175f
C965 VCC 5_bit_dac_0[0].4_bit_dac_0[1].VREFH 0.14f
C966 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5.84e-19
C967 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 0.00375f
C968 a_1556_12686# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 4.09e-19
C969 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H a_1556_11458# 4.83e-19
C970 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.579f
C971 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 0.24f
C972 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].D0 0.132f
C973 5_bit_dac_0[0].switch_n_3v3_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].VOUT 0.0853f
C974 switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 1.26e-20
C975 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.622f
C976 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.463f
C977 a_1556_17598# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 6.04e-19
C978 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 4.15e-19
C979 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 0.132f
C980 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.037f
C981 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 4.81e-19
C982 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].VOUT switch_n_3v3_0.D6 4.32e-20
C983 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.088f
C984 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00189f
C985 5_bit_dac_0[1].VOUT switch_n_3v3_0.D7 0.0126f
C986 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.138f
C987 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 1.06e-19
C988 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].D1 2.51e-20
C989 a_1556_15142# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 1.21e-20
C990 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.218f
C991 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 0.14f
C992 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5.59e-19
C993 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.DX_ 1.34e-20
C994 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.00832f
C995 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 4.25e-19
C996 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D6 1.72e-19
C997 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.0199f
C998 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3.36e-19
C999 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 1.79e-20
C1000 5_bit_dac_0[1].4_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.635f
C1001 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 1.85e-19
C1002 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00805f
C1003 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 1.46e-19
C1004 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H D0_BUF 0.24f
C1005 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH switch_n_3v3_0.D6 6.1e-19
C1006 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 6.14e-19
C1007 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT D1_BUF 1.81e-20
C1008 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.504f
C1009 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.00114f
C1010 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 1.06e-19
C1011 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.805f
C1012 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 4.15e-19
C1013 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5.84e-19
C1014 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L a_1556_13914# 0.403f
C1015 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.037f
C1016 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 3.68e-19
C1017 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH switch_n_3v3_0.D6 6.67e-19
C1018 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.138f
C1019 a_1556_18826# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.296f
C1020 5_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.14f
C1021 D5 switch_n_3v3_0.D7 0.0521f
C1022 a_1556_5318# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0892f
C1023 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3.38e-20
C1024 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].D1 0.219f
C1025 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 1.85e-19
C1026 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 0.544f
C1027 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.315f
C1028 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.312f
C1029 5_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 0.0904f
C1030 a_1556_7774# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.0331f
C1031 D4_BUF switch_n_3v3_0.D6 0.0301f
C1032 a_1556_2862# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.296f
C1033 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.00114f
C1034 switch_n_3v3_0.D4 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00595f
C1035 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 0.044f
C1036 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.504f
C1037 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 0.712f
C1038 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.243f
C1039 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 0.00379f
C1040 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT switch_n_3v3_0.D6 0.0258f
C1041 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VOUT D3_BUF 0.15f
C1042 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.394f
C1043 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ switch_n_3v3_0.D7 0.0268f
C1044 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L a_1556_4090# 1.29e-19
C1045 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00805f
C1046 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 0.00237f
C1047 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0551f
C1048 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH switch_n_3v3_0.D6 6.67e-19
C1049 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT switch_n_3v3_0.D6 0.027f
C1050 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.00213f
C1051 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.0104f
C1052 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D7 1.45e-19
C1053 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT switch_n_3v3_0.D7 0.0265f
C1054 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].D1 0.0757f
C1055 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 switch_n_3v3_0.D6 1.79e-20
C1056 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 0.0124f
C1057 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 8.92e-19
C1058 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0801f
C1059 a_1556_2862# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.0331f
C1060 5_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.129f
C1061 5_bit_dac_0[0].4_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3.36e-19
C1062 switch_n_3v3_0.D4 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00116f
C1063 switch_n_3v3_0.D4 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00517f
C1064 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.514f
C1065 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.DX_ 3.68e-19
C1066 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH a_1556_2862# 0.175f
C1067 D3 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.017f
C1068 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0172f
C1069 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VOUT switch_n_3v3_0.D3 0.15f
C1070 a_1556_11458# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 6.04e-19
C1071 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 4.58e-19
C1072 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 0.255f
C1073 D3_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.00213f
C1074 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH a_1556_11458# 2.68e-20
C1075 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.0104f
C1076 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.39f
C1077 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.DX_ switch_n_3v3_0.D2 6.07e-19
C1078 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ D3 1.03e-19
C1079 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 9.82e-21
C1080 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 D4 0.0888f
C1081 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT D4 0.0547f
C1082 5_bit_dac_0[0].switch_n_3v3_0.D3 D4_BUF 1.25f
C1083 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH a_1556_17598# 9.57e-20
C1084 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH D5 8.21e-19
C1085 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VREFH a_1556_16370# 0.337f
C1086 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.0018f
C1087 D3 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.DX_ 0.0904f
C1088 5_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.037f
C1089 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 1.18f
C1090 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH a_1556_12686# 0.175f
C1091 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH a_1556_6546# 2.68e-20
C1092 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 0.359f
C1093 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.128f
C1094 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 2.09e-21
C1095 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 1.8e-19
C1096 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.00805f
C1097 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0701f
C1098 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0927f
C1099 5_bit_dac_0[0].switch_n_3v3_0.DX_ switch_n_3v3_0.D6 2.54e-19
C1100 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].D0 0.472f
C1101 5_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.00183f
C1102 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.312f
C1103 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.0107f
C1104 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.579f
C1105 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 1.7e-19
C1106 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[0].switch_n_3v3_0.D2 0.219f
C1107 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH switch_n_3v3_0.D6 6.67e-19
C1108 5_bit_dac_0[1].4_bit_dac_0[1].VOUT 5_bit_dac_0[1].VOUT 0.323f
C1109 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.312f
C1110 5_bit_dac_0[1].4_bit_dac_0[0].VOUT switch_n_3v3_0.D2 1.79e-20
C1111 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 0.339f
C1112 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.236f
C1113 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 4.25e-19
C1114 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 0.236f
C1115 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L a_1556_2862# 1.29e-19
C1116 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D6 1.72e-19
C1117 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 D5 2.05e-20
C1118 5_bit_dac_0[1].4_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 0.0104f
C1119 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].VOUT 2.49e-22
C1120 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.24f
C1121 5_bit_dac_0[1].4_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.205f
C1122 switch_n_3v3_0.D4 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00517f
C1123 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT D4 0.0234f
C1124 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 2.07e-19
C1125 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.037f
C1126 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.714f
C1127 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.39f
C1128 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.0104f
C1129 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.13f
C1130 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.00379f
C1131 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.291f
C1132 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 9.82e-21
C1133 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 1.06e-19
C1134 a_1556_12686# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 0.325f
C1135 switch_n_3v3_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 9.82e-21
C1136 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 0.00164f
C1137 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.805f
C1138 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ D2 0.0222f
C1139 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.622f
C1140 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH switch_n_3v3_0.D6 6.1e-19
C1141 5_bit_dac_0[0].4_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.DX_ 0.236f
C1142 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 1.85e-19
C1143 5_bit_dac_0[1].4_bit_dac_0[1].VOUT D5 2.82e-20
C1144 switch_n_3v3_0.D4 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.0271f
C1145 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 2.34e-21
C1146 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ VOUT 5.19e-19
C1147 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.0551f
C1148 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.463f
C1149 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.622f
C1150 a_1556_6546# 5_bit_dac_0[0].4_bit_dac_0[0].D0 0.00365f
C1151 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 a_1556_5318# 0.0981f
C1152 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.544f
C1153 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].D1 6.11e-19
C1154 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.111f
C1155 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.037f
C1156 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].switch_n_3v3_0.DX_ 1.03e-19
C1157 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.0259f
C1158 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].VOUT 2.78e-22
C1159 switch_n_3v3_0.D4 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 4.04e-19
C1160 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 0.0155f
C1161 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.00577f
C1162 a_1556_5318# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.0331f
C1163 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.265f
C1164 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].D0 1.9e-19
C1165 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 0.14f
C1166 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 1.06e-19
C1167 5_bit_dac_0[1].4_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.00319f
C1168 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 0.00164f
C1169 VCC D4_BUF 0.5f
C1170 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.00577f
C1171 VCC a_1556_11458# 0.713f
C1172 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0668f
C1173 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH a_1556_18826# 0.175f
C1174 a_1556_4090# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.296f
C1175 5_bit_dac_0[0].VOUT D4_BUF 0.0748f
C1176 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.177f
C1177 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.529f
C1178 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 0.00237f
C1179 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 0.0155f
C1180 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH switch_n_3v3_0.D6 6.67e-19
C1181 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 0.00426f
C1182 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H a_1556_15142# 0.397f
C1183 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 a_1556_406# 0.0981f
C1184 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 2.38e-19
C1185 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 8.92e-19
C1186 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.765f
C1187 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.622f
C1188 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 0.472f
C1189 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.322f
C1190 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.00577f
C1191 a_1556_17598# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.0331f
C1192 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 0.797f
C1193 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VOUT switch_n_3v3_0.D7 0.0191f
C1194 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L VREFL 0.482f
C1195 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.0259f
C1196 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 0.14f
C1197 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL switch_n_3v3_0.D7 0.00143f
C1198 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].VOUT switch_n_3v3_0.D6 4.32e-20
C1199 switch_n_3v3_0.D4 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.0135f
C1200 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.0035f
C1201 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.0757f
C1202 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.68e-19
C1203 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0801f
C1204 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00189f
C1205 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 4.25e-19
C1206 5_bit_dac_0[1].switch_n_3v3_0.D3 switch_n_3v3_0.D7 0.0924f
C1207 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 1.46e-19
C1208 a_1556_4090# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.325f
C1209 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 0.0104f
C1210 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_406# 0.00538f
C1211 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 0.00426f
C1212 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3.82e-19
C1213 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.0757f
C1214 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.DX_ switch_n_3v3_0.D7 0.0268f
C1215 VCC D0_BUF 0.732f
C1216 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 0.0757f
C1217 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0801f
C1218 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 a_1556_15142# 0.003f
C1219 5_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 3.54e-19
C1220 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ D3 0.00594f
C1221 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 3.62e-20
C1222 switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00872f
C1223 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.189f
C1224 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH a_1556_15142# 0.337f
C1225 D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.111f
C1226 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.0018f
C1227 switch_n_3v3_0.D4 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.0293f
C1228 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 7.75e-19
C1229 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 3.62e-20
C1230 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.48e-19
C1231 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D7 1.45e-19
C1232 switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 0.628f
C1233 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 3.23e-20
C1234 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 switch_n_3v3_0.D6 1.79e-20
C1235 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VOUT VOUT 0.00378f
C1236 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.38f
C1237 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 0.00237f
C1238 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].D1 1.85e-19
C1239 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.00577f
C1240 a_1556_10230# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2.93e-19
C1241 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.291f
C1242 5_bit_dac_0[1].switch_n_3v3_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 0.0104f
C1243 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.14f
C1244 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 0.219f
C1245 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.349f
C1246 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 6.14e-19
C1247 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0145f
C1248 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 0.0757f
C1249 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.265f
C1250 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5.89e-20
C1251 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.DX_ 1.79e-20
C1252 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 1.9e-19
C1253 VCC 5_bit_dac_0[0].switch_n_3v3_0.DX_ 0.71f
C1254 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 0.236f
C1255 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH a_1556_2862# 9.57e-20
C1256 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L D0 0.253f
C1257 5_bit_dac_0[1].4_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.347f
C1258 5_bit_dac_0[0].VOUT 5_bit_dac_0[0].switch_n_3v3_0.DX_ 0.258f
C1259 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 0.177f
C1260 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.504f
C1261 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.622f
C1262 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 0.00375f
C1263 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT D1_BUF 0.0757f
C1264 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 2.49e-22
C1265 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.544f
C1266 5_bit_dac_0[1].4_bit_dac_0[0].VOUT switch_n_3v3_0.D7 0.00725f
C1267 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.236f
C1268 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.0172f
C1269 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 0.0124f
C1270 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.0824f
C1271 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 3.47e-20
C1272 D4 switch_n_3v3_0.D6 0.0328f
C1273 D5_BUF D3_BUF 0.0301f
C1274 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.714f
C1275 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 2.07e-19
C1276 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0927f
C1277 5_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 1.75e-20
C1278 a_1556_10230# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.00365f
C1279 5_bit_dac_0[0].D0 a_1556_9002# 0.0981f
C1280 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].VOUT 2.49e-22
C1281 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.0104f
C1282 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 1.06f
C1283 5_bit_dac_0[1].switch_n_3v3_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00394f
C1284 D0_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5.84e-19
C1285 5_bit_dac_0[0].4_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.00183f
C1286 D3_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 0.177f
C1287 switch_n_3v3_0.D2 D5_BUF 0.0385f
C1288 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.544f
C1289 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 2.49e-22
C1290 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 D3_BUF 4.43e-21
C1291 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.236f
C1292 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 0.219f
C1293 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.00143f
C1294 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.622f
C1295 5_bit_dac_0[1].4_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 9.68e-20
C1296 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 0.0858f
C1297 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH switch_n_3v3_0.D7 4.71e-19
C1298 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.DX_ switch_n_3v3_0.D6 2.54e-19
C1299 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 2.29e-20
C1300 5_bit_dac_0[1].4_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 3.7e-20
C1301 switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00476f
C1302 switch_n_3v3_0.D4 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.0271f
C1303 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 3.38e-20
C1304 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 a_1556_7774# 0.003f
C1305 5_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00476f
C1306 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 3.54e-19
C1307 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 1.85e-19
C1308 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VOUT switch_n_3v3_0.D6 4.36e-20
C1309 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 1.8e-19
C1310 5_bit_dac_0[0].4_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.00262f
C1311 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].D1 0.00375f
C1312 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.00319f
C1313 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.38f
C1314 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT D5_BUF 0.00514f
C1315 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.404f
C1316 5_bit_dac_0[1].VOUT VOUT 0.466f
C1317 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 1.79e-20
C1318 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0551f
C1319 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2.66e-20
C1320 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 2.29e-20
C1321 5_bit_dac_0[0].4_bit_dac_0[0].D1 switch_n_3v3_0.D7 1.57e-20
C1322 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 3.08e-20
C1323 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 0.00262f
C1324 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_10230# 0.00538f
C1325 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.0261f
C1326 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.00819f
C1327 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 1.06f
C1328 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.00114f
C1329 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.DX_ 0.125f
C1330 D2_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00476f
C1331 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 3.82e-19
C1332 5_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 0.0326f
C1333 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.302f
C1334 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.622f
C1335 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.0923f
C1336 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.0579f
C1337 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.00319f
C1338 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 4.15e-19
C1339 switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0269f
C1340 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].D1 0.219f
C1341 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 2.38e-19
C1342 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.088f
C1343 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 0.339f
C1344 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[1].VOUT 0.0743f
C1345 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.0261f
C1346 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 3.38e-20
C1347 D4_BUF D2_BUF 0.0295f
C1348 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D7 1.45e-19
C1349 D5 VOUT 2.49e-20
C1350 5_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 0.00514f
C1351 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 switch_n_3v3_0.D6 1.79e-20
C1352 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.579f
C1353 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.DX_ 0.0904f
C1354 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0801f
C1355 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.DX_ 7.51e-19
C1356 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00473f
C1357 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.00123f
C1358 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.805f
C1359 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 7.75e-19
C1360 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].D1 0.00237f
C1361 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.0107f
C1362 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.005f
C1363 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0102f
C1364 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.037f
C1365 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH switch_n_3v3_0.D7 4.71e-19
C1366 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 9.68e-20
C1367 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ D5 1.8e-19
C1368 5_bit_dac_0[0].4_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.005f
C1369 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.291f
C1370 5_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00476f
C1371 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.349f
C1372 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ D4 2.51e-19
C1373 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 3.82e-19
C1374 5_bit_dac_0[0].4_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.176f
C1375 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3.36e-19
C1376 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L a_1556_1634# 0.403f
C1377 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 0.793f
C1378 switch_n_3v3_0.D4 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.0056f
C1379 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 0.315f
C1380 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 0.00105f
C1381 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H a_1556_13914# 4.83e-19
C1382 a_1556_15142# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 4.09e-19
C1383 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 2.66e-20
C1384 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5.89e-20
C1385 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 3.62e-20
C1386 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.00379f
C1387 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.13f
C1388 5_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[0].D1 0.0189f
C1389 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VOUT D4 2.38e-20
C1390 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.00319f
C1391 VCC a_1556_6546# 0.713f
C1392 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.00349f
C1393 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D3 8.04e-20
C1394 5_bit_dac_0[0].4_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.00319f
C1395 5_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.0211f
C1396 5_bit_dac_0[1].4_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].VOUT 0.34f
C1397 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.00183f
C1398 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3.53e-19
C1399 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5.59e-19
C1400 5_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.176f
C1401 5_bit_dac_0[0].4_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 0.0353f
C1402 5_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.138f
C1403 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.00832f
C1404 5_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 0.0905f
C1405 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0927f
C1406 switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0269f
C1407 VCC D4 0.434f
C1408 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0172f
C1409 switch_n_3v3_0.D4 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.0547f
C1410 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].D0 0.00349f
C1411 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.13f
C1412 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.00379f
C1413 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 1.9e-19
C1414 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH a_1556_13914# 1.97e-19
C1415 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00306f
C1416 5_bit_dac_0[0].4_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.404f
C1417 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0927f
C1418 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 2.49e-22
C1419 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 1.85e-19
C1420 D5_BUF switch_n_3v3_0.D7 0.0408f
C1421 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL D5 0.00306f
C1422 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.0172f
C1423 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 3.62e-20
C1424 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.00819f
C1425 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 9.68e-20
C1426 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.347f
C1427 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.394f
C1428 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT switch_n_3v3_0.D6 0.027f
C1429 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 0.0179f
C1430 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D7 1.45e-19
C1431 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.347f
C1432 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 switch_n_3v3_0.D6 1.79e-20
C1433 5_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3.53e-19
C1434 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH switch_n_3v3_0.D7 4.71e-19
C1435 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.00491f
C1436 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.836f
C1437 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 3.47e-20
C1438 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 0.0744f
C1439 VCC 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.DX_ 0.712f
C1440 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.00577f
C1441 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5.55e-20
C1442 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.635f
C1443 switch_n_3v3_0.D4 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 2.52e-20
C1444 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.00143f
C1445 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.111f
C1446 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ D1_BUF 6.11e-19
C1447 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].VOUT switch_n_3v3_0.D7 0.0133f
C1448 5_bit_dac_0[1].4_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].D0 1.06f
C1449 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 7.75e-19
C1450 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 switch_n_3v3_0.D7 1.57e-20
C1451 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 4.97e-19
C1452 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VOUT D5 3.8e-20
C1453 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 0.524f
C1454 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].VREFH 0.0124f
C1455 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.00164f
C1456 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.347f
C1457 5_bit_dac_0[0].4_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.544f
C1458 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.315f
C1459 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.322f
C1460 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.613f
C1461 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.115f
C1462 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 3.7e-20
C1463 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L a_1556_16370# 0.403f
C1464 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.00491f
C1465 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.38f
C1466 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.115f
C1467 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 D5 2.05e-20
C1468 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 switch_n_3v3_0.D6 0.0618f
C1469 5_bit_dac_0[1].4_bit_dac_0[0].D1 switch_n_3v3_0.D7 1.57e-20
C1470 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.265f
C1471 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 2.07e-19
C1472 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.579f
C1473 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 0.00375f
C1474 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 4.97e-19
C1475 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5.55e-20
C1476 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT switch_n_3v3_0.D7 0.0324f
C1477 a_1556_18826# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 1.21e-20
C1478 switch_n_3v3_0.D4 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 2.38e-20
C1479 a_1556_9002# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 4.09e-19
C1480 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H a_1556_7774# 4.83e-19
C1481 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.68e-19
C1482 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 0.0104f
C1483 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_1634# 0.00538f
C1484 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 1.18f
C1485 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.229f
C1486 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 2.05e-20
C1487 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 1.9e-19
C1488 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.265f
C1489 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00473f
C1490 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 8.97e-19
C1491 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 3.11e-20
C1492 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH a_1556_6546# 9.57e-20
C1493 VREFL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0551f
C1494 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 1.46e-19
C1495 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 0.797f
C1496 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2.66e-20
C1497 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.347f
C1498 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL switch_n_3v3_0.D6 0.00202f
C1499 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.579f
C1500 D4_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00517f
C1501 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 2.96e-19
C1502 D5_BUF 5_bit_dac_0[0].switch_n_3v3_0.D2 0.0616f
C1503 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5.55e-20
C1504 a_1556_6546# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 6.04e-19
C1505 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 0.00375f
C1506 5_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.0222f
C1507 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 7.75e-19
C1508 switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 0.0026f
C1509 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH a_1556_1634# 0.175f
C1510 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.DX_ switch_n_3v3_0.D7 0.0268f
C1511 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].D1 0.219f
C1512 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.0129f
C1513 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.236f
C1514 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH D1_BUF 0.00375f
C1515 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 4.25e-19
C1516 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00872f
C1517 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH a_1556_1634# 9.57e-20
C1518 a_1556_11458# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 2.93e-19
C1519 a_1556_12686# a_1556_11458# 0.00981f
C1520 VCC 5_bit_dac_0[1].4_bit_dac_0[1].VREFH 0.14f
C1521 5_bit_dac_0[1].VOUT D5 2.86e-19
C1522 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 D0_BUF 0.124f
C1523 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.805f
C1524 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].D0 1.9e-19
C1525 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.265f
C1526 5_bit_dac_0[0].4_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.13f
C1527 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[0].switch_n_3v3_0.D3 0.631f
C1528 5_bit_dac_0[0].4_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.00491f
C1529 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.00379f
C1530 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.229f
C1531 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.0211f
C1532 5_bit_dac_0[1].switch_n_3v3_0.D2 switch_n_3v3_0.D7 0.0916f
C1533 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VREFH a_1556_5318# 1.97e-19
C1534 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 1.81e-20
C1535 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.229f
C1536 switch_n_3v3_0.D4 switch_n_3v3_0.D2 0.0617f
C1537 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 a_1556_12686# 0.003f
C1538 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D4 7.1e-20
C1539 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH a_1556_12686# 0.337f
C1540 VREFL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 4.97e-19
C1541 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.0018f
C1542 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH a_1556_9002# 2.68e-20
C1543 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL D0_BUF 0.00349f
C1544 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].D1 0.00237f
C1545 D4_BUF 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 0.0895f
C1546 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.177f
C1547 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.0129f
C1548 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.229f
C1549 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 0.00262f
C1550 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 VREFL 3.54e-19
C1551 D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 1.9e-19
C1552 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 D2_BUF 0.00779f
C1553 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.00819f
C1554 switch_n_3v3_0.D4 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.0263f
C1555 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL D4 0.00517f
C1556 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0269f
C1557 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.051f
C1558 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0172f
C1559 5_bit_dac_0[0].4_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 3.96e-20
C1560 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.312f
C1561 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 0.219f
C1562 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.579f
C1563 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.514f
C1564 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 0.0104f
C1565 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.176f
C1566 VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.0579f
C1567 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.0923f
C1568 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.DX_ 1.34e-20
C1569 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL switch_n_3v3_0.D6 0.00202f
C1570 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ D4 1.33e-19
C1571 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.774f
C1572 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 4.25e-19
C1573 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H a_1556_13914# 0.397f
C1574 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 1.18f
C1575 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 a_1556_10230# 0.003f
C1576 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].D1 0.044f
C1577 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 0.797f
C1578 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH a_1556_10230# 0.337f
C1579 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.128f
C1580 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL switch_n_3v3_0.D7 0.00143f
C1581 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.0018f
C1582 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].D1 3.54e-19
C1583 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 8.92e-19
C1584 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.472f
C1585 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.322f
C1586 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.DX_ D4 1.33e-19
C1587 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.DX_ 5_bit_dac_0[0].switch_n_3v3_0.D2 6.07e-19
C1588 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.482f
C1589 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.24f
C1590 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2.66e-20
C1591 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ D5 2.07e-19
C1592 switch_n_3v3_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 6.07e-19
C1593 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.229f
C1594 a_1556_12686# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0892f
C1595 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.00368f
C1596 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.00491f
C1597 5_bit_dac_0[1].4_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 1.05e-19
C1598 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.128f
C1599 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 0.00379f
C1600 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.13f
C1601 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.302f
C1602 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.DX_ D2_BUF 6.07e-19
C1603 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2.66e-20
C1604 VCC 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 0.779f
C1605 switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.0607f
C1606 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_11458# 0.00538f
C1607 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].switch_n_3v3_0.DX_ 1.79e-20
C1608 5_bit_dac_0[1].4_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.00107f
C1609 5_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 0.00197f
C1610 a_1556_17598# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2.93e-19
C1611 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5.55e-20
C1612 5_bit_dac_0[0].switch_n_3v3_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 6.07e-19
C1613 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].D0 0.544f
C1614 switch_n_3v3_0.D3 switch_n_3v3_0.D6 0.0625f
C1615 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 7.75e-19
C1616 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.00123f
C1617 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 VREFL 0.544f
C1618 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D6 1.72e-19
C1619 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00473f
C1620 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.38f
C1621 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5.19e-20
C1622 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00805f
C1623 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 1.26e-20
C1624 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[1].switch_n_3v3_0.D2 0.0155f
C1625 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.404f
C1626 5_bit_dac_0[1].4_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.544f
C1627 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH a_1556_11458# 0.175f
C1628 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 3.62e-20
C1629 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00805f
C1630 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 3.38e-20
C1631 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 4.97e-19
C1632 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL switch_n_3v3_0.D6 0.00202f
C1633 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.312f
C1634 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.347f
C1635 D4_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00517f
C1636 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5.89e-20
C1637 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 0.0858f
C1638 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 switch_n_3v3_0.D7 1.57e-20
C1639 5_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 4.97e-19
C1640 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH switch_n_3v3_0.D6 6.67e-19
C1641 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3.53e-19
C1642 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 8.92e-19
C1643 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH a_1556_16370# 9.57e-20
C1644 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 1.34e-20
C1645 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.00114f
C1646 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[1].switch_n_3v3_0.D3 4.43e-21
C1647 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.291f
C1648 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 0.552f
C1649 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.0551f
C1650 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00476f
C1651 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00394f
C1652 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].D0 4.97e-19
C1653 a_1556_9002# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0892f
C1654 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 4.97e-19
C1655 switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 3.08e-20
C1656 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.125f
C1657 5_bit_dac_0[1].4_bit_dac_0[1].VOUT 5_bit_dac_0[1].switch_n_3v3_0.D2 0.0034f
C1658 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 6.11e-19
C1659 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.111f
C1660 switch_n_3v3_0.D4 switch_n_3v3_0.D7 0.0925f
C1661 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 1.06f
C1662 5_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.0579f
C1663 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 1.34e-20
C1664 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.0923f
C1665 5_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.48e-19
C1666 VCC a_1556_10230# 0.713f
C1667 a_1556_4090# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 2.93e-19
C1668 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 switch_n_3v3_0.D6 0.0618f
C1669 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.635f
C1670 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH a_1556_4090# 9.57e-20
C1671 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 0.00262f
C1672 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT switch_n_3v3_0.D6 0.0258f
C1673 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H a_1556_6546# 0.397f
C1674 switch_n_3v3_0.D3 5_bit_dac_0[0].switch_n_3v3_0.D3 0.0618f
C1675 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 3.38e-20
C1676 switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.00594f
C1677 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.635f
C1678 D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.0255f
C1679 5_bit_dac_0[1].4_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 0.302f
C1680 5_bit_dac_0[1].4_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.0824f
C1681 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 3.38e-20
C1682 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 0.219f
C1683 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3.82e-19
C1684 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.00114f
C1685 D2 D3 0.398f
C1686 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.579f
C1687 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.045f
C1688 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00123f
C1689 a_1556_17598# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.00365f
C1690 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 a_1556_16370# 0.0981f
C1691 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.312f
C1692 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 4.15e-19
C1693 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.635f
C1694 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.00368f
C1695 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.00213f
C1696 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].VOUT 5.4e-19
C1697 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L a_1556_12686# 0.403f
C1698 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 0.044f
C1699 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.00819f
C1700 a_1556_4090# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0331f
C1701 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ D4 2.51e-19
C1702 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.312f
C1703 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].switch_n_3v3_0.DX_ 3.68e-19
C1704 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 3.47e-20
C1705 switch_n_3v3_0.D4 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 2.51e-19
C1706 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00123f
C1707 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.045f
C1708 5_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.DX_ 0.0139f
C1709 5_bit_dac_0[0].4_bit_dac_0[0].VOUT switch_n_3v3_0.D6 4.7e-20
C1710 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 2.38e-19
C1711 switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 1.03e-19
C1712 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 0.0026f
C1713 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L a_1556_5318# 1.29e-19
C1714 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.482f
C1715 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.00105f
C1716 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 6.14e-19
C1717 a_1556_7774# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 0.325f
C1718 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT switch_n_3v3_0.D6 0.0234f
C1719 switch_n_3v3_0.D4 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 2.52e-20
C1720 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.00832f
C1721 5_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 0.0104f
C1722 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.13f
C1723 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].D0 0.00379f
C1724 switch_n_3v3_0.D4 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.00147f
C1725 5_bit_dac_0[1].4_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.037f
C1726 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.00832f
C1727 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5.89e-20
C1728 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL D5 0.00306f
C1729 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.027f
C1730 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 1.18f
C1731 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 3.62e-20
C1732 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.0199f
C1733 5_bit_dac_0[1].switch_n_3v3_0.D3 D5 0.0849f
C1734 switch_n_3v3_0.D4 5_bit_dac_0[0].switch_n_3v3_0.D2 0.0361f
C1735 5_bit_dac_0[1].switch_n_3v3_0.DX_ switch_n_3v3_0.D7 0.0268f
C1736 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 0.0026f
C1737 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L a_1556_406# 1.29e-19
C1738 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].D0 2.29e-20
C1739 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.635f
C1740 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.0923f
C1741 switch_n_3v3_0.D3 switch_n_3v3_0.DX_ 1.03e-19
C1742 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.128f
C1743 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.0579f
C1744 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 2.34e-21
C1745 D5_BUF VOUT 0.0719f
C1746 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.DX_ D5 1.8e-19
C1747 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.312f
C1748 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.651f
C1749 5_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].VOUT 0.88f
C1750 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H VREFL 0.138f
C1751 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D2 0.00132f
C1752 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.836f
C1753 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 switch_n_3v3_0.D3 0.631f
C1754 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.0057f
C1755 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.579f
C1756 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_6546# 0.00538f
C1757 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.0211f
C1758 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 6.14e-19
C1759 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 0.00262f
C1760 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.00117f
C1761 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.00819f
C1762 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 1.06f
C1763 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.128f
C1764 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ D5_BUF 6.07e-19
C1765 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L a_1556_4090# 0.403f
C1766 VCC switch_n_3v3_0.D3 0.773f
C1767 D1 D3 2.93e-21
C1768 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.132f
C1769 5_bit_dac_0[0].4_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.0057f
C1770 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.714f
C1771 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[0].VOUT 2.04e-20
C1772 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0701f
C1773 switch_n_3v3_0.D3 5_bit_dac_0[0].VOUT 1.11e-21
C1774 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.00213f
C1775 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.0035f
C1776 VCC VREFH 0.0022f
C1777 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 9.82e-21
C1778 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.0222f
C1779 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.48e-19
C1780 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.0035f
C1781 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.312f
C1782 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 9.82e-21
C1783 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5.84e-19
C1784 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH a_1556_15142# 9.57e-20
C1785 a_1556_5318# 5_bit_dac_0[0].4_bit_dac_0[0].D1 6.04e-19
C1786 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[1].VOUT 2.82e-20
C1787 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.347f
C1788 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.622f
C1789 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 6.11e-19
C1790 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.111f
C1791 5_bit_dac_0[1].4_bit_dac_0[0].VOUT D5 4.14e-20
C1792 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 0.0744f
C1793 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.00117f
C1794 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.0035f
C1795 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.189f
C1796 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 9.82e-21
C1797 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.0035f
C1798 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.312f
C1799 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.651f
C1800 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.DX_ 3.53e-19
C1801 5_bit_dac_0[1].4_bit_dac_0[1].VOUT switch_n_3v3_0.D4 0.15f
C1802 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0102f
C1803 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H D0 0.117f
C1804 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 0.0988f
C1805 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0018f
C1806 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.48e-19
C1807 D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3.53e-19
C1808 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.482f
C1809 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.0104f
C1810 a_1556_7774# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0892f
C1811 VCC 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 0.779f
C1812 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.552f
C1813 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.00577f
C1814 D4_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 1.33e-19
C1815 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L a_1556_9002# 1.29e-19
C1816 a_1556_15142# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2.93e-19
C1817 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.579f
C1818 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.00183f
C1819 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0824f
C1820 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.482f
C1821 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 0.552f
C1822 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT switch_n_3v3_0.D6 0.0258f
C1823 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 9.82e-21
C1824 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.0035f
C1825 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH a_1556_5318# 9.57e-20
C1826 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 0.14f
C1827 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VOUT D5_BUF 1.79e-20
C1828 5_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3.36e-19
C1829 5_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 1.48e-19
C1830 5_bit_dac_0[1].4_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.48e-19
C1831 5_bit_dac_0[1].4_bit_dac_0[1].VREFH a_1556_12686# 1.97e-19
C1832 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 0.0988f
C1833 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 3.62e-20
C1834 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ D4_BUF 7.1e-20
C1835 VCC 5_bit_dac_0[0].4_bit_dac_0[0].VOUT 0.452f
C1836 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.24f
C1837 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.00114f
C1838 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.322f
C1839 5_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].VOUT 0.369f
C1840 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.189f
C1841 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL switch_n_3v3_0.D7 0.00143f
C1842 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].VOUT 0.252f
C1843 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.771f
C1844 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.00819f
C1845 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.0035f
C1846 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 1.06e-19
C1847 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 2.34e-21
C1848 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 0.00112f
C1849 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 2.51e-20
C1850 a_1556_13914# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 1.21e-20
C1851 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH a_1556_406# 9.57e-20
C1852 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.00183f
C1853 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.472f
C1854 5_bit_dac_0[1].4_bit_dac_0[1].VOUT 5_bit_dac_0[1].switch_n_3v3_0.DX_ 0.124f
C1855 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.115f
C1856 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.027f
C1857 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ D5 2.07e-19
C1858 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5.84e-19
C1859 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT D4_BUF 0.00505f
C1860 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VREFH a_1556_17598# 2.68e-20
C1861 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.229f
C1862 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.39f
C1863 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 6.14e-19
C1864 D3 switch_n_3v3_0.D7 0.0518f
C1865 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.315f
C1866 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D7 1.45e-19
C1867 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 switch_n_3v3_0.D6 1.79e-20
C1868 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH a_1556_4090# 0.175f
C1869 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 0.00112f
C1870 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].switch_n_3v3_0.D3 0.00505f
C1871 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.229f
C1872 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3.53e-19
C1873 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 0.00426f
C1874 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 1.81e-20
C1875 D4 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.0115f
C1876 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5.89e-20
C1877 VCC 5_bit_dac_0[0].4_bit_dac_0[0].D0 1.18f
C1878 5_bit_dac_0[0].switch_n_3v3_0.D3 switch_n_3v3_0.D6 0.0625f
C1879 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 1.9e-19
C1880 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D6 1.72e-19
C1881 a_1556_10230# 5_bit_dac_0[0].D1 6.04e-19
C1882 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 0.255f
C1883 5_bit_dac_0[0].4_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 2.66e-20
C1884 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].VREFH 0.0124f
C1885 D4_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.0259f
C1886 5_bit_dac_0[1].VOUT D5_BUF 0.15f
C1887 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 a_1556_11458# 0.003f
C1888 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 3.7e-20
C1889 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.48e-19
C1890 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0269f
C1891 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].D0 0.00164f
C1892 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.312f
C1893 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.00819f
C1894 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 6.14e-19
C1895 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.579f
C1896 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.115f
C1897 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.307f
C1898 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].switch_n_3v3_0.DX_ 1.79e-20
C1899 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 1.81e-20
C1900 a_1556_15142# a_1556_13914# 0.00981f
C1901 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.088f
C1902 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 0.24f
C1903 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 0.044f
C1904 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 1.7e-19
C1905 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.138f
C1906 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.DX_ 0.0904f
C1907 5_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.129f
C1908 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH switch_n_3v3_0.D7 5.14e-19
C1909 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 3.54e-19
C1910 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 0.0155f
C1911 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.00368f
C1912 a_1556_9002# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 6.04e-19
C1913 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.205f
C1914 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 8.92e-19
C1915 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.037f
C1916 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3.38e-20
C1917 5_bit_dac_0[1].4_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 2.66e-20
C1918 5_bit_dac_0[0].4_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0551f
C1919 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ switch_n_3v3_0.D6 2.54e-19
C1920 D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 2.96e-19
C1921 5_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00805f
C1922 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 3.54e-19
C1923 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 0.0988f
C1924 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 1.7e-19
C1925 D5 D5_BUF 0.0466f
C1926 a_1556_10230# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.0331f
C1927 D3_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00189f
C1928 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.0018f
C1929 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00143f
C1930 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D6 1.72e-19
C1931 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].switch_n_3v3_0.DX_ 0.00373f
C1932 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 0.0124f
C1933 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH D3 0.00189f
C1934 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.129f
C1935 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 9.68e-20
C1936 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.00368f
C1937 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH D5 8.21e-19
C1938 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].switch_n_3v3_0.D3 8.04e-20
C1939 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.205f
C1940 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[1].switch_n_3v3_0.D2 1.48e-19
C1941 5_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.00134f
C1942 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00143f
C1943 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 3.62e-20
C1944 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VOUT switch_n_3v3_0.D6 4.36e-20
C1945 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 0.219f
C1946 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.129f
C1947 5_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.0179f
C1948 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[0].VOUT 2.04e-20
C1949 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 1.8e-19
C1950 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 0.0124f
C1951 a_1556_17598# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0892f
C1952 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0018f
C1953 switch_n_3v3_0.DX_ switch_n_3v3_0.D6 2.54e-19
C1954 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.00319f
C1955 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.529f
C1956 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L D1 0.00319f
C1957 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0018f
C1958 D4_BUF D3_BUF 0.929f
C1959 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5.59e-19
C1960 D4_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 2.51e-19
C1961 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 switch_n_3v3_0.D6 0.0618f
C1962 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.0199f
C1963 5_bit_dac_0[1].4_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.DX_ 0.236f
C1964 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.00819f
C1965 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.DX_ 3.53e-19
C1966 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.39f
C1967 5_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.00489f
C1968 switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0145f
C1969 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.322f
C1970 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.00832f
C1971 switch_n_3v3_0.D4 VOUT 1.74e-20
C1972 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 1.18f
C1973 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.176f
C1974 a_1556_2862# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 6.04e-19
C1975 5_bit_dac_0[1].4_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.00183f
C1976 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].D0 0.472f
C1977 VCC switch_n_3v3_0.D6 0.823f
C1978 5_bit_dac_0[1].4_bit_dac_0[0].D1 D5 2.05e-20
C1979 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 6.14e-19
C1980 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.005f
C1981 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[0].switch_n_3v3_0.D3 6.07e-19
C1982 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0018f
C1983 5_bit_dac_0[0].VOUT switch_n_3v3_0.D6 2.25e-20
C1984 5_bit_dac_0[0].4_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.482f
C1985 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.314f
C1986 switch_n_3v3_0.D3 5_bit_dac_0[0].D1 3.54e-20
C1987 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0102f
C1988 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ switch_n_3v3_0.D7 0.0268f
C1989 switch_n_3v3_0.D4 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 1.33e-19
C1990 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.00123f
C1991 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00473f
C1992 a_1556_10230# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.296f
C1993 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT D5 0.0259f
C1994 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.504f
C1995 a_1556_7774# a_1556_6546# 0.00981f
C1996 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H a_1556_16370# 0.397f
C1997 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].D0 0.315f
C1998 5_bit_dac_0[1].4_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3.38e-20
C1999 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00805f
C2000 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].D0 0.0179f
C2001 a_1556_13914# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.296f
C2002 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].D1 4.15e-19
C2003 5_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].VOUT 1.22e-20
C2004 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.189f
C2005 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.472f
C2006 D4_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 4.04e-19
C2007 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.13f
C2008 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.125f
C2009 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 0.0026f
C2010 switch_n_3v3_0.D4 5_bit_dac_0[0].4_bit_dac_0[1].VOUT 2.76e-19
C2011 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.48e-19
C2012 D3 5_bit_dac_0[1].4_bit_dac_0[1].VOUT 6.19e-19
C2013 5_bit_dac_0[0].4_bit_dac_0[0].VOUT D2_BUF 1.79e-20
C2014 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.005f
C2015 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.0035f
C2016 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 1.34e-20
C2017 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 6.11e-19
C2018 5_bit_dac_0[1].4_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.111f
C2019 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.00114f
C2020 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 0.797f
C2021 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.DX_ 3.68e-19
C2022 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.291f
C2023 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.635f
C2024 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 0.14f
C2025 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.13f
C2026 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 0.00379f
C2027 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.0035f
C2028 a_1556_2862# a_1556_1634# 0.00981f
C2029 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 1.85e-19
C2030 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.0129f
C2031 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0102f
C2032 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0018f
C2033 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.48e-19
C2034 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.314f
C2035 VCC 5_bit_dac_0[0].switch_n_3v3_0.D3 0.773f
C2036 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.714f
C2037 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.68e-19
C2038 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.394f
C2039 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 1.9e-19
C2040 5_bit_dac_0[0].VOUT 5_bit_dac_0[0].switch_n_3v3_0.D3 3.76e-20
C2041 5_bit_dac_0[1].switch_n_3v3_0.D2 D5 0.0616f
C2042 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 0.0104f
C2043 a_1556_406# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0892f
C2044 a_1556_406# D1_BUF 6.04e-19
C2045 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 2.38e-19
C2046 VCC 5_bit_dac_0[1].4_bit_dac_0[0].D0 1.18f
C2047 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 0.00262f
C2048 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.14f
C2049 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.00123f
C2050 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00473f
C2051 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.00832f
C2052 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.836f
C2053 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.115f
C2054 switch_n_3v3_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 0.0104f
C2055 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.00349f
C2056 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L D0_BUF 1.9e-19
C2057 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.0102f
C2058 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.0107f
C2059 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 VREFH 0.0104f
C2060 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].D0 0.00379f
C2061 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.13f
C2062 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.00368f
C2063 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 2.34e-21
C2064 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.00164f
C2065 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 0.0104f
C2066 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].VOUT switch_n_3v3_0.D7 0.0133f
C2067 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 0.712f
C2068 switch_n_3v3_0.D4 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 2.45e-20
C2069 5_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.0222f
C2070 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH a_1556_12686# 9.57e-20
C2071 VREFL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.005f
C2072 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 1.81e-20
C2073 a_1556_15142# 5_bit_dac_0[1].4_bit_dac_0[0].D1 6.04e-19
C2074 5_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 0.0144f
C2075 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.00832f
C2076 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.303f
C2077 switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.0211f
C2078 5_bit_dac_0[0].switch_n_3v3_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 0.0104f
C2079 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.0179f
C2080 switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.0119f
C2081 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.714f
C2082 a_1556_12686# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 1.21e-20
C2083 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 2.51e-20
C2084 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D7 1.45e-19
C2085 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 1.46e-19
C2086 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.39f
C2087 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 2.38e-19
C2088 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 switch_n_3v3_0.D6 1.79e-20
C2089 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL D5 0.00306f
C2090 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00163f
C2091 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.511f
C2092 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 1.34e-20
C2093 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH switch_n_3v3_0.D7 4.71e-19
C2094 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.00183f
C2095 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.0107f
C2096 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].D1 1.85e-19
C2097 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L a_1556_406# 0.403f
C2098 a_1556_12686# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2.93e-19
C2099 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 0.523f
C2100 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.0211f
C2101 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.229f
C2102 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 1.81e-20
C2103 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3.36e-19
C2104 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H a_1556_9002# 0.397f
C2105 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.236f
C2106 switch_n_3v3_0.D4 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 2.69e-19
C2107 VCC switch_n_3v3_0.DX_ 0.712f
C2108 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 0.00262f
C2109 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 0.359f
C2110 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].VREFH 0.0104f
C2111 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH switch_n_3v3_0.D7 5.14e-19
C2112 switch_n_3v3_0.DX_ 5_bit_dac_0[0].VOUT 0.0853f
C2113 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH a_1556_10230# 9.57e-20
C2114 VCC 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 0.779f
C2115 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.0551f
C2116 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.236f
C2117 switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.017f
C2118 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.404f
C2119 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 3.23e-20
C2120 5_bit_dac_0[0].4_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.205f
C2121 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 1.46e-19
C2122 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.0923f
C2123 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.0579f
C2124 a_1556_11458# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.325f
C2125 D4_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00517f
C2126 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.177f
C2127 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.805f
C2128 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 9.82e-21
C2129 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5.55e-20
C2130 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL switch_n_3v3_0.D6 0.00202f
C2131 D4_BUF switch_n_3v3_0.D7 0.0406f
C2132 5_bit_dac_0[1].4_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 0.0353f
C2133 VCC 5_bit_dac_0[0].VOUT 0.614f
C2134 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT switch_n_3v3_0.D7 0.0324f
C2135 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH D4 0.00116f
C2136 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 0.359f
C2137 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L a_1556_17598# 1.29e-19
C2138 D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 9.68e-20
C2139 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH D1_BUF 3.54e-19
C2140 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5.89e-20
C2141 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.0261f
C2142 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0145f
C2143 a_1556_5318# a_1556_4090# 0.00981f
C2144 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ switch_n_3v3_0.D6 2.54e-19
C2145 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.0551f
C2146 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 4.97e-19
C2147 switch_n_3v3_0.D4 5_bit_dac_0[1].VOUT 0.0732f
C2148 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH switch_n_3v3_0.D7 5.14e-19
C2149 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT switch_n_3v3_0.D7 0.0397f
C2150 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.00368f
C2151 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 3.08e-20
C2152 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 switch_n_3v3_0.D7 1.57e-20
C2153 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.111f
C2154 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0927f
C2155 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 6.11e-19
C2156 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 1.06e-19
C2157 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.205f
C2158 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.00143f
C2159 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.DX_ switch_n_3v3_0.D6 2.54e-19
C2160 D2_BUF switch_n_3v3_0.D6 0.0293f
C2161 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 2.07e-19
C2162 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 1.46e-19
C2163 D2 D4 0.0322f
C2164 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5.55e-20
C2165 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.482f
C2166 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.DX_ 7.51e-19
C2167 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].switch_n_3v3_0.D2 0.00132f
C2168 5_bit_dac_0[1].4_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00805f
C2169 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.236f
C2170 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0018f
C2171 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.189f
C2172 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 6.14e-19
C2173 5_bit_dac_0[1].4_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.132f
C2174 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[0].D1 3.54e-20
C2175 D3_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 2.79e-20
C2176 5_bit_dac_0[1].4_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.482f
C2177 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.00105f
C2178 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.111f
C2179 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 6.11e-19
C2180 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.051f
C2181 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.005f
C2182 VCC VREFL 0.144f
C2183 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.0607f
C2184 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0018f
C2185 switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.0204f
C2186 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].D0 0.00379f
C2187 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.13f
C2188 switch_n_3v3_0.D4 D5 2.5f
C2189 5_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.005f
C2190 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.128f
C2191 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.697f
C2192 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.482f
C2193 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH D0_BUF 0.00105f
C2194 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_15142# 0.00538f
C2195 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.00143f
C2196 D4_BUF 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 2.09e-21
C2197 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.DX_ 7.51e-19
C2198 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.00832f
C2199 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.579f
C2200 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.005f
C2201 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0102f
C2202 D1_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.632f
C2203 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.005f
C2204 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.00164f
C2205 5_bit_dac_0[0].switch_n_3v3_0.D2 D4_BUF 0.0391f
C2206 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.115f
C2207 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.005f
C2208 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.176f
C2209 5_bit_dac_0[0].switch_n_3v3_0.DX_ switch_n_3v3_0.D7 0.0268f
C2210 5_bit_dac_0[1].VREFH a_1556_10230# 2.68e-20
C2211 switch_n_3v3_0.D4 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 1.33e-19
C2212 5_bit_dac_0[0].4_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 0.00231f
C2213 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.00114f
C2214 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3.36e-19
C2215 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.39f
C2216 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.00183f
C2217 switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 2.69e-19
C2218 5_bit_dac_0[1].4_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 0.45f
C2219 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH switch_n_3v3_0.D7 5.14e-19
C2220 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.13f
C2221 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 8.21e-19
C2222 switch_n_3v3_0.D4 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 2.51e-19
C2223 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3.53e-19
C2224 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 2.51e-20
C2225 a_1556_1634# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 1.21e-20
C2226 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 1.79e-20
C2227 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D7 1.45e-19
C2228 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ switch_n_3v3_0.D3 6.07e-19
C2229 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.836f
C2230 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.322f
C2231 5_bit_dac_0[1].switch_n_3v3_0.DX_ 5_bit_dac_0[1].VOUT 0.244f
C2232 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.303f
C2233 a_1556_4090# a_1556_2862# 0.00981f
C2234 5_bit_dac_0[0].D1 switch_n_3v3_0.D6 1.79e-20
C2235 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].D0 0.315f
C2236 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L a_1556_18826# 0.403f
C2237 5_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0701f
C2238 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.00577f
C2239 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.322f
C2240 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ D4 0.0056f
C2241 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.DX_ D3_BUF 0.219f
C2242 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].switch_n_3v3_0.D2 1.29f
C2243 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 7.75e-19
C2244 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[0].D1 2.05e-20
C2245 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.24f
C2246 5_bit_dac_0[1].4_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.00927f
C2247 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 0.797f
C2248 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.DX_ 1.79e-20
C2249 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 8.92e-19
C2250 D1 D4 1.41e-21
C2251 5_bit_dac_0[0].4_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.111f
C2252 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 6.11e-19
C2253 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L a_1556_16370# 1.29e-19
C2254 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00163f
C2255 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.511f
C2256 VCC D0 0.407f
C2257 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5.55e-20
C2258 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.0261f
C2259 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 1.81e-20
C2260 5_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.404f
C2261 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 D2 0.0026f
C2262 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H a_1556_12686# 0.397f
C2263 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 1.18f
C2264 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.0102f
C2265 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH switch_n_3v3_0.D7 4.71e-19
C2266 a_1556_7774# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2.93e-19
C2267 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.236f
C2268 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 2.29e-20
C2269 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.189f
C2270 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.132f
C2271 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].D1 0.044f
C2272 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 0.255f
C2273 5_bit_dac_0[1].switch_n_3v3_0.DX_ D5 1.8e-19
C2274 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.138f
C2275 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L a_1556_7774# 0.403f
C2276 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].D1 3.54e-19
C2277 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.0104f
C2278 5_bit_dac_0[0].switch_n_3v3_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 9.82e-21
C2279 a_1556_11458# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0331f
C2280 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.DX_ 0.0104f
C2281 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3.36e-19
C2282 a_1556_16370# 5_bit_dac_0[1].4_bit_dac_0[0].D0 0.00365f
C2283 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 a_1556_15142# 0.0981f
C2284 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 1.81e-20
C2285 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.312f
C2286 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.00368f
C2287 5_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.544f
C2288 5_bit_dac_0[1].4_bit_dac_0[0].D1 a_1556_13914# 0.003f
C2289 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].VOUT 0.00174f
C2290 a_1556_16370# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0331f
C2291 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.68e-19
C2292 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 1.7e-19
C2293 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.DX_ 0.125f
C2294 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.0018f
C2295 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL D3 0.0269f
C2296 5_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].switch_n_3v3_0.DX_ 3.53e-19
C2297 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.132f
C2298 switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.0295f
C2299 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.291f
C2300 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH switch_n_3v3_0.D7 5.14e-19
C2301 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0269f
C2302 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.00117f
C2303 5_bit_dac_0[1].4_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.00262f
C2304 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D6 1.72e-19
C2305 5_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].VOUT 6.06e-19
C2306 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 8.21e-19
C2307 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 0.712f
C2308 a_1556_1634# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0331f
C2309 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5.84e-19
C2310 D0 VREFL 0.77f
C2311 5_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.13f
C2312 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.514f
C2313 VCC D2_BUF 0.337f
C2314 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].VOUT switch_n_3v3_0.D7 0.0133f
C2315 VCC 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.DX_ 0.712f
C2316 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].VOUT 0.00119f
C2317 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2.66e-20
C2318 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.00692f
C2319 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2.38e-19
C2320 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 2.51e-20
C2321 a_1556_16370# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 1.21e-20
C2322 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 7.75e-19
C2323 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 2.96e-19
C2324 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.00123f
C2325 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00473f
C2326 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL switch_n_3v3_0.D6 0.00202f
C2327 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.472f
C2328 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.00183f
C2329 5_bit_dac_0[0].4_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 9.68e-20
C2330 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.302f
C2331 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.045f
C2332 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00123f
C2333 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH D1_BUF 1.85e-19
C2334 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.0551f
C2335 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.265f
C2336 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 1.9e-19
C2337 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_7774# 0.00538f
C2338 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL switch_n_3v3_0.D6 0.00202f
C2339 5_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00872f
C2340 a_1556_5318# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.296f
C2341 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 D3 4.81e-19
C2342 D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 0.0384f
C2343 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.037f
C2344 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 4.25e-19
C2345 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 4.15e-19
C2346 VREFL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 2.66e-20
C2347 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.511f
C2348 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 4.97e-19
C2349 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0018f
C2350 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 switch_n_3v3_0.D7 1.57e-20
C2351 D4_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 7.43e-20
C2352 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.051f
C2353 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 0.0124f
C2354 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.302f
C2355 a_1556_6546# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0331f
C2356 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.115f
C2357 VCC a_1556_16370# 0.713f
C2358 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 a_1556_7774# 0.0981f
C2359 a_1556_9002# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 0.00365f
C2360 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.00164f
C2361 5_bit_dac_0[0].D1 switch_n_3v3_0.DX_ 1.34e-20
C2362 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 0.00375f
C2363 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL switch_n_3v3_0.D6 0.00202f
C2364 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 switch_n_3v3_0.D6 0.0618f
C2365 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH switch_n_3v3_0.D6 6.1e-19
C2366 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 2.07e-19
C2367 switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.249f
C2368 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.0035f
C2369 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.394f
C2370 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00805f
C2371 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5.89e-20
C2372 D4 switch_n_3v3_0.D7 0.0519f
C2373 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.404f
C2374 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 3.8e-20
C2375 5_bit_dac_0[0].4_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2.38e-19
C2376 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.00832f
C2377 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 2.05e-20
C2378 VCC 5_bit_dac_0[0].D1 0.797f
C2379 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.303f
C2380 switch_n_3v3_0.D4 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00517f
C2381 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.176f
C2382 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 5_bit_dac_0[0].switch_n_3v3_0.D2 0.0719f
C2383 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 6.11e-19
C2384 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.111f
C2385 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H a_1556_9002# 4.83e-19
C2386 5_bit_dac_0[1].switch_n_3v3_0.D3 switch_n_3v3_0.D4 1.25f
C2387 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 0.0744f
C2388 D0_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.347f
C2389 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.00577f
C2390 5_bit_dac_0[0].4_bit_dac_0[1].VREFH a_1556_5318# 2.68e-20
C2391 D0_BUF D1_BUF 0.00262f
C2392 switch_n_3v3_0.D4 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.DX_ 1.33e-19
C2393 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00394f
C2394 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 1.7e-19
C2395 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0801f
C2396 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.0104f
C2397 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 0.315f
C2398 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 1.06e-19
C2399 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.DX_ switch_n_3v3_0.D7 0.0268f
C2400 5_bit_dac_0[0].4_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.132f
C2401 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.205f
C2402 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VOUT switch_n_3v3_0.D7 0.0191f
C2403 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 D1 0.0179f
C2404 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.805f
C2405 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 0.0124f
C2406 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 a_1556_6546# 0.003f
C2407 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 1.34e-20
C2408 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 0.628f
C2409 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.0204f
C2410 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.128f
C2411 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 6.14e-19
C2412 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.836f
C2413 D3 D5 0.0324f
C2414 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 3.62e-20
C2415 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ D5 2.07e-19
C2416 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 0.00237f
C2417 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.312f
C2418 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.514f
C2419 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL switch_n_3v3_0.D6 0.00202f
C2420 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.0923f
C2421 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.0579f
C2422 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 2.66e-20
C2423 5_bit_dac_0[1].4_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3.36e-19
C2424 switch_n_3v3_0.D4 5_bit_dac_0[1].4_bit_dac_0[0].VOUT 0.177f
C2425 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5.55e-20
C2426 switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 0.0694f
C2427 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 1.17f
C2428 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 4.25e-19
C2429 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.714f
C2430 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.DX_ 1.8e-19
C2431 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0102f
C2432 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.00805f
C2433 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 a_1556_1634# 0.003f
C2434 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH a_1556_17598# 0.175f
C2435 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L D0_BUF 0.315f
C2436 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH D4 0.00116f
C2437 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3.53e-19
C2438 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT switch_n_3v3_0.D6 0.027f
C2439 D4_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.0271f
C2440 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 0.544f
C2441 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00394f
C2442 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 switch_n_3v3_0.D7 1.57e-20
C2443 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 0.00349f
C2444 switch_n_3v3_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00394f
C2445 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 1.06f
C2446 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.312f
C2447 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].switch_n_3v3_0.DX_ 1.03e-19
C2448 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL switch_n_3v3_0.D6 0.00202f
C2449 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 1.7e-19
C2450 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H a_1556_5318# 0.397f
C2451 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.291f
C2452 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ switch_n_3v3_0.D6 2.54e-19
C2453 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 4.15e-19
C2454 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.DX_ 0.0104f
C2455 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH D5 8.97e-19
C2456 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.236f
C2457 switch_n_3v3_0.D4 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00116f
C2458 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VREFH a_1556_15142# 1.97e-19
C2459 5_bit_dac_0[0].4_bit_dac_0[1].VREFH a_1556_2862# 1.97e-19
C2460 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.312f
C2461 VCC a_1556_12686# 0.713f
C2462 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 D4 2.52e-20
C2463 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].VOUT 3.47e-20
C2464 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 0.132f
C2465 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 0.00349f
C2466 switch_n_3v3_0.D4 5_bit_dac_0[0].4_bit_dac_0[0].D1 4.72e-19
C2467 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5.59e-19
C2468 a_1556_17598# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 0.325f
C2469 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.805f
C2470 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 0.00375f
C2471 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 0.0124f
C2472 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00476f
C2473 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_16370# 0.00538f
C2474 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL switch_n_3v3_0.D6 0.00202f
C2475 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5.55e-20
C2476 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[1].VOUT 1.47e-19
C2477 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 a_1556_17598# 0.003f
C2478 5_bit_dac_0[0].4_bit_dac_0[1].VOUT D4_BUF 0.15f
C2479 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 switch_n_3v3_0.D3 4.43e-21
C2480 5_bit_dac_0[0].4_bit_dac_0[0].D1 a_1556_4090# 0.003f
C2481 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 0.219f
C2482 5_bit_dac_0[0].4_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 1.05e-19
C2483 5_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].D1 0.0189f
C2484 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VREFH a_1556_2862# 2.68e-20
C2485 VCC 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 0.776f
C2486 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.622f
C2487 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.312f
C2488 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.205f
C2489 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.189f
C2490 5_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 1.79e-20
C2491 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.249f
C2492 5_bit_dac_0[1].4_bit_dac_0[1].VOUT D4 2.76e-19
C2493 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.349f
C2494 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.0035f
C2495 5_bit_dac_0[1].switch_n_3v3_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].VOUT 0.0853f
C2496 5_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 2.96e-19
C2497 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.0261f
C2498 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.176f
C2499 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 8.92e-19
C2500 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00805f
C2501 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0269f
C2502 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 3.82e-19
C2503 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 0.00164f
C2504 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.48e-19
C2505 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 7.75e-19
C2506 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.0018f
C2507 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT switch_n_3v3_0.D6 0.027f
C2508 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.504f
C2509 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.176f
C2510 a_1556_18826# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0331f
C2511 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00805f
C2512 5_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.00319f
C2513 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT switch_n_3v3_0.D7 0.0397f
C2514 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].VOUT 2.49e-22
C2515 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 0.00237f
C2516 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.394f
C2517 switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0701f
C2518 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 switch_n_3v3_0.D7 1.57e-20
C2519 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ D5 1.8e-19
C2520 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.39f
C2521 switch_n_3v3_0.D4 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00116f
C2522 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.394f
C2523 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H D1 0.037f
C2524 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 1.06f
C2525 switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 2.78e-19
C2526 a_1556_13914# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0331f
C2527 5_bit_dac_0[1].4_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 3.96e-20
C2528 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0801f
C2529 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.291f
C2530 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.0018f
C2531 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 D1_BUF 0.0392f
C2532 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.051f
C2533 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].D0 0.315f
C2534 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].D1 4.15e-19
C2535 5_bit_dac_0[1].4_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.0579f
C2536 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.0923f
C2537 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 0.0104f
C2538 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.68e-19
C2539 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00872f
C2540 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00473f
C2541 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.00114f
C2542 a_1556_6546# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.325f
C2543 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.129f
C2544 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 3.7e-20
C2545 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].VOUT 0.0157f
C2546 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.00491f
C2547 5_bit_dac_0[1].4_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.38f
C2548 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.302f
C2549 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.312f
C2550 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].D0 0.24f
C2551 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.322f
C2552 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.00319f
C2553 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 switch_n_3v3_0.D7 0.0916f
C2554 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.0579f
C2555 5_bit_dac_0[0].4_bit_dac_0[1].VOUT 5_bit_dac_0[0].switch_n_3v3_0.DX_ 0.124f
C2556 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.0923f
C2557 a_1556_18826# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 0.00365f
C2558 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 2.05e-20
C2559 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 a_1556_17598# 0.0981f
C2560 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 5_bit_dac_0[1].VOUT 0.00366f
C2561 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 1.06e-19
C2562 D2 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 0.0694f
C2563 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 0.00112f
C2564 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.128f
C2565 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].VREFH 0.0988f
C2566 a_1556_18826# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 6.04e-19
C2567 5_bit_dac_0[0].4_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5.84e-19
C2568 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].VREFH 0.0988f
C2569 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.312f
C2570 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 0.0757f
C2571 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 a_1556_12686# 0.0981f
C2572 a_1556_13914# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 0.00365f
C2573 switch_n_3v3_0.D3 switch_n_3v3_0.D2 1.29f
C2574 5_bit_dac_0[0].4_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.00927f
C2575 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.836f
C2576 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.00368f
C2577 D3_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 2.09e-21
C2578 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT switch_n_3v3_0.D6 0.027f
C2579 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.774f
C2580 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0927f
C2581 D4_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.233f
C2582 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 0.219f
C2583 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0102f
C2584 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 1.85e-19
C2585 switch_n_3v3_0.D4 D5_BUF 2.51f
C2586 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.322f
C2587 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.00319f
C2588 5_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.00406f
C2589 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.0172f
C2590 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL switch_n_3v3_0.D7 0.00143f
C2591 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.312f
C2592 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.347f
C2593 switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0668f
C2594 D3 5_bit_dac_0[1].switch_n_3v3_0.D3 0.0618f
C2595 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 0.712f
C2596 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.DX_ 1.79e-20
C2597 switch_n_3v3_0.D4 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00116f
C2598 5_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 0.0026f
C2599 5_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0668f
C2600 5_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.347f
C2601 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 4.15e-19
C2602 switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.0265f
C2603 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.125f
C2604 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 0.00132f
C2605 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].D0 2.29e-20
C2606 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].VOUT D5 3.8e-20
C2607 a_1556_4090# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 1.21e-20
C2608 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.291f
C2609 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 2.51e-20
C2610 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.347f
C2611 D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.134f
C2612 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H a_1556_2862# 0.397f
C2613 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 a_1556_10230# 0.0981f
C2614 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 1.06f
C2615 D2_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0668f
C2616 a_1556_11458# 5_bit_dac_0[0].D0 0.00365f
C2617 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.051f
C2618 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.00368f
C2619 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 1.18f
C2620 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.0757f
C2621 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 0.0189f
C2622 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.0757f
C2623 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.312f
C2624 5_bit_dac_0[1].4_bit_dac_0[0].D1 switch_n_3v3_0.D4 2.7e-21
C2625 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ switch_n_3v3_0.D6 2.54e-19
C2626 VREFL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 3.7e-20
C2627 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 2.78e-22
C2628 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[0].switch_n_3v3_0.D2 0.0694f
C2629 switch_n_3v3_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.0199f
C2630 5_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.0404f
C2631 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.229f
C2632 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.00319f
C2633 switch_n_3v3_0.D4 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.0259f
C2634 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 2.09e-21
C2635 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.0757f
C2636 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 1.79e-20
C2637 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 0.00237f
C2638 D1 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 1.48e-19
C2639 5_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.00491f
C2640 D5 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0011f
C2641 5_bit_dac_0[0].4_bit_dac_0[0].VOUT D3_BUF 0.0719f
C2642 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00805f
C2643 a_1556_18826# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.325f
C2644 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.511f
C2645 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00163f
C2646 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.771f
C2647 5_bit_dac_0[0].4_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 0.45f
C2648 5_bit_dac_0[1].4_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.0745f
C2649 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.0579f
C2650 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.0923f
C2651 5_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.123f
C2652 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH a_1556_406# 0.175f
C2653 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5.55e-20
C2654 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL switch_n_3v3_0.D7 0.00143f
C2655 5_bit_dac_0[0].switch_n_3v3_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.0143f
C2656 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D6 1.72e-19
C2657 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 D2_BUF 0.0694f
C2658 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.00114f
C2659 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 2.51e-20
C2660 a_1556_7774# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 1.21e-20
C2661 5_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0668f
C2662 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT D5 0.0259f
C2663 switch_n_3v3_0.D4 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.DX_ 1.33e-19
C2664 5_bit_dac_0[0].4_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.635f
C2665 VCC 5_bit_dac_0[1].VREFH 0.14f
C2666 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 2.38e-19
C2667 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH a_1556_2862# 0.337f
C2668 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT D5 0.027f
C2669 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L a_1556_11458# 0.403f
C2670 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 D5 2.05e-20
C2671 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.394f
C2672 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ D4_BUF 6.07e-19
C2673 5_bit_dac_0[0].4_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 0.0174f
C2674 5_bit_dac_0[1].switch_n_3v3_0.D2 switch_n_3v3_0.D4 0.0391f
C2675 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.0757f
C2676 D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.48e-19
C2677 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H a_1556_17598# 4.83e-19
C2678 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT switch_n_3v3_0.D6 0.0258f
C2679 D4_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.02f
C2680 D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.0057f
C2681 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.0018f
C2682 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 1.9e-19
C2683 5_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.635f
C2684 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.005f
C2685 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.0199f
C2686 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.514f
C2687 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 2.34e-21
C2688 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.128f
C2689 5_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5.84e-19
C2690 5_bit_dac_0[1].4_bit_dac_0[0].D1 5_bit_dac_0[1].switch_n_3v3_0.DX_ 1.34e-20
C2691 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3.36e-19
C2692 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT switch_n_3v3_0.DX_ 3.68e-19
C2693 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.229f
C2694 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 3.74e-19
C2695 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5.59e-19
C2696 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 0.219f
C2697 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.14f
C2698 switch_n_3v3_0.D3 switch_n_3v3_0.D7 0.0924f
C2699 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 4.58e-19
C2700 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D7 1.45e-19
C2701 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 2.29e-20
C2702 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 4.15e-19
C2703 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 switch_n_3v3_0.D6 1.79e-20
C2704 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.394f
C2705 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.115f
C2706 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3.53e-19
C2707 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.38f
C2708 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH switch_n_3v3_0.D6 6.1e-19
C2709 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT switch_n_3v3_0.D6 0.0258f
C2710 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.771f
C2711 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 1.9e-19
C2712 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.38f
C2713 5_bit_dac_0[1].4_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.265f
C2714 5_bit_dac_0[0].4_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].D1 1.7e-19
C2715 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.00832f
C2716 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].VOUT 0.00112f
C2717 5_bit_dac_0[1].4_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.138f
C2718 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.579f
C2719 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL switch_n_3v3_0.D7 0.00143f
C2720 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5.84e-19
C2721 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ D3 0.00213f
C2722 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT D0_BUF 2.29e-20
C2723 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 0.00375f
C2724 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.0172f
C2725 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH switch_n_3v3_0.D7 5.14e-19
C2726 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.00368f
C2727 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 3.68e-19
C2728 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 0.24f
C2729 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.0102f
C2730 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH D5 8.97e-19
C2731 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.00349f
C2732 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.205f
C2733 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.38f
C2734 D2 switch_n_3v3_0.D6 0.0325f
C2735 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.0265f
C2736 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.463f
C2737 VCC a_1556_7774# 0.713f
C2738 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 2.29e-20
C2739 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ D5 0.00535f
C2740 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0551f
C2741 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 3.7e-20
C2742 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[0].switch_n_3v3_0.DX_ 0.0104f
C2743 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 3.7e-20
C2744 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 0.044f
C2745 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL D4 0.00517f
C2746 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VOUT switch_n_3v3_0.D6 4.36e-20
C2747 switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.00213f
C2748 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH a_1556_10230# 0.175f
C2749 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.236f
C2750 5_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].switch_n_3v3_0.DX_ 3.53e-19
C2751 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.68e-19
C2752 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.00368f
C2753 5_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0551f
C2754 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 switch_n_3v3_0.D7 0.0916f
C2755 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT switch_n_3v3_0.D7 0.0324f
C2756 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.00143f
C2757 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 0.698f
C2758 switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 4.81e-19
C2759 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 8.92e-19
C2760 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.0607f
C2761 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H a_1556_18826# 0.397f
C2762 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.00832f
C2763 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.00143f
C2764 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00306f
C2765 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.68e-19
C2766 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.805f
C2767 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0102f
C2768 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 7.75e-19
C2769 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5.84e-19
C2770 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 0.177f
C2771 D3_BUF switch_n_3v3_0.D6 0.0299f
C2772 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].D0 0.00164f
C2773 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.38f
C2774 a_1556_17598# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 4.09e-19
C2775 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.205f
C2776 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H a_1556_16370# 4.83e-19
C2777 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D6 1.72e-19
C2778 switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 2.96e-19
C2779 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.291f
C2780 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 0.544f
C2781 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 D4 2.52e-20
C2782 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 9.68e-20
C2783 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].D1 0.00237f
C2784 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.714f
C2785 5_bit_dac_0[0].4_bit_dac_0[0].VOUT switch_n_3v3_0.D7 0.00725f
C2786 switch_n_3v3_0.D4 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 2.52e-20
C2787 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 1.9e-19
C2788 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.265f
C2789 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.322f
C2790 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0701f
C2791 switch_n_3v3_0.D2 switch_n_3v3_0.D6 0.0618f
C2792 a_1556_6546# a_1556_5318# 0.00981f
C2793 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH D5 8.97e-19
C2794 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VREFH a_1556_11458# 0.337f
C2795 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.0551f
C2796 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.0018f
C2797 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT switch_n_3v3_0.D7 0.036f
C2798 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D6 1.72e-19
C2799 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 5_bit_dac_0[0].switch_n_3v3_0.D3 0.15f
C2800 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 0.359f
C2801 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 3.62e-20
C2802 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0927f
C2803 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L a_1556_15142# 1.29e-19
C2804 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.0261f
C2805 5_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.482f
C2806 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.00105f
C2807 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0927f
C2808 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ switch_n_3v3_0.D6 2.54e-19
C2809 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 0.00375f
C2810 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT switch_n_3v3_0.D6 0.0258f
C2811 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 1.9e-19
C2812 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.265f
C2813 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.552f
C2814 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 0.00349f
C2815 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 0.0988f
C2816 D4_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 2.38e-20
C2817 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.394f
C2818 5_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.0181f
C2819 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00476f
C2820 a_1556_1634# a_1556_406# 0.00981f
C2821 a_1556_16370# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 2.93e-19
C2822 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 3.62e-20
C2823 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 1.46e-19
C2824 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.DX_ 3.68e-19
C2825 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH a_1556_7774# 0.175f
C2826 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.635f
C2827 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0927f
C2828 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 4.25e-19
C2829 5_bit_dac_0[0].switch_n_3v3_0.D3 D3_BUF 0.0618f
C2830 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.00368f
C2831 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 0.236f
C2832 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 switch_n_3v3_0.D2 0.0155f
C2833 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.00594f
C2834 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 0.0189f
C2835 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3.36e-19
C2836 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].switch_n_3v3_0.D3 0.00505f
C2837 D4 5_bit_dac_0[1].VOUT 2.07e-20
C2838 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 0.255f
C2839 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.303f
C2840 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].D0 0.472f
C2841 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 0.00237f
C2842 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.0923f
C2843 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.0579f
C2844 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.635f
C2845 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 0.797f
C2846 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.13f
C2847 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.0295f
C2848 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.00379f
C2849 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 3.38e-20
C2850 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.529f
C2851 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 1.06e-19
C2852 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.622f
C2853 D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 1.75e-20
C2854 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 3.11e-20
C2855 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.0018f
C2856 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0102f
C2857 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].VOUT 2.78e-22
C2858 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 3.62e-20
C2859 5_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 3.12e-19
C2860 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.00692f
C2861 D4_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 2.51e-19
C2862 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.DX_ 3.68e-19
C2863 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 0.0026f
C2864 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.00692f
C2865 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 0.00262f
C2866 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.00819f
C2867 5_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[0].VOUT 6.06e-19
C2868 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.005f
C2869 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 1.03e-19
C2870 5_bit_dac_0[1].4_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5.84e-19
C2871 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 0.044f
C2872 switch_n_3v3_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 5.19e-19
C2873 VOUT 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 1.79e-20
C2874 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.514f
C2875 5_bit_dac_0[0].4_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 1.9e-19
C2876 VCC D2 0.333f
C2877 5_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 0.0867f
C2878 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5.89e-20
C2879 5_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.0057f
C2880 a_1556_12686# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.296f
C2881 D4 D5 2.27f
C2882 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 1.7e-19
C2883 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0927f
C2884 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.00692f
C2885 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.0018f
C2886 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L a_1556_7774# 1.29e-19
C2887 switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 0.0904f
C2888 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 0.523f
C2889 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[1].VOUT 6.12e-19
C2890 5_bit_dac_0[1].switch_n_3v3_0.DX_ switch_n_3v3_0.D4 0.219f
C2891 5_bit_dac_0[1].4_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.0295f
C2892 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.48e-19
C2893 a_1556_15142# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0892f
C2894 5_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 0.0534f
C2895 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VREFH a_1556_6546# 0.337f
C2896 5_bit_dac_0[1].VREFH 5_bit_dac_0[0].D1 1.7e-19
C2897 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].D1 6.11e-19
C2898 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.111f
C2899 5_bit_dac_0[0].switch_n_3v3_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 4.09e-19
C2900 5_bit_dac_0[1].4_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.213f
C2901 a_1556_12686# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.0331f
C2902 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.39f
C2903 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.315f
C2904 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.404f
C2905 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].VOUT 6.12e-19
C2906 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.0104f
C2907 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00163f
C2908 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 0.00164f
C2909 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.511f
C2910 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.38f
C2911 a_1556_10230# a_1556_9002# 0.00981f
C2912 5_bit_dac_0[0].4_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.347f
C2913 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH a_1556_1634# 2.68e-20
C2914 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VOUT D5 3.23e-20
C2915 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.00213f
C2916 VCC D3_BUF 0.396f
C2917 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 2.34e-21
C2918 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.0824f
C2919 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT switch_n_3v3_0.D7 0.0324f
C2920 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.714f
C2921 switch_n_3v3_0.D2 switch_n_3v3_0.DX_ 3.53e-19
C2922 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VREFH a_1556_1634# 0.337f
C2923 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.38f
C2924 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 9.82e-21
C2925 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.00692f
C2926 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL switch_n_3v3_0.D6 0.00202f
C2927 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 switch_n_3v3_0.D2 0.0694f
C2928 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5.55e-20
C2929 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5.59e-19
C2930 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 1.9e-19
C2931 5_bit_dac_0[0].4_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.265f
C2932 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ D2_BUF 0.219f
C2933 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 3.82e-19
C2934 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.045f
C2935 switch_n_3v3_0.D6 switch_n_3v3_0.D7 9.44f
C2936 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00123f
C2937 5_bit_dac_0[0].4_bit_dac_0[0].D1 D4_BUF 2.7e-21
C2938 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5.55e-20
C2939 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].VOUT 0.0157f
C2940 VCC switch_n_3v3_0.D2 0.779f
C2941 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 4.25e-19
C2942 5_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.205f
C2943 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0668f
C2944 switch_n_3v3_0.D2 5_bit_dac_0[0].VOUT 5.38e-19
C2945 a_1556_9002# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.296f
C2946 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT switch_n_3v3_0.DX_ 7.51e-19
C2947 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.714f
C2948 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 9.82e-21
C2949 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.0824f
C2950 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 0.00237f
C2951 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.0057f
C2952 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].D1 1.81e-20
C2953 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 2.96e-19
C2954 a_1556_13914# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 6.04e-19
C2955 VCC D1 0.459f
C2956 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH a_1556_13914# 2.68e-20
C2957 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 0.712f
C2958 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.39f
C2959 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 0.472f
C2960 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.533f
C2961 5_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 0.00149f
C2962 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5.89e-20
C2963 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 D5 2.05e-20
C2964 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 0.00262f
C2965 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.00819f
C2966 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.291f
C2967 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.0035f
C2968 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].VOUT 0.0065f
C2969 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 1.06f
C2970 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.0757f
C2971 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH D0_BUF 0.472f
C2972 VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 7.62e-19
C2973 a_1556_9002# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.325f
C2974 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.045f
C2975 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00123f
C2976 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 switch_n_3v3_0.D7 1.57e-20
C2977 a_1556_1634# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 2.93e-19
C2978 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.511f
C2979 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00163f
C2980 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D6 1.72e-19
C2981 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.0035f
C2982 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.482f
C2983 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 0.0757f
C2984 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 0.00105f
C2985 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.544f
C2986 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.00193f
C2987 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.017f
C2988 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.00183f
C2989 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 0.472f
C2990 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 1.06f
C2991 5_bit_dac_0[0].switch_n_3v3_0.D3 switch_n_3v3_0.D7 0.0924f
C2992 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 0.00375f
C2993 5_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3.38e-20
C2994 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D7 1.45e-19
C2995 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 switch_n_3v3_0.D6 1.79e-20
C2996 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00163f
C2997 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.511f
C2998 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH switch_n_3v3_0.D6 6.67e-19
C2999 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.0551f
C3000 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.0102f
C3001 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].VOUT 7.93e-20
C3002 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.68e-19
C3003 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 0.00237f
C3004 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00473f
C3005 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.00123f
C3006 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH switch_n_3v3_0.D6 6.1e-19
C3007 D1 VREFL 1.7e-19
C3008 5_bit_dac_0[0].switch_n_3v3_0.D2 switch_n_3v3_0.D6 0.0618f
C3009 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 2.07e-19
C3010 switch_n_3v3_0.D4 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.0115f
C3011 5_bit_dac_0[0].4_bit_dac_0[0].D1 5_bit_dac_0[0].switch_n_3v3_0.DX_ 1.34e-20
C3012 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 1.9e-19
C3013 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.265f
C3014 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[1].switch_n_3v3_0.D2 0.219f
C3015 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L a_1556_17598# 0.403f
C3016 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH a_1556_7774# 9.57e-20
C3017 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 8.21e-19
C3018 a_1556_7774# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 4.09e-19
C3019 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H a_1556_6546# 4.83e-19
C3020 5_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 2.66e-20
C3021 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ switch_n_3v3_0.D7 0.0268f
C3022 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL a_1556_4090# 0.00538f
C3023 switch_n_3v3_0.D3 VOUT 1.45e-20
C3024 D5_BUF 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 2.09e-21
C3025 D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 0.0904f
C3026 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.0104f
C3027 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3.82e-19
C3028 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].VOUT 2.78e-22
C3029 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.115f
C3030 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.00114f
C3031 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT D5 0.027f
C3032 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D7 1.45e-19
C3033 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 switch_n_3v3_0.D6 1.79e-20
C3034 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0801f
C3035 switch_n_3v3_0.D4 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 2.51e-19
C3036 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.00123f
C3037 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00473f
C3038 switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 3.74e-19
C3039 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H a_1556_1634# 4.83e-19
C3040 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL a_1556_5318# 0.00538f
C3041 a_1556_2862# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 4.09e-19
C3042 D5_BUF D4_BUF 2.18f
C3043 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[0].switch_n_3v3_0.D3 4.43e-21
C3044 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 0.219f
C3045 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].D0 0.132f
C3046 5_bit_dac_0[0].4_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0801f
C3047 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.00193f
C3048 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VOUT switch_n_3v3_0.D7 0.0191f
C3049 D4_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 2.51e-19
C3050 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00394f
C3051 switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[1].VOUT 6.19e-19
C3052 switch_n_3v3_0.DX_ switch_n_3v3_0.D7 0.0268f
C3053 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 0.219f
C3054 5_bit_dac_0[0].4_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.0824f
C3055 a_1556_11458# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0892f
C3056 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 a_1556_2862# 0.003f
C3057 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00394f
C3058 5_bit_dac_0[1].switch_n_3v3_0.D3 D4 1.25f
C3059 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 8.97e-19
C3060 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 3.54e-19
C3061 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].switch_n_3v3_0.D2 1.29f
C3062 D4_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 2.45e-20
C3063 a_1556_16370# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0892f
C3064 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 switch_n_3v3_0.D7 0.0916f
C3065 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 1.18f
C3066 D4_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 2.52e-20
C3067 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.394f
C3068 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.472f
C3069 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.38f
C3070 5_bit_dac_0[1].4_bit_dac_0[1].VOUT switch_n_3v3_0.D6 4.1e-20
C3071 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.312f
C3072 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 1.79e-20
C3073 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H D1_BUF 0.00237f
C3074 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.836f
C3075 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.00164f
C3076 5_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 9.68e-20
C3077 VCC switch_n_3v3_0.D7 2.1f
C3078 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].D0 0.24f
C3079 5_bit_dac_0[1].4_bit_dac_0[1].VREFH a_1556_15142# 2.68e-20
C3080 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00143f
C3081 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 3.53e-19
C3082 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.39f
C3083 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.DX_ 0.125f
C3084 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH a_1556_6546# 1.97e-19
C3085 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00394f
C3086 5_bit_dac_0[0].VOUT switch_n_3v3_0.D7 0.00551f
C3087 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 0.143f
C3088 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.0824f
C3089 a_1556_1634# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0892f
C3090 5_bit_dac_0[0].4_bit_dac_0[1].VREFH a_1556_4090# 0.337f
C3091 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L a_1556_6546# 0.403f
C3092 D3_BUF D2_BUF 0.307f
C3093 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.836f
C3094 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.189f
C3095 a_1556_10230# 5_bit_dac_0[0].D0 0.325f
C3096 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 5_bit_dac_0[1].switch_n_3v3_0.D2 0.0719f
C3097 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.805f
C3098 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 0.0904f
C3099 a_1556_7774# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.296f
C3100 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 2.78e-19
C3101 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.836f
C3102 5_bit_dac_0[0].4_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.00583f
C3103 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH a_1556_1634# 1.97e-19
C3104 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.00491f
C3105 5_bit_dac_0[1].4_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.0057f
C3106 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].D0 0.0179f
C3107 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.DX_ 0.125f
C3108 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.205f
C3109 5_bit_dac_0[1].4_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 0.044f
C3110 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].D0 0.544f
C3111 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.00491f
C3112 D4 5_bit_dac_0[1].4_bit_dac_0[0].VOUT 1.26e-20
C3113 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.205f
C3114 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 4.25e-19
C3115 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.349f
C3116 VCC a_1556_17598# 0.713f
C3117 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L a_1556_12686# 1.29e-19
C3118 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.714f
C3119 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.0261f
C3120 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.00692f
C3121 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.805f
C3122 D5_BUF 5_bit_dac_0[0].switch_n_3v3_0.DX_ 1.8e-19
C3123 switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 0.177f
C3124 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 0.0904f
C3125 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 2.49e-22
C3126 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00394f
C3127 5_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2.38e-19
C3128 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.00491f
C3129 a_1556_6546# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0892f
C3130 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 0.797f
C3131 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.622f
C3132 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VREFL 0.0988f
C3133 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH switch_n_3v3_0.D6 3.83e-20
C3134 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ D5_BUF 6.33e-20
C3135 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0018f
C3136 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00123f
C3137 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.045f
C3138 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 0.00105f
C3139 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 0.219f
C3140 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.404f
C3141 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 3.62e-20
C3142 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 9.82e-21
C3143 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.622f
C3144 5_bit_dac_0[0].4_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].VOUT 0.34f
C3145 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.312f
C3146 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00143f
C3147 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0018f
C3148 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 1.46e-19
C3149 VCC 5_bit_dac_0[0].switch_n_3v3_0.D2 0.779f
C3150 5_bit_dac_0[1].4_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 0.546f
C3151 a_1556_1634# D0_BUF 0.00365f
C3152 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ switch_n_3v3_0.D4 6.07e-19
C3153 5_bit_dac_0[0].VOUT 5_bit_dac_0[0].switch_n_3v3_0.D2 3.6e-20
C3154 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0668f
C3155 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L a_1556_10230# 1.29e-19
C3156 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.00183f
C3157 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.0261f
C3158 5_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.132f
C3159 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H a_1556_4090# 4.83e-19
C3160 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 0.291f
C3161 a_1556_5318# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 4.09e-19
C3162 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 8.21e-19
C3163 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 2.34e-21
C3164 5_bit_dac_0[1].4_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.404f
C3165 5_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.14f
C3166 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 2.34e-21
C3167 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0927f
C3168 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 1.9e-19
C3169 5_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 0.0026f
C3170 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00473f
C3171 VREFL a_1556_17598# 1.97e-19
C3172 5_bit_dac_0[1].4_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3.53e-19
C3173 switch_n_3v3_0.D2 5_bit_dac_0[0].D1 0.0189f
C3174 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.00491f
C3175 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 6.14e-19
C3176 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.037f
C3177 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 0.797f
C3178 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.504f
C3179 a_1556_12686# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 6.04e-19
C3180 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 switch_n_3v3_0.D7 1.57e-20
C3181 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 1.85e-19
C3182 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 0.14f
C3183 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 0.0179f
C3184 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 9.68e-20
C3185 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].VOUT 0.546f
C3186 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH D0 0.00555f
C3187 5_bit_dac_0[1].VOUT switch_n_3v3_0.D3 0.00191f
C3188 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.39f
C3189 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 0.0189f
C3190 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].D1 0.0757f
C3191 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5.59e-19
C3192 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].D0 0.00349f
C3193 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.303f
C3194 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ D4 2.51e-19
C3195 VCC a_1556_18826# 0.713f
C3196 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00473f
C3197 VCC 5_bit_dac_0[1].4_bit_dac_0[1].VOUT 0.775f
C3198 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.836f
C3199 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH a_1556_6546# 0.175f
C3200 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 1.85e-19
C3201 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 3.8e-20
C3202 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.613f
C3203 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H a_1556_11458# 0.397f
C3204 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL switch_n_3v3_0.D7 0.00143f
C3205 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 9.68e-20
C3206 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.249f
C3207 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.404f
C3208 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ 5_bit_dac_0[1].switch_n_3v3_0.DX_ 0.0104f
C3209 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 0.00375f
C3210 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ switch_n_3v3_0.D7 0.0268f
C3211 switch_n_3v3_0.D3 D5 0.0318f
C3212 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].VOUT switch_n_3v3_0.D4 1.79e-20
C3213 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ D5 2.07e-19
C3214 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 3.7e-20
C3215 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.00819f
C3216 a_1556_4090# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 4.09e-19
C3217 D3_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0269f
C3218 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H a_1556_2862# 4.83e-19
C3219 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 0.0104f
C3220 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 0.044f
C3221 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0172f
C3222 5_bit_dac_0[1].4_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.176f
C3223 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 1.06e-19
C3224 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0801f
C3225 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 1.81e-20
C3226 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 4.25e-19
C3227 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT switch_n_3v3_0.D6 0.027f
C3228 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.DX_ switch_n_3v3_0.D7 0.0268f
C3229 D2_BUF switch_n_3v3_0.D7 0.0399f
C3230 5_bit_dac_0[0].4_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.213f
C3231 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 2.05e-20
C3232 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].VOUT 0.017f
C3233 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL D5 0.00306f
C3234 switch_n_3v3_0.D4 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 2.51e-19
C3235 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 1.85e-19
C3236 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0172f
C3237 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH a_1556_5318# 0.337f
C3238 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5.89e-20
C3239 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].switch_n_3v3_0.D2 0.0155f
C3240 VOUT switch_n_3v3_0.D6 2.3e-20
C3241 a_1556_18826# VREFL 0.337f
C3242 a_1556_17598# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.296f
C3243 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.189f
C3244 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.315f
C3245 5_bit_dac_0[0].4_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 3.38e-20
C3246 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.00379f
C3247 5_bit_dac_0[1].4_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.13f
C3248 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.0104f
C3249 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.189f
C3250 5_bit_dac_0[1].4_bit_dac_0[1].VREFH a_1556_13914# 0.337f
C3251 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 0.044f
C3252 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.0018f
C3253 switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.129f
C3254 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH a_1556_9002# 1.97e-19
C3255 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 4.25e-19
C3256 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].VOUT 0.00119f
C3257 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.349f
C3258 switch_n_3v3_0.D4 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.00127f
C3259 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ switch_n_3v3_0.D6 2.54e-19
C3260 a_1556_2862# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0892f
C3261 VCC 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 1.18f
C3262 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].VOUT 0.00174f
C3263 5_bit_dac_0[1].VREFH a_1556_7774# 1.97e-19
C3264 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.635f
C3265 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.603f
C3266 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.805f
C3267 VCC D1_BUF 0.317f
C3268 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH a_1556_406# 0.337f
C3269 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0801f
C3270 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00473f
C3271 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 D3_BUF 0.631f
C3272 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.0211f
C3273 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.189f
C3274 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 D5 0.0616f
C3275 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT D5 0.0259f
C3276 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 0.219f
C3277 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.836f
C3278 switch_n_3v3_0.D4 D4_BUF 0.0541f
C3279 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VREFH a_1556_406# 1.97e-19
C3280 5_bit_dac_0[0].4_bit_dac_0[1].VOUT switch_n_3v3_0.D6 4.1e-20
C3281 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00163f
C3282 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VREFH a_1556_10230# 1.97e-19
C3283 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.302f
C3284 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 0.0858f
C3285 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.68e-19
C3286 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH a_1556_16370# 1.97e-19
C3287 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 2.69e-19
C3288 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH a_1556_4090# 2.68e-20
C3289 5_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0145f
C3290 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 4.97e-19
C3291 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.00491f
C3292 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5.59e-19
C3293 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 9.82e-21
C3294 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.DX_ 1.8e-19
C3295 switch_n_3v3_0.D4 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.00127f
C3296 switch_n_3v3_0.D4 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.233f
C3297 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.00832f
C3298 D3 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.00213f
C3299 switch_n_3v3_0.D4 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 2.52e-20
C3300 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00143f
C3301 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 5_bit_dac_0[1].switch_n_3v3_0.DX_ 1.05e-19
C3302 a_1556_1634# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 6.04e-19
C3303 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 1.34e-20
C3304 5_bit_dac_0[0].D1 switch_n_3v3_0.D7 1.57e-20
C3305 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.051f
C3306 a_1556_5318# 5_bit_dac_0[0].4_bit_dac_0[0].D0 0.325f
C3307 D0 a_1556_18826# 0.0975f
C3308 a_1556_15142# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.0331f
C3309 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 1.06e-19
C3310 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 0.219f
C3311 5_bit_dac_0[1].4_bit_dac_0[0].D1 D4 4.72e-19
C3312 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 0.0858f
C3313 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 4.15e-19
C3314 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.DX_ 1.34e-20
C3315 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 2.66e-20
C3316 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 4.25e-19
C3317 5_bit_dac_0[0].4_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 0.044f
C3318 a_1556_17598# a_1556_16370# 0.00981f
C3319 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.189f
C3320 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.29f
C3321 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT D5 0.0234f
C3322 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL switch_n_3v3_0.D6 0.00202f
C3323 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 8.92e-19
C3324 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.312f
C3325 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.115f
C3326 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.482f
C3327 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 1.48e-19
C3328 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0927f
C3329 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ D1_BUF 0.219f
C3330 a_1556_406# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.296f
C3331 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.0129f
C3332 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[1].VOUT 0.0743f
C3333 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.315f
C3334 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 1.9e-19
C3335 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00872f
C3336 a_1556_18826# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 2.93e-19
C3337 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 0.0988f
C3338 VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 1.05e-19
C3339 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.511f
C3340 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.00163f
C3341 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH a_1556_11458# 9.57e-20
C3342 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.00832f
C3343 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VOUT switch_n_3v3_0.D6 4.32e-20
C3344 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 6.11e-19
C3345 5_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.111f
C3346 a_1556_16370# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 4.09e-19
C3347 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H a_1556_15142# 4.83e-19
C3348 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 2.34e-21
C3349 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5.84e-19
C3350 switch_n_3v3_0.D4 5_bit_dac_0[0].switch_n_3v3_0.DX_ 0.0904f
C3351 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.13f
C3352 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 0.00379f
C3353 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.00349f
C3354 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.463f
C3355 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].VOUT 5.16e-19
C3356 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.00491f
C3357 switch_n_3v3_0.D4 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.00127f
C3358 VCC a_1556_9002# 0.713f
C3359 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.00105f
C3360 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ switch_n_3v3_0.D7 1.45e-19
C3361 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.205f
C3362 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 0.0988f
C3363 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 switch_n_3v3_0.D6 1.79e-20
C3364 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.579f
C3365 switch_n_3v3_0.D4 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 3.75e-19
C3366 5_bit_dac_0[1].switch_n_3v3_0.D2 D4 0.0361f
C3367 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].VOUT 0.252f
C3368 5_bit_dac_0[1].switch_n_3v3_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.0143f
C3369 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].VOUT 5.16e-19
C3370 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 0.00262f
C3371 switch_n_3v3_0.DX_ VOUT 0.236f
C3372 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 7.75e-19
C3373 VCC 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.77f
C3374 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.0261f
C3375 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT switch_n_3v3_0.D6 0.027f
C3376 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.0102f
C3377 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.472f
C3378 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 4.25e-19
C3379 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL switch_n_3v3_0.D7 0.00143f
C3380 a_1556_16370# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 6.04e-19
C3381 5_bit_dac_0[0].4_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 0.0579f
C3382 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 0.0923f
C3383 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[0].D1 4.15e-19
C3384 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 3.38e-20
C3385 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH a_1556_16370# 2.68e-20
C3386 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.00105f
C3387 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.404f
C3388 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 2.38e-19
C3389 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ switch_n_3v3_0.DX_ 0.0104f
C3390 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.39f
C3391 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5.89e-20
C3392 a_1556_12686# 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 0.00365f
C3393 VCC VOUT 0.394f
C3394 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 a_1556_11458# 0.0981f
C3395 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.00368f
C3396 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.322f
C3397 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 0.0904f
C3398 VOUT 5_bit_dac_0[0].VOUT 0.31f
C3399 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL switch_n_3v3_0.D7 0.00143f
C3400 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.322f
C3401 5_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT 0.00117f
C3402 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].D0 4.97e-19
C3403 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VOUT 0.552f
C3404 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 7.75e-19
C3405 a_1556_17598# 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 1.21e-20
C3406 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 2.51e-20
C3407 VCC 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ 0.712f
C3408 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.00476f
C3409 5_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VOUT 1.75e-20
C3410 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 0.0179f
C3411 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00394f
C3412 5_bit_dac_0[1].switch_n_3v3_0.D3 switch_n_3v3_0.D3 0.0618f
C3413 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.037f
C3414 a_1556_4090# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 0.0892f
C3415 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 0.00594f
C3416 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 0.544f
C3417 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5.59e-19
C3418 5_bit_dac_0[1].VOUT switch_n_3v3_0.D6 3.73e-20
C3419 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H 3.62e-20
C3420 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 1.06f
C3421 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 4.25e-19
C3422 5_bit_dac_0[1].4_bit_dac_0[1].VREFH 5_bit_dac_0[1].4_bit_dac_0[0].D1 1.7e-19
C3423 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.404f
C3424 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 3.36e-19
C3425 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 1.68e-19
C3426 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL D4 0.00517f
C3427 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.DX_ switch_n_3v3_0.D3 0.219f
C3428 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 9.68e-20
C3429 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.DX_ 1.79e-20
C3430 VCC 5_bit_dac_0[0].4_bit_dac_0[1].VOUT 0.735f
C3431 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.129f
C3432 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.236f
C3433 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 2.66e-20
C3434 5_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].VOUT 1.52f
C3435 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 switch_n_3v3_0.D7 0.0916f
C3436 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL switch_n_3v3_0.D7 0.00143f
C3437 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH switch_n_3v3_0.D7 4.71e-19
C3438 switch_n_3v3_0.D4 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 2.09e-21
C3439 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 2.05e-20
C3440 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 0.0057f
C3441 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.128f
C3442 5_bit_dac_0[0].switch_n_3v3_0.D3 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.0295f
C3443 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H 0.037f
C3444 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 1.46e-19
C3445 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.0172f
C3446 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 0.219f
C3447 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 1.06e-19
C3448 D2_BUF 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 1.98e-19
C3449 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].D1 0.00375f
C3450 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 7.75e-19
C3451 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 5_bit_dac_0[0].D0 0.0179f
C3452 switch_n_3v3_0.D4 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 2.45e-20
C3453 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 0.24f
C3454 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L 9.68e-20
C3455 D3 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].VOUT 1.26e-20
C3456 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH 5_bit_dac_0[0].D0 0.544f
C3457 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.322f
C3458 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5.59e-19
C3459 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 0.044f
C3460 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.0018f
C3461 switch_n_3v3_0.D2 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.14f
C3462 D5 switch_n_3v3_0.D6 4.78f
C3463 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.00473f
C3464 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 1.46e-19
C3465 a_1556_9002# 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH 0.0331f
C3466 5_bit_dac_0[1].4_bit_dac_0[0].VOUT switch_n_3v3_0.D3 0.0719f
C3467 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 5_bit_dac_0[1].switch_n_3v3_0.D3 0.631f
C3468 5_bit_dac_0[1].switch_n_3v3_0.D3 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 0.0265f
C3469 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH 0.00577f
C3470 VCC 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL 0.312f
C3471 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.189f
C3472 5_bit_dac_0[0].4_bit_dac_0[1].VREFH 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H 3.7e-20
C3473 D5_BUF 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 0.067f
C3474 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.111f
C3475 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 6.11e-19
C3476 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT 5_bit_dac_0[1].4_bit_dac_0[0].D1 1.81e-20
C3477 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH 0.347f
C3478 a_1556_2862# 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 0.325f
C3479 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VOUT switch_n_3v3_0.DX_ 1.05e-19
C3480 D4_BUF 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.0135f
C3481 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL 0.0172f
C3482 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT 0.0134f
C3483 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ switch_n_3v3_0.D6 2.54e-19
C3484 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VOUT 1.85e-20
C3485 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H a_1556_1634# 0.397f
C3486 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ 0.00819f
C3487 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH 3.82e-19
R0 D0_BUF.n15 D0_BUF.n0 400.238
R1 D0_BUF.n3 D0_BUF.n2 292.5
R2 D0_BUF.n17 D0_BUF.n16 153.333
R3 D0_BUF D0_BUF.n17 105.785
R4 D0_BUF.n0 D0_BUF.t2 83.8685
R5 D0_BUF.n16 D0_BUF.t5 80.9765
R6 D0_BUF.n16 D0_BUF.t3 57.8405
R7 D0_BUF.n0 D0_BUF.t4 54.9485
R8 D0_BUF.n5 D0_BUF.t1 47.274
R9 D0_BUF.n2 D0_BUF.t0 27.6955
R10 D0_BUF.n17 D0_BUF.n15 23.9595
R11 D0_BUF.n11 D0_BUF.n3 13.177
R12 D0_BUF.n8 D0_BUF.n3 13.177
R13 D0_BUF.n11 D0_BUF.n10 9.3005
R14 D0_BUF.n9 D0_BUF.n8 9.3005
R15 D0_BUF.n6 D0_BUF.n5 9.3005
R16 D0_BUF.n7 D0_BUF.n4 9.3005
R17 D0_BUF.n12 D0_BUF.n1 9.3005
R18 D0_BUF.n14 D0_BUF.n13 9.3005
R19 D0_BUF.n13 D0_BUF.n2 9.02061
R20 D0_BUF.n6 D0_BUF.n2 9.0206
R21 D0_BUF.n13 D0_BUF.n12 6.02403
R22 D0_BUF.n7 D0_BUF.n6 6.02403
R23 D0_BUF.n15 D0_BUF 5.08342
R24 D0_BUF D0_BUF.n14 2.37139
R25 D0_BUF.n12 D0_BUF.n11 0.376971
R26 D0_BUF.n8 D0_BUF.n7 0.376971
R27 D0_BUF.n10 D0_BUF.n9 0.190717
R28 D0_BUF.n14 D0_BUF.n1 0.0439783
R29 D0_BUF.n5 D0_BUF.n4 0.0439783
R30 D0_BUF.n10 D0_BUF.n1 0.00321739
R31 D0_BUF.n9 D0_BUF.n4 0.00321739
R32 VCC.n426 VCC.t282 4282.54
R33 VCC.n978 VCC.t136 4282.54
R34 VCC.n1536 VCC.t1 4282.54
R35 VCC.n2087 VCC.t47 4282.54
R36 VCC.n2645 VCC.t200 4282.54
R37 VCC.n3196 VCC.t273 4282.54
R38 VCC.n3754 VCC.t101 4282.54
R39 VCC.n4305 VCC.t267 4282.54
R40 VCC.n4863 VCC.t118 4282.54
R41 VCC.n5414 VCC.t10 4282.54
R42 VCC.n5971 VCC.t239 4282.54
R43 VCC.n6521 VCC.t87 4282.54
R44 VCC.n7078 VCC.t310 4282.54
R45 VCC.n7628 VCC.t37 4282.54
R46 VCC.n8185 VCC.t297 4282.54
R47 VCC.n8548 VCC.t129 4282.54
R48 VCC.t254 VCC.t283 1149.1
R49 VCC.t31 VCC.t133 1149.1
R50 VCC.t26 VCC.t0 1149.1
R51 VCC.t23 VCC.t44 1149.1
R52 VCC.t189 VCC.t197 1149.1
R53 VCC.t97 VCC.t272 1149.1
R54 VCC.t271 VCC.t98 1149.1
R55 VCC.t302 VCC.t266 1149.1
R56 VCC.t111 VCC.t115 1149.1
R57 VCC.t225 VCC.t7 1149.1
R58 VCC.t247 VCC.t240 1149.1
R59 VCC.t167 VCC.t84 1149.1
R60 VCC.t110 VCC.t307 1149.1
R61 VCC.t71 VCC.t38 1149.1
R62 VCC.t220 VCC.t296 1149.1
R63 VCC.t67 VCC.t128 1149.1
R64 VCC.t282 VCC.t254 978.443
R65 VCC.t136 VCC.t31 978.443
R66 VCC.t1 VCC.t26 978.443
R67 VCC.t47 VCC.t23 978.443
R68 VCC.t200 VCC.t189 978.443
R69 VCC.t273 VCC.t97 978.443
R70 VCC.t101 VCC.t271 978.443
R71 VCC.t267 VCC.t302 978.443
R72 VCC.t118 VCC.t111 978.443
R73 VCC.t10 VCC.t225 978.443
R74 VCC.t239 VCC.t247 978.443
R75 VCC.t87 VCC.t167 978.443
R76 VCC.t310 VCC.t110 978.443
R77 VCC.t37 VCC.t71 978.443
R78 VCC.t297 VCC.t220 978.443
R79 VCC.t129 VCC.t67 978.443
R80 VCC.t283 VCC.t251 972.755
R81 VCC.t133 VCC.t28 972.755
R82 VCC.t0 VCC.t27 972.755
R83 VCC.t44 VCC.t20 972.755
R84 VCC.t197 VCC.t190 972.755
R85 VCC.t272 VCC.t94 972.755
R86 VCC.t98 VCC.t268 972.755
R87 VCC.t266 VCC.t303 972.755
R88 VCC.t115 VCC.t112 972.755
R89 VCC.t7 VCC.t222 972.755
R90 VCC.t240 VCC.t244 972.755
R91 VCC.t84 VCC.t168 972.755
R92 VCC.t307 VCC.t107 972.755
R93 VCC.t38 VCC.t72 972.755
R94 VCC.t296 VCC.t217 972.755
R95 VCC.t128 VCC.t68 972.755
R96 VCC.t251 VCC.n425 723.087
R97 VCC.t28 VCC.n977 723.087
R98 VCC.t27 VCC.n1535 723.087
R99 VCC.t20 VCC.n2086 723.087
R100 VCC.t190 VCC.n2644 723.087
R101 VCC.t94 VCC.n3195 723.087
R102 VCC.t268 VCC.n3753 723.087
R103 VCC.t303 VCC.n4304 723.087
R104 VCC.t112 VCC.n4862 723.087
R105 VCC.t222 VCC.n5413 723.087
R106 VCC.t244 VCC.n5970 723.087
R107 VCC.t168 VCC.n6520 723.087
R108 VCC.t107 VCC.n7077 723.087
R109 VCC.t72 VCC.n7627 723.087
R110 VCC.t217 VCC.n8184 723.087
R111 VCC.t68 VCC.n8547 723.087
R112 VCC.t151 VCC.t261 571.485
R113 VCC.t211 VCC.t250 571.485
R114 VCC.t146 VCC.t304 571.485
R115 VCC.t257 VCC.t104 571.485
R116 VCC.t17 VCC.t137 571.485
R117 VCC.t34 VCC.t6 571.485
R118 VCC.t90 VCC.t210 571.485
R119 VCC.t145 VCC.t49 571.485
R120 VCC.t229 VCC.t194 571.485
R121 VCC.t313 VCC.t228 571.485
R122 VCC.t127 VCC.t184 571.485
R123 VCC.t183 VCC.t291 571.485
R124 VCC.t93 VCC.t180 571.485
R125 VCC.t177 VCC.t286 571.485
R126 VCC.t204 VCC.t75 571.485
R127 VCC.t122 VCC.t201 571.485
R128 VCC.t163 VCC.t158 571.485
R129 VCC.t258 VCC.t58 571.485
R130 VCC.t171 VCC.t142 571.485
R131 VCC.t241 VCC.t232 571.485
R132 VCC.t164 VCC.t193 571.485
R133 VCC.t81 VCC.t52 571.485
R134 VCC.t221 VCC.t61 571.485
R135 VCC.t132 VCC.t14 571.485
R136 VCC.t62 VCC.t155 571.485
R137 VCC.t205 VCC.t43 571.485
R138 VCC.t48 VCC.t11 571.485
R139 VCC.t119 VCC.t281 571.485
R140 VCC.t278 VCC.t214 571.485
R141 VCC.t174 VCC.t80 571.485
R142 VCC.t55 VCC.t154 571.485
R143 VCC.n122 VCC.t211 544.823
R144 VCC.n674 VCC.t257 544.823
R145 VCC.n1231 VCC.t17 544.823
R146 VCC.n1783 VCC.t145 544.823
R147 VCC.n2340 VCC.t229 544.823
R148 VCC.n2892 VCC.t183 544.823
R149 VCC.n3449 VCC.t93 544.823
R150 VCC.n4001 VCC.t122 544.823
R151 VCC.n4558 VCC.t163 544.823
R152 VCC.n5110 VCC.t241 544.823
R153 VCC.n5666 VCC.t164 544.823
R154 VCC.n6217 VCC.t132 544.823
R155 VCC.n6773 VCC.t62 544.823
R156 VCC.n7324 VCC.t119 544.823
R157 VCC.n7880 VCC.t278 544.823
R158 VCC.n8431 VCC.t55 544.823
R159 VCC.n209 VCC.t151 542.996
R160 VCC.n761 VCC.t146 542.996
R161 VCC.n1319 VCC.t34 542.996
R162 VCC.n1870 VCC.t90 542.996
R163 VCC.n2428 VCC.t313 542.996
R164 VCC.n2979 VCC.t127 542.996
R165 VCC.n3537 VCC.t177 542.996
R166 VCC.n4088 VCC.t204 542.996
R167 VCC.n4646 VCC.t258 542.996
R168 VCC.n5197 VCC.t171 542.996
R169 VCC.n5754 VCC.t81 542.996
R170 VCC.n6304 VCC.t221 542.996
R171 VCC.n6861 VCC.t205 542.996
R172 VCC.n7411 VCC.t48 542.996
R173 VCC.n7968 VCC.t174 542.996
R174 VCC.n209 VCC.n194 187.349
R175 VCC.n123 VCC.n122 187.349
R176 VCC.n426 VCC.n79 187.349
R177 VCC.n761 VCC.n746 187.349
R178 VCC.n675 VCC.n674 187.349
R179 VCC.n978 VCC.n631 187.349
R180 VCC.n1232 VCC.n1231 187.349
R181 VCC.n1536 VCC.n1188 187.349
R182 VCC.n1319 VCC.n1304 187.349
R183 VCC.n1870 VCC.n1855 187.349
R184 VCC.n1784 VCC.n1783 187.349
R185 VCC.n2087 VCC.n1740 187.349
R186 VCC.n2341 VCC.n2340 187.349
R187 VCC.n2645 VCC.n2297 187.349
R188 VCC.n2428 VCC.n2413 187.349
R189 VCC.n2979 VCC.n2964 187.349
R190 VCC.n2893 VCC.n2892 187.349
R191 VCC.n3196 VCC.n2849 187.349
R192 VCC.n3450 VCC.n3449 187.349
R193 VCC.n3754 VCC.n3406 187.349
R194 VCC.n3537 VCC.n3522 187.349
R195 VCC.n4088 VCC.n4073 187.349
R196 VCC.n4002 VCC.n4001 187.349
R197 VCC.n4305 VCC.n3958 187.349
R198 VCC.n4559 VCC.n4558 187.349
R199 VCC.n4863 VCC.n4515 187.349
R200 VCC.n4646 VCC.n4631 187.349
R201 VCC.n5197 VCC.n5182 187.349
R202 VCC.n5111 VCC.n5110 187.349
R203 VCC.n5414 VCC.n5067 187.349
R204 VCC.n5667 VCC.n5666 187.349
R205 VCC.n5971 VCC.n5623 187.349
R206 VCC.n5754 VCC.n5739 187.349
R207 VCC.n6304 VCC.n6289 187.349
R208 VCC.n6218 VCC.n6217 187.349
R209 VCC.n6521 VCC.n6174 187.349
R210 VCC.n6774 VCC.n6773 187.349
R211 VCC.n7078 VCC.n6730 187.349
R212 VCC.n6861 VCC.n6846 187.349
R213 VCC.n7411 VCC.n7396 187.349
R214 VCC.n7325 VCC.n7324 187.349
R215 VCC.n7628 VCC.n7281 187.349
R216 VCC.n7881 VCC.n7880 187.349
R217 VCC.n8185 VCC.n7837 187.349
R218 VCC.n7968 VCC.n7953 187.349
R219 VCC.n8432 VCC.n8431 187.349
R220 VCC.n8548 VCC.n8388 187.349
R221 VCC.n231 VCC.n230 185
R222 VCC.n230 VCC.n229 185
R223 VCC.n270 VCC.n269 185
R224 VCC.n269 VCC.n268 185
R225 VCC.n286 VCC.n140 185
R226 VCC.n290 VCC.n140 185
R227 VCC.n292 VCC.n141 185
R228 VCC.n292 VCC.n291 185
R229 VCC.n271 VCC.n143 185
R230 VCC.n143 VCC.n142 185
R231 VCC.n210 VCC.n208 185
R232 VCC.n183 VCC.n182 185
R233 VCC.n182 VCC.n181 185
R234 VCC.n225 VCC.n224 185
R235 VCC.n226 VCC.n225 185
R236 VCC.n180 VCC.n178 185
R237 VCC.n228 VCC.n180 185
R238 VCC.n359 VCC.n358 185
R239 VCC.n360 VCC.n359 185
R240 VCC.n92 VCC.n91 185
R241 VCC.n395 VCC.n92 185
R242 VCC.n416 VCC.n415 185
R243 VCC.n417 VCC.n416 185
R244 VCC.n414 VCC.n80 185
R245 VCC.n418 VCC.n80 185
R246 VCC.n398 VCC.n397 185
R247 VCC.n397 VCC.n396 185
R248 VCC.n427 VCC.n81 185
R249 VCC.n121 VCC.n120 185
R250 VCC.n119 VCC.n118 185
R251 VCC.n336 VCC.n119 185
R252 VCC.n339 VCC.n338 185
R253 VCC.n338 VCC.n337 185
R254 VCC.n107 VCC.n106 185
R255 VCC.n361 VCC.n107 185
R256 VCC.n546 VCC.n545 185
R257 VCC.n547 VCC.n546 185
R258 VCC.n421 VCC.n56 185
R259 VCC.n419 VCC.n56 185
R260 VCC.n493 VCC.n39 185
R261 VCC.n494 VCC.n493 185
R262 VCC.n21 VCC.n20 185
R263 VCC.n526 VCC.n21 185
R264 VCC.n529 VCC.n528 185
R265 VCC.n528 VCC.n527 185
R266 VCC.n24 VCC.n23 185
R267 VCC.n23 VCC.n22 185
R268 VCC.n498 VCC.n497 185
R269 VCC.n497 VCC.n496 185
R270 VCC.n492 VCC.n491 185
R271 VCC.n492 VCC.n41 185
R272 VCC.n475 VCC.n474 185
R273 VCC.n474 VCC.n473 185
R274 VCC.n55 VCC.n54 185
R275 VCC.n471 VCC.n55 185
R276 VCC.n423 VCC.n422 185
R277 VCC.n423 VCC.n420 185
R278 VCC.n4 VCC.n3 185
R279 VCC.n783 VCC.n782 185
R280 VCC.n782 VCC.n781 185
R281 VCC.n822 VCC.n821 185
R282 VCC.n821 VCC.n820 185
R283 VCC.n838 VCC.n692 185
R284 VCC.n842 VCC.n692 185
R285 VCC.n844 VCC.n693 185
R286 VCC.n844 VCC.n843 185
R287 VCC.n823 VCC.n695 185
R288 VCC.n695 VCC.n694 185
R289 VCC.n762 VCC.n760 185
R290 VCC.n735 VCC.n734 185
R291 VCC.n734 VCC.n733 185
R292 VCC.n777 VCC.n776 185
R293 VCC.n778 VCC.n777 185
R294 VCC.n732 VCC.n730 185
R295 VCC.n780 VCC.n732 185
R296 VCC.n911 VCC.n910 185
R297 VCC.n912 VCC.n911 185
R298 VCC.n644 VCC.n643 185
R299 VCC.n947 VCC.n644 185
R300 VCC.n968 VCC.n967 185
R301 VCC.n969 VCC.n968 185
R302 VCC.n966 VCC.n632 185
R303 VCC.n970 VCC.n632 185
R304 VCC.n950 VCC.n949 185
R305 VCC.n949 VCC.n948 185
R306 VCC.n979 VCC.n633 185
R307 VCC.n673 VCC.n672 185
R308 VCC.n671 VCC.n670 185
R309 VCC.n888 VCC.n671 185
R310 VCC.n891 VCC.n890 185
R311 VCC.n890 VCC.n889 185
R312 VCC.n659 VCC.n658 185
R313 VCC.n913 VCC.n659 185
R314 VCC.n973 VCC.n608 185
R315 VCC.n971 VCC.n608 185
R316 VCC.n607 VCC.n606 185
R317 VCC.n1023 VCC.n607 185
R318 VCC.n1044 VCC.n1043 185
R319 VCC.n1044 VCC.n593 185
R320 VCC.n576 VCC.n575 185
R321 VCC.n575 VCC.n574 185
R322 VCC.n1081 VCC.n1080 185
R323 VCC.n1080 VCC.n1079 185
R324 VCC.n1100 VCC.n1099 185
R325 VCC.n1101 VCC.n1100 185
R326 VCC.n1050 VCC.n1049 185
R327 VCC.n1049 VCC.n1048 185
R328 VCC.n1027 VCC.n1026 185
R329 VCC.n1026 VCC.n1025 185
R330 VCC.n1045 VCC.n591 185
R331 VCC.n1046 VCC.n1045 185
R332 VCC.n573 VCC.n572 185
R333 VCC.n1078 VCC.n573 185
R334 VCC.n558 VCC.n557 185
R335 VCC.n975 VCC.n974 185
R336 VCC.n975 VCC.n972 185
R337 VCC.n1531 VCC.n1530 185
R338 VCC.n1530 VCC.n1529 185
R339 VCC.n1579 VCC.n1578 185
R340 VCC.n1580 VCC.n1579 185
R341 VCC.n1162 VCC.n1160 185
R342 VCC.n1584 VCC.n1162 185
R343 VCC.n1142 VCC.n1135 185
R344 VCC.n1620 VCC.n1142 185
R345 VCC.n1650 VCC.n1649 185
R346 VCC.n1651 VCC.n1650 185
R347 VCC.n1654 VCC.n1112 185
R348 VCC.n1654 VCC.n1653 185
R349 VCC.n1116 VCC.n1115 185
R350 VCC.n1115 VCC.n1114 185
R351 VCC.n1618 VCC.n1617 185
R352 VCC.n1619 VCC.n1618 185
R353 VCC.n1582 VCC.n1145 185
R354 VCC.n1583 VCC.n1582 185
R355 VCC.n1161 VCC.n1159 185
R356 VCC.n1581 VCC.n1161 185
R357 VCC.n1656 VCC.n1655 185
R358 VCC.n1533 VCC.n1532 185
R359 VCC.n1533 VCC.n1528 185
R360 VCC.n1448 VCC.n1447 185
R361 VCC.n1447 VCC.n1446 185
R362 VCC.n1216 VCC.n1215 185
R363 VCC.n1470 VCC.n1216 185
R364 VCC.n1201 VCC.n1200 185
R365 VCC.n1504 VCC.n1201 185
R366 VCC.n1525 VCC.n1524 185
R367 VCC.n1526 VCC.n1525 185
R368 VCC.n1523 VCC.n1189 185
R369 VCC.n1527 VCC.n1189 185
R370 VCC.n1468 VCC.n1467 185
R371 VCC.n1469 VCC.n1468 185
R372 VCC.n1228 VCC.n1227 185
R373 VCC.n1445 VCC.n1228 185
R374 VCC.n1507 VCC.n1506 185
R375 VCC.n1506 VCC.n1505 185
R376 VCC.n1537 VCC.n1190 185
R377 VCC.n1230 VCC.n1229 185
R378 VCC.n1335 VCC.n1334 185
R379 VCC.n1336 VCC.n1335 185
R380 VCC.n1290 VCC.n1288 185
R381 VCC.n1338 VCC.n1290 185
R382 VCC.n1380 VCC.n1379 185
R383 VCC.n1379 VCC.n1378 185
R384 VCC.n1396 VCC.n1250 185
R385 VCC.n1400 VCC.n1250 185
R386 VCC.n1402 VCC.n1251 185
R387 VCC.n1402 VCC.n1401 185
R388 VCC.n1341 VCC.n1340 185
R389 VCC.n1340 VCC.n1339 185
R390 VCC.n1293 VCC.n1292 185
R391 VCC.n1292 VCC.n1291 185
R392 VCC.n1381 VCC.n1253 185
R393 VCC.n1253 VCC.n1252 185
R394 VCC.n1320 VCC.n1318 185
R395 VCC.n1892 VCC.n1891 185
R396 VCC.n1891 VCC.n1890 185
R397 VCC.n1931 VCC.n1930 185
R398 VCC.n1930 VCC.n1929 185
R399 VCC.n1947 VCC.n1801 185
R400 VCC.n1951 VCC.n1801 185
R401 VCC.n1953 VCC.n1802 185
R402 VCC.n1953 VCC.n1952 185
R403 VCC.n1932 VCC.n1804 185
R404 VCC.n1804 VCC.n1803 185
R405 VCC.n1871 VCC.n1869 185
R406 VCC.n1844 VCC.n1843 185
R407 VCC.n1843 VCC.n1842 185
R408 VCC.n1886 VCC.n1885 185
R409 VCC.n1887 VCC.n1886 185
R410 VCC.n1841 VCC.n1839 185
R411 VCC.n1889 VCC.n1841 185
R412 VCC.n2020 VCC.n2019 185
R413 VCC.n2021 VCC.n2020 185
R414 VCC.n1753 VCC.n1752 185
R415 VCC.n2056 VCC.n1753 185
R416 VCC.n2077 VCC.n2076 185
R417 VCC.n2078 VCC.n2077 185
R418 VCC.n2075 VCC.n1741 185
R419 VCC.n2079 VCC.n1741 185
R420 VCC.n2059 VCC.n2058 185
R421 VCC.n2058 VCC.n2057 185
R422 VCC.n2088 VCC.n1742 185
R423 VCC.n1782 VCC.n1781 185
R424 VCC.n1780 VCC.n1779 185
R425 VCC.n1997 VCC.n1780 185
R426 VCC.n2000 VCC.n1999 185
R427 VCC.n1999 VCC.n1998 185
R428 VCC.n1768 VCC.n1767 185
R429 VCC.n2022 VCC.n1768 185
R430 VCC.n2082 VCC.n1717 185
R431 VCC.n2080 VCC.n1717 185
R432 VCC.n1716 VCC.n1715 185
R433 VCC.n2132 VCC.n1716 185
R434 VCC.n2153 VCC.n2152 185
R435 VCC.n2153 VCC.n1702 185
R436 VCC.n1685 VCC.n1684 185
R437 VCC.n1684 VCC.n1683 185
R438 VCC.n2190 VCC.n2189 185
R439 VCC.n2189 VCC.n2188 185
R440 VCC.n2209 VCC.n2208 185
R441 VCC.n2210 VCC.n2209 185
R442 VCC.n2159 VCC.n2158 185
R443 VCC.n2158 VCC.n2157 185
R444 VCC.n2136 VCC.n2135 185
R445 VCC.n2135 VCC.n2134 185
R446 VCC.n2154 VCC.n1700 185
R447 VCC.n2155 VCC.n2154 185
R448 VCC.n1682 VCC.n1681 185
R449 VCC.n2187 VCC.n1682 185
R450 VCC.n1667 VCC.n1666 185
R451 VCC.n2084 VCC.n2083 185
R452 VCC.n2084 VCC.n2081 185
R453 VCC.n2640 VCC.n2639 185
R454 VCC.n2639 VCC.n2638 185
R455 VCC.n2688 VCC.n2687 185
R456 VCC.n2689 VCC.n2688 185
R457 VCC.n2271 VCC.n2269 185
R458 VCC.n2693 VCC.n2271 185
R459 VCC.n2251 VCC.n2244 185
R460 VCC.n2729 VCC.n2251 185
R461 VCC.n2759 VCC.n2758 185
R462 VCC.n2760 VCC.n2759 185
R463 VCC.n2763 VCC.n2221 185
R464 VCC.n2763 VCC.n2762 185
R465 VCC.n2225 VCC.n2224 185
R466 VCC.n2224 VCC.n2223 185
R467 VCC.n2727 VCC.n2726 185
R468 VCC.n2728 VCC.n2727 185
R469 VCC.n2691 VCC.n2254 185
R470 VCC.n2692 VCC.n2691 185
R471 VCC.n2270 VCC.n2268 185
R472 VCC.n2690 VCC.n2270 185
R473 VCC.n2765 VCC.n2764 185
R474 VCC.n2642 VCC.n2641 185
R475 VCC.n2642 VCC.n2637 185
R476 VCC.n2557 VCC.n2556 185
R477 VCC.n2556 VCC.n2555 185
R478 VCC.n2325 VCC.n2324 185
R479 VCC.n2579 VCC.n2325 185
R480 VCC.n2310 VCC.n2309 185
R481 VCC.n2613 VCC.n2310 185
R482 VCC.n2634 VCC.n2633 185
R483 VCC.n2635 VCC.n2634 185
R484 VCC.n2632 VCC.n2298 185
R485 VCC.n2636 VCC.n2298 185
R486 VCC.n2577 VCC.n2576 185
R487 VCC.n2578 VCC.n2577 185
R488 VCC.n2337 VCC.n2336 185
R489 VCC.n2554 VCC.n2337 185
R490 VCC.n2616 VCC.n2615 185
R491 VCC.n2615 VCC.n2614 185
R492 VCC.n2646 VCC.n2299 185
R493 VCC.n2339 VCC.n2338 185
R494 VCC.n2444 VCC.n2443 185
R495 VCC.n2445 VCC.n2444 185
R496 VCC.n2399 VCC.n2397 185
R497 VCC.n2447 VCC.n2399 185
R498 VCC.n2489 VCC.n2488 185
R499 VCC.n2488 VCC.n2487 185
R500 VCC.n2505 VCC.n2359 185
R501 VCC.n2509 VCC.n2359 185
R502 VCC.n2511 VCC.n2360 185
R503 VCC.n2511 VCC.n2510 185
R504 VCC.n2450 VCC.n2449 185
R505 VCC.n2449 VCC.n2448 185
R506 VCC.n2402 VCC.n2401 185
R507 VCC.n2401 VCC.n2400 185
R508 VCC.n2490 VCC.n2362 185
R509 VCC.n2362 VCC.n2361 185
R510 VCC.n2429 VCC.n2427 185
R511 VCC.n3001 VCC.n3000 185
R512 VCC.n3000 VCC.n2999 185
R513 VCC.n3040 VCC.n3039 185
R514 VCC.n3039 VCC.n3038 185
R515 VCC.n3056 VCC.n2910 185
R516 VCC.n3060 VCC.n2910 185
R517 VCC.n3062 VCC.n2911 185
R518 VCC.n3062 VCC.n3061 185
R519 VCC.n3041 VCC.n2913 185
R520 VCC.n2913 VCC.n2912 185
R521 VCC.n2980 VCC.n2978 185
R522 VCC.n2953 VCC.n2952 185
R523 VCC.n2952 VCC.n2951 185
R524 VCC.n2995 VCC.n2994 185
R525 VCC.n2996 VCC.n2995 185
R526 VCC.n2950 VCC.n2948 185
R527 VCC.n2998 VCC.n2950 185
R528 VCC.n3129 VCC.n3128 185
R529 VCC.n3130 VCC.n3129 185
R530 VCC.n2862 VCC.n2861 185
R531 VCC.n3165 VCC.n2862 185
R532 VCC.n3186 VCC.n3185 185
R533 VCC.n3187 VCC.n3186 185
R534 VCC.n3184 VCC.n2850 185
R535 VCC.n3188 VCC.n2850 185
R536 VCC.n3168 VCC.n3167 185
R537 VCC.n3167 VCC.n3166 185
R538 VCC.n3197 VCC.n2851 185
R539 VCC.n2891 VCC.n2890 185
R540 VCC.n2889 VCC.n2888 185
R541 VCC.n3106 VCC.n2889 185
R542 VCC.n3109 VCC.n3108 185
R543 VCC.n3108 VCC.n3107 185
R544 VCC.n2877 VCC.n2876 185
R545 VCC.n3131 VCC.n2877 185
R546 VCC.n3191 VCC.n2826 185
R547 VCC.n3189 VCC.n2826 185
R548 VCC.n2825 VCC.n2824 185
R549 VCC.n3241 VCC.n2825 185
R550 VCC.n3262 VCC.n3261 185
R551 VCC.n3262 VCC.n2811 185
R552 VCC.n2794 VCC.n2793 185
R553 VCC.n2793 VCC.n2792 185
R554 VCC.n3299 VCC.n3298 185
R555 VCC.n3298 VCC.n3297 185
R556 VCC.n3318 VCC.n3317 185
R557 VCC.n3319 VCC.n3318 185
R558 VCC.n3268 VCC.n3267 185
R559 VCC.n3267 VCC.n3266 185
R560 VCC.n3245 VCC.n3244 185
R561 VCC.n3244 VCC.n3243 185
R562 VCC.n3263 VCC.n2809 185
R563 VCC.n3264 VCC.n3263 185
R564 VCC.n2791 VCC.n2790 185
R565 VCC.n3296 VCC.n2791 185
R566 VCC.n2776 VCC.n2775 185
R567 VCC.n3193 VCC.n3192 185
R568 VCC.n3193 VCC.n3190 185
R569 VCC.n3749 VCC.n3748 185
R570 VCC.n3748 VCC.n3747 185
R571 VCC.n3797 VCC.n3796 185
R572 VCC.n3798 VCC.n3797 185
R573 VCC.n3380 VCC.n3378 185
R574 VCC.n3802 VCC.n3380 185
R575 VCC.n3360 VCC.n3353 185
R576 VCC.n3838 VCC.n3360 185
R577 VCC.n3868 VCC.n3867 185
R578 VCC.n3869 VCC.n3868 185
R579 VCC.n3872 VCC.n3330 185
R580 VCC.n3872 VCC.n3871 185
R581 VCC.n3334 VCC.n3333 185
R582 VCC.n3333 VCC.n3332 185
R583 VCC.n3836 VCC.n3835 185
R584 VCC.n3837 VCC.n3836 185
R585 VCC.n3800 VCC.n3363 185
R586 VCC.n3801 VCC.n3800 185
R587 VCC.n3379 VCC.n3377 185
R588 VCC.n3799 VCC.n3379 185
R589 VCC.n3874 VCC.n3873 185
R590 VCC.n3751 VCC.n3750 185
R591 VCC.n3751 VCC.n3746 185
R592 VCC.n3666 VCC.n3665 185
R593 VCC.n3665 VCC.n3664 185
R594 VCC.n3434 VCC.n3433 185
R595 VCC.n3688 VCC.n3434 185
R596 VCC.n3419 VCC.n3418 185
R597 VCC.n3722 VCC.n3419 185
R598 VCC.n3743 VCC.n3742 185
R599 VCC.n3744 VCC.n3743 185
R600 VCC.n3741 VCC.n3407 185
R601 VCC.n3745 VCC.n3407 185
R602 VCC.n3686 VCC.n3685 185
R603 VCC.n3687 VCC.n3686 185
R604 VCC.n3446 VCC.n3445 185
R605 VCC.n3663 VCC.n3446 185
R606 VCC.n3725 VCC.n3724 185
R607 VCC.n3724 VCC.n3723 185
R608 VCC.n3755 VCC.n3408 185
R609 VCC.n3448 VCC.n3447 185
R610 VCC.n3553 VCC.n3552 185
R611 VCC.n3554 VCC.n3553 185
R612 VCC.n3508 VCC.n3506 185
R613 VCC.n3556 VCC.n3508 185
R614 VCC.n3598 VCC.n3597 185
R615 VCC.n3597 VCC.n3596 185
R616 VCC.n3614 VCC.n3468 185
R617 VCC.n3618 VCC.n3468 185
R618 VCC.n3620 VCC.n3469 185
R619 VCC.n3620 VCC.n3619 185
R620 VCC.n3559 VCC.n3558 185
R621 VCC.n3558 VCC.n3557 185
R622 VCC.n3511 VCC.n3510 185
R623 VCC.n3510 VCC.n3509 185
R624 VCC.n3599 VCC.n3471 185
R625 VCC.n3471 VCC.n3470 185
R626 VCC.n3538 VCC.n3536 185
R627 VCC.n4110 VCC.n4109 185
R628 VCC.n4109 VCC.n4108 185
R629 VCC.n4149 VCC.n4148 185
R630 VCC.n4148 VCC.n4147 185
R631 VCC.n4165 VCC.n4019 185
R632 VCC.n4169 VCC.n4019 185
R633 VCC.n4171 VCC.n4020 185
R634 VCC.n4171 VCC.n4170 185
R635 VCC.n4150 VCC.n4022 185
R636 VCC.n4022 VCC.n4021 185
R637 VCC.n4089 VCC.n4087 185
R638 VCC.n4062 VCC.n4061 185
R639 VCC.n4061 VCC.n4060 185
R640 VCC.n4104 VCC.n4103 185
R641 VCC.n4105 VCC.n4104 185
R642 VCC.n4059 VCC.n4057 185
R643 VCC.n4107 VCC.n4059 185
R644 VCC.n4238 VCC.n4237 185
R645 VCC.n4239 VCC.n4238 185
R646 VCC.n3971 VCC.n3970 185
R647 VCC.n4274 VCC.n3971 185
R648 VCC.n4295 VCC.n4294 185
R649 VCC.n4296 VCC.n4295 185
R650 VCC.n4293 VCC.n3959 185
R651 VCC.n4297 VCC.n3959 185
R652 VCC.n4277 VCC.n4276 185
R653 VCC.n4276 VCC.n4275 185
R654 VCC.n4306 VCC.n3960 185
R655 VCC.n4000 VCC.n3999 185
R656 VCC.n3998 VCC.n3997 185
R657 VCC.n4215 VCC.n3998 185
R658 VCC.n4218 VCC.n4217 185
R659 VCC.n4217 VCC.n4216 185
R660 VCC.n3986 VCC.n3985 185
R661 VCC.n4240 VCC.n3986 185
R662 VCC.n4300 VCC.n3935 185
R663 VCC.n4298 VCC.n3935 185
R664 VCC.n3934 VCC.n3933 185
R665 VCC.n4350 VCC.n3934 185
R666 VCC.n4371 VCC.n4370 185
R667 VCC.n4371 VCC.n3920 185
R668 VCC.n3903 VCC.n3902 185
R669 VCC.n3902 VCC.n3901 185
R670 VCC.n4408 VCC.n4407 185
R671 VCC.n4407 VCC.n4406 185
R672 VCC.n4427 VCC.n4426 185
R673 VCC.n4428 VCC.n4427 185
R674 VCC.n4377 VCC.n4376 185
R675 VCC.n4376 VCC.n4375 185
R676 VCC.n4354 VCC.n4353 185
R677 VCC.n4353 VCC.n4352 185
R678 VCC.n4372 VCC.n3918 185
R679 VCC.n4373 VCC.n4372 185
R680 VCC.n3900 VCC.n3899 185
R681 VCC.n4405 VCC.n3900 185
R682 VCC.n3885 VCC.n3884 185
R683 VCC.n4302 VCC.n4301 185
R684 VCC.n4302 VCC.n4299 185
R685 VCC.n4858 VCC.n4857 185
R686 VCC.n4857 VCC.n4856 185
R687 VCC.n4906 VCC.n4905 185
R688 VCC.n4907 VCC.n4906 185
R689 VCC.n4489 VCC.n4487 185
R690 VCC.n4911 VCC.n4489 185
R691 VCC.n4469 VCC.n4462 185
R692 VCC.n4947 VCC.n4469 185
R693 VCC.n4977 VCC.n4976 185
R694 VCC.n4978 VCC.n4977 185
R695 VCC.n4981 VCC.n4439 185
R696 VCC.n4981 VCC.n4980 185
R697 VCC.n4443 VCC.n4442 185
R698 VCC.n4442 VCC.n4441 185
R699 VCC.n4945 VCC.n4944 185
R700 VCC.n4946 VCC.n4945 185
R701 VCC.n4909 VCC.n4472 185
R702 VCC.n4910 VCC.n4909 185
R703 VCC.n4488 VCC.n4486 185
R704 VCC.n4908 VCC.n4488 185
R705 VCC.n4983 VCC.n4982 185
R706 VCC.n4860 VCC.n4859 185
R707 VCC.n4860 VCC.n4855 185
R708 VCC.n4775 VCC.n4774 185
R709 VCC.n4774 VCC.n4773 185
R710 VCC.n4543 VCC.n4542 185
R711 VCC.n4797 VCC.n4543 185
R712 VCC.n4528 VCC.n4527 185
R713 VCC.n4831 VCC.n4528 185
R714 VCC.n4852 VCC.n4851 185
R715 VCC.n4853 VCC.n4852 185
R716 VCC.n4850 VCC.n4516 185
R717 VCC.n4854 VCC.n4516 185
R718 VCC.n4795 VCC.n4794 185
R719 VCC.n4796 VCC.n4795 185
R720 VCC.n4555 VCC.n4554 185
R721 VCC.n4772 VCC.n4555 185
R722 VCC.n4834 VCC.n4833 185
R723 VCC.n4833 VCC.n4832 185
R724 VCC.n4864 VCC.n4517 185
R725 VCC.n4557 VCC.n4556 185
R726 VCC.n4662 VCC.n4661 185
R727 VCC.n4663 VCC.n4662 185
R728 VCC.n4617 VCC.n4615 185
R729 VCC.n4665 VCC.n4617 185
R730 VCC.n4707 VCC.n4706 185
R731 VCC.n4706 VCC.n4705 185
R732 VCC.n4723 VCC.n4577 185
R733 VCC.n4727 VCC.n4577 185
R734 VCC.n4729 VCC.n4578 185
R735 VCC.n4729 VCC.n4728 185
R736 VCC.n4668 VCC.n4667 185
R737 VCC.n4667 VCC.n4666 185
R738 VCC.n4620 VCC.n4619 185
R739 VCC.n4619 VCC.n4618 185
R740 VCC.n4708 VCC.n4580 185
R741 VCC.n4580 VCC.n4579 185
R742 VCC.n4647 VCC.n4645 185
R743 VCC.n5219 VCC.n5218 185
R744 VCC.n5218 VCC.n5217 185
R745 VCC.n5258 VCC.n5257 185
R746 VCC.n5257 VCC.n5256 185
R747 VCC.n5274 VCC.n5128 185
R748 VCC.n5278 VCC.n5128 185
R749 VCC.n5280 VCC.n5129 185
R750 VCC.n5280 VCC.n5279 185
R751 VCC.n5259 VCC.n5131 185
R752 VCC.n5131 VCC.n5130 185
R753 VCC.n5198 VCC.n5196 185
R754 VCC.n5171 VCC.n5170 185
R755 VCC.n5170 VCC.n5169 185
R756 VCC.n5213 VCC.n5212 185
R757 VCC.n5214 VCC.n5213 185
R758 VCC.n5168 VCC.n5166 185
R759 VCC.n5216 VCC.n5168 185
R760 VCC.n5347 VCC.n5346 185
R761 VCC.n5348 VCC.n5347 185
R762 VCC.n5080 VCC.n5079 185
R763 VCC.n5383 VCC.n5080 185
R764 VCC.n5404 VCC.n5403 185
R765 VCC.n5405 VCC.n5404 185
R766 VCC.n5402 VCC.n5068 185
R767 VCC.n5406 VCC.n5068 185
R768 VCC.n5386 VCC.n5385 185
R769 VCC.n5385 VCC.n5384 185
R770 VCC.n5415 VCC.n5069 185
R771 VCC.n5109 VCC.n5108 185
R772 VCC.n5107 VCC.n5106 185
R773 VCC.n5324 VCC.n5107 185
R774 VCC.n5327 VCC.n5326 185
R775 VCC.n5326 VCC.n5325 185
R776 VCC.n5095 VCC.n5094 185
R777 VCC.n5349 VCC.n5095 185
R778 VCC.n5409 VCC.n5044 185
R779 VCC.n5407 VCC.n5044 185
R780 VCC.n5043 VCC.n5042 185
R781 VCC.n5459 VCC.n5043 185
R782 VCC.n5480 VCC.n5479 185
R783 VCC.n5480 VCC.n5029 185
R784 VCC.n5012 VCC.n5011 185
R785 VCC.n5011 VCC.n5010 185
R786 VCC.n5517 VCC.n5516 185
R787 VCC.n5516 VCC.n5515 185
R788 VCC.n5536 VCC.n5535 185
R789 VCC.n5537 VCC.n5536 185
R790 VCC.n5486 VCC.n5485 185
R791 VCC.n5485 VCC.n5484 185
R792 VCC.n5463 VCC.n5462 185
R793 VCC.n5462 VCC.n5461 185
R794 VCC.n5481 VCC.n5027 185
R795 VCC.n5482 VCC.n5481 185
R796 VCC.n5009 VCC.n5008 185
R797 VCC.n5514 VCC.n5009 185
R798 VCC.n4994 VCC.n4993 185
R799 VCC.n5411 VCC.n5410 185
R800 VCC.n5411 VCC.n5408 185
R801 VCC.n5966 VCC.n5965 185
R802 VCC.n5965 VCC.n5964 185
R803 VCC.n6014 VCC.n6013 185
R804 VCC.n6015 VCC.n6014 185
R805 VCC.n5597 VCC.n5595 185
R806 VCC.n6019 VCC.n5597 185
R807 VCC.n5577 VCC.n5570 185
R808 VCC.n6055 VCC.n5577 185
R809 VCC.n6085 VCC.n6084 185
R810 VCC.n6086 VCC.n6085 185
R811 VCC.n6089 VCC.n5547 185
R812 VCC.n6089 VCC.n6088 185
R813 VCC.n5551 VCC.n5550 185
R814 VCC.n5550 VCC.n5549 185
R815 VCC.n6053 VCC.n6052 185
R816 VCC.n6054 VCC.n6053 185
R817 VCC.n6017 VCC.n5580 185
R818 VCC.n6018 VCC.n6017 185
R819 VCC.n5596 VCC.n5594 185
R820 VCC.n6016 VCC.n5596 185
R821 VCC.n6091 VCC.n6090 185
R822 VCC.n5968 VCC.n5967 185
R823 VCC.n5968 VCC.n5963 185
R824 VCC.n5883 VCC.n5882 185
R825 VCC.n5882 VCC.n5881 185
R826 VCC.n5651 VCC.n5650 185
R827 VCC.n5905 VCC.n5651 185
R828 VCC.n5636 VCC.n5635 185
R829 VCC.n5939 VCC.n5636 185
R830 VCC.n5960 VCC.n5959 185
R831 VCC.n5961 VCC.n5960 185
R832 VCC.n5958 VCC.n5624 185
R833 VCC.n5962 VCC.n5624 185
R834 VCC.n5903 VCC.n5902 185
R835 VCC.n5904 VCC.n5903 185
R836 VCC.n5663 VCC.n5662 185
R837 VCC.n5880 VCC.n5663 185
R838 VCC.n5942 VCC.n5941 185
R839 VCC.n5941 VCC.n5940 185
R840 VCC.n5972 VCC.n5625 185
R841 VCC.n5665 VCC.n5664 185
R842 VCC.n5770 VCC.n5769 185
R843 VCC.n5771 VCC.n5770 185
R844 VCC.n5725 VCC.n5723 185
R845 VCC.n5773 VCC.n5725 185
R846 VCC.n5815 VCC.n5814 185
R847 VCC.n5814 VCC.n5813 185
R848 VCC.n5831 VCC.n5685 185
R849 VCC.n5835 VCC.n5685 185
R850 VCC.n5837 VCC.n5686 185
R851 VCC.n5837 VCC.n5836 185
R852 VCC.n5776 VCC.n5775 185
R853 VCC.n5775 VCC.n5774 185
R854 VCC.n5728 VCC.n5727 185
R855 VCC.n5727 VCC.n5726 185
R856 VCC.n5816 VCC.n5688 185
R857 VCC.n5688 VCC.n5687 185
R858 VCC.n5755 VCC.n5753 185
R859 VCC.n6326 VCC.n6325 185
R860 VCC.n6325 VCC.n6324 185
R861 VCC.n6365 VCC.n6364 185
R862 VCC.n6364 VCC.n6363 185
R863 VCC.n6381 VCC.n6235 185
R864 VCC.n6385 VCC.n6235 185
R865 VCC.n6387 VCC.n6236 185
R866 VCC.n6387 VCC.n6386 185
R867 VCC.n6366 VCC.n6238 185
R868 VCC.n6238 VCC.n6237 185
R869 VCC.n6305 VCC.n6303 185
R870 VCC.n6278 VCC.n6277 185
R871 VCC.n6277 VCC.n6276 185
R872 VCC.n6320 VCC.n6319 185
R873 VCC.n6321 VCC.n6320 185
R874 VCC.n6275 VCC.n6273 185
R875 VCC.n6323 VCC.n6275 185
R876 VCC.n6454 VCC.n6453 185
R877 VCC.n6455 VCC.n6454 185
R878 VCC.n6187 VCC.n6186 185
R879 VCC.n6490 VCC.n6187 185
R880 VCC.n6511 VCC.n6510 185
R881 VCC.n6512 VCC.n6511 185
R882 VCC.n6509 VCC.n6175 185
R883 VCC.n6513 VCC.n6175 185
R884 VCC.n6493 VCC.n6492 185
R885 VCC.n6492 VCC.n6491 185
R886 VCC.n6522 VCC.n6176 185
R887 VCC.n6216 VCC.n6215 185
R888 VCC.n6214 VCC.n6213 185
R889 VCC.n6431 VCC.n6214 185
R890 VCC.n6434 VCC.n6433 185
R891 VCC.n6433 VCC.n6432 185
R892 VCC.n6202 VCC.n6201 185
R893 VCC.n6456 VCC.n6202 185
R894 VCC.n6516 VCC.n6151 185
R895 VCC.n6514 VCC.n6151 185
R896 VCC.n6150 VCC.n6149 185
R897 VCC.n6566 VCC.n6150 185
R898 VCC.n6587 VCC.n6586 185
R899 VCC.n6587 VCC.n6136 185
R900 VCC.n6119 VCC.n6118 185
R901 VCC.n6118 VCC.n6117 185
R902 VCC.n6624 VCC.n6623 185
R903 VCC.n6623 VCC.n6622 185
R904 VCC.n6643 VCC.n6642 185
R905 VCC.n6644 VCC.n6643 185
R906 VCC.n6593 VCC.n6592 185
R907 VCC.n6592 VCC.n6591 185
R908 VCC.n6570 VCC.n6569 185
R909 VCC.n6569 VCC.n6568 185
R910 VCC.n6588 VCC.n6134 185
R911 VCC.n6589 VCC.n6588 185
R912 VCC.n6116 VCC.n6115 185
R913 VCC.n6621 VCC.n6116 185
R914 VCC.n6101 VCC.n6100 185
R915 VCC.n6518 VCC.n6517 185
R916 VCC.n6518 VCC.n6515 185
R917 VCC.n7073 VCC.n7072 185
R918 VCC.n7072 VCC.n7071 185
R919 VCC.n7121 VCC.n7120 185
R920 VCC.n7122 VCC.n7121 185
R921 VCC.n6704 VCC.n6702 185
R922 VCC.n7126 VCC.n6704 185
R923 VCC.n6684 VCC.n6677 185
R924 VCC.n7162 VCC.n6684 185
R925 VCC.n7192 VCC.n7191 185
R926 VCC.n7193 VCC.n7192 185
R927 VCC.n7196 VCC.n6654 185
R928 VCC.n7196 VCC.n7195 185
R929 VCC.n6658 VCC.n6657 185
R930 VCC.n6657 VCC.n6656 185
R931 VCC.n7160 VCC.n7159 185
R932 VCC.n7161 VCC.n7160 185
R933 VCC.n7124 VCC.n6687 185
R934 VCC.n7125 VCC.n7124 185
R935 VCC.n6703 VCC.n6701 185
R936 VCC.n7123 VCC.n6703 185
R937 VCC.n7198 VCC.n7197 185
R938 VCC.n7075 VCC.n7074 185
R939 VCC.n7075 VCC.n7070 185
R940 VCC.n6990 VCC.n6989 185
R941 VCC.n6989 VCC.n6988 185
R942 VCC.n6758 VCC.n6757 185
R943 VCC.n7012 VCC.n6758 185
R944 VCC.n6743 VCC.n6742 185
R945 VCC.n7046 VCC.n6743 185
R946 VCC.n7067 VCC.n7066 185
R947 VCC.n7068 VCC.n7067 185
R948 VCC.n7065 VCC.n6731 185
R949 VCC.n7069 VCC.n6731 185
R950 VCC.n7010 VCC.n7009 185
R951 VCC.n7011 VCC.n7010 185
R952 VCC.n6770 VCC.n6769 185
R953 VCC.n6987 VCC.n6770 185
R954 VCC.n7049 VCC.n7048 185
R955 VCC.n7048 VCC.n7047 185
R956 VCC.n7079 VCC.n6732 185
R957 VCC.n6772 VCC.n6771 185
R958 VCC.n6877 VCC.n6876 185
R959 VCC.n6878 VCC.n6877 185
R960 VCC.n6832 VCC.n6830 185
R961 VCC.n6880 VCC.n6832 185
R962 VCC.n6922 VCC.n6921 185
R963 VCC.n6921 VCC.n6920 185
R964 VCC.n6938 VCC.n6792 185
R965 VCC.n6942 VCC.n6792 185
R966 VCC.n6944 VCC.n6793 185
R967 VCC.n6944 VCC.n6943 185
R968 VCC.n6883 VCC.n6882 185
R969 VCC.n6882 VCC.n6881 185
R970 VCC.n6835 VCC.n6834 185
R971 VCC.n6834 VCC.n6833 185
R972 VCC.n6923 VCC.n6795 185
R973 VCC.n6795 VCC.n6794 185
R974 VCC.n6862 VCC.n6860 185
R975 VCC.n7433 VCC.n7432 185
R976 VCC.n7432 VCC.n7431 185
R977 VCC.n7472 VCC.n7471 185
R978 VCC.n7471 VCC.n7470 185
R979 VCC.n7488 VCC.n7342 185
R980 VCC.n7492 VCC.n7342 185
R981 VCC.n7494 VCC.n7343 185
R982 VCC.n7494 VCC.n7493 185
R983 VCC.n7473 VCC.n7345 185
R984 VCC.n7345 VCC.n7344 185
R985 VCC.n7412 VCC.n7410 185
R986 VCC.n7385 VCC.n7384 185
R987 VCC.n7384 VCC.n7383 185
R988 VCC.n7427 VCC.n7426 185
R989 VCC.n7428 VCC.n7427 185
R990 VCC.n7382 VCC.n7380 185
R991 VCC.n7430 VCC.n7382 185
R992 VCC.n7561 VCC.n7560 185
R993 VCC.n7562 VCC.n7561 185
R994 VCC.n7294 VCC.n7293 185
R995 VCC.n7597 VCC.n7294 185
R996 VCC.n7618 VCC.n7617 185
R997 VCC.n7619 VCC.n7618 185
R998 VCC.n7616 VCC.n7282 185
R999 VCC.n7620 VCC.n7282 185
R1000 VCC.n7600 VCC.n7599 185
R1001 VCC.n7599 VCC.n7598 185
R1002 VCC.n7629 VCC.n7283 185
R1003 VCC.n7323 VCC.n7322 185
R1004 VCC.n7321 VCC.n7320 185
R1005 VCC.n7538 VCC.n7321 185
R1006 VCC.n7541 VCC.n7540 185
R1007 VCC.n7540 VCC.n7539 185
R1008 VCC.n7309 VCC.n7308 185
R1009 VCC.n7563 VCC.n7309 185
R1010 VCC.n7623 VCC.n7258 185
R1011 VCC.n7621 VCC.n7258 185
R1012 VCC.n7257 VCC.n7256 185
R1013 VCC.n7673 VCC.n7257 185
R1014 VCC.n7694 VCC.n7693 185
R1015 VCC.n7694 VCC.n7243 185
R1016 VCC.n7226 VCC.n7225 185
R1017 VCC.n7225 VCC.n7224 185
R1018 VCC.n7731 VCC.n7730 185
R1019 VCC.n7730 VCC.n7729 185
R1020 VCC.n7750 VCC.n7749 185
R1021 VCC.n7751 VCC.n7750 185
R1022 VCC.n7700 VCC.n7699 185
R1023 VCC.n7699 VCC.n7698 185
R1024 VCC.n7677 VCC.n7676 185
R1025 VCC.n7676 VCC.n7675 185
R1026 VCC.n7695 VCC.n7241 185
R1027 VCC.n7696 VCC.n7695 185
R1028 VCC.n7223 VCC.n7222 185
R1029 VCC.n7728 VCC.n7223 185
R1030 VCC.n7208 VCC.n7207 185
R1031 VCC.n7625 VCC.n7624 185
R1032 VCC.n7625 VCC.n7622 185
R1033 VCC.n8180 VCC.n8179 185
R1034 VCC.n8179 VCC.n8178 185
R1035 VCC.n8228 VCC.n8227 185
R1036 VCC.n8229 VCC.n8228 185
R1037 VCC.n7811 VCC.n7809 185
R1038 VCC.n8233 VCC.n7811 185
R1039 VCC.n7791 VCC.n7784 185
R1040 VCC.n8269 VCC.n7791 185
R1041 VCC.n8299 VCC.n8298 185
R1042 VCC.n8300 VCC.n8299 185
R1043 VCC.n8303 VCC.n7761 185
R1044 VCC.n8303 VCC.n8302 185
R1045 VCC.n7765 VCC.n7764 185
R1046 VCC.n7764 VCC.n7763 185
R1047 VCC.n8267 VCC.n8266 185
R1048 VCC.n8268 VCC.n8267 185
R1049 VCC.n8231 VCC.n7794 185
R1050 VCC.n8232 VCC.n8231 185
R1051 VCC.n7810 VCC.n7808 185
R1052 VCC.n8230 VCC.n7810 185
R1053 VCC.n8305 VCC.n8304 185
R1054 VCC.n8182 VCC.n8181 185
R1055 VCC.n8182 VCC.n8177 185
R1056 VCC.n8097 VCC.n8096 185
R1057 VCC.n8096 VCC.n8095 185
R1058 VCC.n7865 VCC.n7864 185
R1059 VCC.n8119 VCC.n7865 185
R1060 VCC.n7850 VCC.n7849 185
R1061 VCC.n8153 VCC.n7850 185
R1062 VCC.n8174 VCC.n8173 185
R1063 VCC.n8175 VCC.n8174 185
R1064 VCC.n8172 VCC.n7838 185
R1065 VCC.n8176 VCC.n7838 185
R1066 VCC.n8117 VCC.n8116 185
R1067 VCC.n8118 VCC.n8117 185
R1068 VCC.n7877 VCC.n7876 185
R1069 VCC.n8094 VCC.n7877 185
R1070 VCC.n8156 VCC.n8155 185
R1071 VCC.n8155 VCC.n8154 185
R1072 VCC.n8186 VCC.n7839 185
R1073 VCC.n7879 VCC.n7878 185
R1074 VCC.n7984 VCC.n7983 185
R1075 VCC.n7985 VCC.n7984 185
R1076 VCC.n7939 VCC.n7937 185
R1077 VCC.n7987 VCC.n7939 185
R1078 VCC.n8029 VCC.n8028 185
R1079 VCC.n8028 VCC.n8027 185
R1080 VCC.n8045 VCC.n7899 185
R1081 VCC.n8049 VCC.n7899 185
R1082 VCC.n8051 VCC.n7900 185
R1083 VCC.n8051 VCC.n8050 185
R1084 VCC.n7990 VCC.n7989 185
R1085 VCC.n7989 VCC.n7988 185
R1086 VCC.n7942 VCC.n7941 185
R1087 VCC.n7941 VCC.n7940 185
R1088 VCC.n8030 VCC.n7902 185
R1089 VCC.n7902 VCC.n7901 185
R1090 VCC.n7969 VCC.n7967 185
R1091 VCC.n8481 VCC.n8480 185
R1092 VCC.n8482 VCC.n8481 185
R1093 VCC.n8401 VCC.n8400 185
R1094 VCC.n8517 VCC.n8401 185
R1095 VCC.n8538 VCC.n8537 185
R1096 VCC.n8539 VCC.n8538 185
R1097 VCC.n8536 VCC.n8389 185
R1098 VCC.n8540 VCC.n8389 185
R1099 VCC.n8520 VCC.n8519 185
R1100 VCC.n8519 VCC.n8518 185
R1101 VCC.n8549 VCC.n8390 185
R1102 VCC.n8430 VCC.n8429 185
R1103 VCC.n8428 VCC.n8427 185
R1104 VCC.n8458 VCC.n8428 185
R1105 VCC.n8461 VCC.n8460 185
R1106 VCC.n8460 VCC.n8459 185
R1107 VCC.n8416 VCC.n8415 185
R1108 VCC.n8483 VCC.n8416 185
R1109 VCC.n8543 VCC.n8365 185
R1110 VCC.n8541 VCC.n8365 185
R1111 VCC.n8364 VCC.n8363 185
R1112 VCC.n8593 VCC.n8364 185
R1113 VCC.n8614 VCC.n8613 185
R1114 VCC.n8614 VCC.n8350 185
R1115 VCC.n8333 VCC.n8332 185
R1116 VCC.n8332 VCC.n8331 185
R1117 VCC.n8651 VCC.n8650 185
R1118 VCC.n8650 VCC.n8649 185
R1119 VCC.n8670 VCC.n8669 185
R1120 VCC.n8671 VCC.n8670 185
R1121 VCC.n8620 VCC.n8619 185
R1122 VCC.n8619 VCC.n8618 185
R1123 VCC.n8597 VCC.n8596 185
R1124 VCC.n8596 VCC.n8595 185
R1125 VCC.n8615 VCC.n8348 185
R1126 VCC.n8616 VCC.n8615 185
R1127 VCC.n8330 VCC.n8329 185
R1128 VCC.n8648 VCC.n8330 185
R1129 VCC.n8315 VCC.n8314 185
R1130 VCC.n8545 VCC.n8544 185
R1131 VCC.n8545 VCC.n8542 185
R1132 VCC.n229 VCC.n227 96.8274
R1133 VCC.n289 VCC.n142 96.8274
R1134 VCC.n360 VCC.n108 96.8274
R1135 VCC.n396 VCC.n82 96.8274
R1136 VCC.n781 VCC.n779 96.8274
R1137 VCC.n841 VCC.n694 96.8274
R1138 VCC.n912 VCC.n660 96.8274
R1139 VCC.n948 VCC.n634 96.8274
R1140 VCC.n1469 VCC.n1217 96.8274
R1141 VCC.n1505 VCC.n1191 96.8274
R1142 VCC.n1339 VCC.n1337 96.8274
R1143 VCC.n1399 VCC.n1252 96.8274
R1144 VCC.n1890 VCC.n1888 96.8274
R1145 VCC.n1950 VCC.n1803 96.8274
R1146 VCC.n2021 VCC.n1769 96.8274
R1147 VCC.n2057 VCC.n1743 96.8274
R1148 VCC.n2578 VCC.n2326 96.8274
R1149 VCC.n2614 VCC.n2300 96.8274
R1150 VCC.n2448 VCC.n2446 96.8274
R1151 VCC.n2508 VCC.n2361 96.8274
R1152 VCC.n2999 VCC.n2997 96.8274
R1153 VCC.n3059 VCC.n2912 96.8274
R1154 VCC.n3130 VCC.n2878 96.8274
R1155 VCC.n3166 VCC.n2852 96.8274
R1156 VCC.n3687 VCC.n3435 96.8274
R1157 VCC.n3723 VCC.n3409 96.8274
R1158 VCC.n3557 VCC.n3555 96.8274
R1159 VCC.n3617 VCC.n3470 96.8274
R1160 VCC.n4108 VCC.n4106 96.8274
R1161 VCC.n4168 VCC.n4021 96.8274
R1162 VCC.n4239 VCC.n3987 96.8274
R1163 VCC.n4275 VCC.n3961 96.8274
R1164 VCC.n4796 VCC.n4544 96.8274
R1165 VCC.n4832 VCC.n4518 96.8274
R1166 VCC.n4666 VCC.n4664 96.8274
R1167 VCC.n4726 VCC.n4579 96.8274
R1168 VCC.n5217 VCC.n5215 96.8274
R1169 VCC.n5277 VCC.n5130 96.8274
R1170 VCC.n5348 VCC.n5096 96.8274
R1171 VCC.n5384 VCC.n5070 96.8274
R1172 VCC.n5904 VCC.n5652 96.8274
R1173 VCC.n5940 VCC.n5626 96.8274
R1174 VCC.n5774 VCC.n5772 96.8274
R1175 VCC.n5834 VCC.n5687 96.8274
R1176 VCC.n6324 VCC.n6322 96.8274
R1177 VCC.n6384 VCC.n6237 96.8274
R1178 VCC.n6455 VCC.n6203 96.8274
R1179 VCC.n6491 VCC.n6177 96.8274
R1180 VCC.n7011 VCC.n6759 96.8274
R1181 VCC.n7047 VCC.n6733 96.8274
R1182 VCC.n6881 VCC.n6879 96.8274
R1183 VCC.n6941 VCC.n6794 96.8274
R1184 VCC.n7431 VCC.n7429 96.8274
R1185 VCC.n7491 VCC.n7344 96.8274
R1186 VCC.n7562 VCC.n7310 96.8274
R1187 VCC.n7598 VCC.n7284 96.8274
R1188 VCC.n8118 VCC.n7866 96.8274
R1189 VCC.n8154 VCC.n7840 96.8274
R1190 VCC.n7988 VCC.n7986 96.8274
R1191 VCC.n8048 VCC.n7901 96.8274
R1192 VCC.n8482 VCC.n8417 96.8274
R1193 VCC.n8518 VCC.n8391 96.8274
R1194 VCC.n266 VCC.n153 95.0005
R1195 VCC.n267 VCC.n266 95.0005
R1196 VCC.n362 VCC.n93 95.0005
R1197 VCC.n394 VCC.n93 95.0005
R1198 VCC.n818 VCC.n705 95.0005
R1199 VCC.n819 VCC.n818 95.0005
R1200 VCC.n914 VCC.n645 95.0005
R1201 VCC.n946 VCC.n645 95.0005
R1202 VCC.n1471 VCC.n1202 95.0005
R1203 VCC.n1503 VCC.n1202 95.0005
R1204 VCC.n1376 VCC.n1263 95.0005
R1205 VCC.n1377 VCC.n1376 95.0005
R1206 VCC.n1927 VCC.n1814 95.0005
R1207 VCC.n1928 VCC.n1927 95.0005
R1208 VCC.n2023 VCC.n1754 95.0005
R1209 VCC.n2055 VCC.n1754 95.0005
R1210 VCC.n2580 VCC.n2311 95.0005
R1211 VCC.n2612 VCC.n2311 95.0005
R1212 VCC.n2485 VCC.n2372 95.0005
R1213 VCC.n2486 VCC.n2485 95.0005
R1214 VCC.n3036 VCC.n2923 95.0005
R1215 VCC.n3037 VCC.n3036 95.0005
R1216 VCC.n3132 VCC.n2863 95.0005
R1217 VCC.n3164 VCC.n2863 95.0005
R1218 VCC.n3689 VCC.n3420 95.0005
R1219 VCC.n3721 VCC.n3420 95.0005
R1220 VCC.n3594 VCC.n3481 95.0005
R1221 VCC.n3595 VCC.n3594 95.0005
R1222 VCC.n4145 VCC.n4032 95.0005
R1223 VCC.n4146 VCC.n4145 95.0005
R1224 VCC.n4241 VCC.n3972 95.0005
R1225 VCC.n4273 VCC.n3972 95.0005
R1226 VCC.n4798 VCC.n4529 95.0005
R1227 VCC.n4830 VCC.n4529 95.0005
R1228 VCC.n4703 VCC.n4590 95.0005
R1229 VCC.n4704 VCC.n4703 95.0005
R1230 VCC.n5254 VCC.n5141 95.0005
R1231 VCC.n5255 VCC.n5254 95.0005
R1232 VCC.n5350 VCC.n5081 95.0005
R1233 VCC.n5382 VCC.n5081 95.0005
R1234 VCC.n5906 VCC.n5637 95.0005
R1235 VCC.n5938 VCC.n5637 95.0005
R1236 VCC.n5811 VCC.n5698 95.0005
R1237 VCC.n5812 VCC.n5811 95.0005
R1238 VCC.n6361 VCC.n6248 95.0005
R1239 VCC.n6362 VCC.n6361 95.0005
R1240 VCC.n6457 VCC.n6188 95.0005
R1241 VCC.n6489 VCC.n6188 95.0005
R1242 VCC.n7013 VCC.n6744 95.0005
R1243 VCC.n7045 VCC.n6744 95.0005
R1244 VCC.n6918 VCC.n6805 95.0005
R1245 VCC.n6919 VCC.n6918 95.0005
R1246 VCC.n7468 VCC.n7355 95.0005
R1247 VCC.n7469 VCC.n7468 95.0005
R1248 VCC.n7564 VCC.n7295 95.0005
R1249 VCC.n7596 VCC.n7295 95.0005
R1250 VCC.n8120 VCC.n7851 95.0005
R1251 VCC.n8152 VCC.n7851 95.0005
R1252 VCC.n8025 VCC.n7912 95.0005
R1253 VCC.n8026 VCC.n8025 95.0005
R1254 VCC.n8484 VCC.n8402 95.0005
R1255 VCC.n8516 VCC.n8402 95.0005
R1256 VCC.n473 VCC.n472 93.2412
R1257 VCC.n495 VCC.n494 93.2412
R1258 VCC.n496 VCC.n495 93.2412
R1259 VCC.n547 VCC.n5 93.2412
R1260 VCC.n1025 VCC.n1024 93.2412
R1261 VCC.n1047 VCC.n1046 93.2412
R1262 VCC.n1048 VCC.n1047 93.2412
R1263 VCC.n1101 VCC.n559 93.2412
R1264 VCC.n1585 VCC.n1581 93.2412
R1265 VCC.n1583 VCC.n1143 93.2412
R1266 VCC.n1619 VCC.n1143 93.2412
R1267 VCC.n1653 VCC.n1652 93.2412
R1268 VCC.n2134 VCC.n2133 93.2412
R1269 VCC.n2156 VCC.n2155 93.2412
R1270 VCC.n2157 VCC.n2156 93.2412
R1271 VCC.n2210 VCC.n1668 93.2412
R1272 VCC.n2694 VCC.n2690 93.2412
R1273 VCC.n2692 VCC.n2252 93.2412
R1274 VCC.n2728 VCC.n2252 93.2412
R1275 VCC.n2762 VCC.n2761 93.2412
R1276 VCC.n3243 VCC.n3242 93.2412
R1277 VCC.n3265 VCC.n3264 93.2412
R1278 VCC.n3266 VCC.n3265 93.2412
R1279 VCC.n3319 VCC.n2777 93.2412
R1280 VCC.n3803 VCC.n3799 93.2412
R1281 VCC.n3801 VCC.n3361 93.2412
R1282 VCC.n3837 VCC.n3361 93.2412
R1283 VCC.n3871 VCC.n3870 93.2412
R1284 VCC.n4352 VCC.n4351 93.2412
R1285 VCC.n4374 VCC.n4373 93.2412
R1286 VCC.n4375 VCC.n4374 93.2412
R1287 VCC.n4428 VCC.n3886 93.2412
R1288 VCC.n4912 VCC.n4908 93.2412
R1289 VCC.n4910 VCC.n4470 93.2412
R1290 VCC.n4946 VCC.n4470 93.2412
R1291 VCC.n4980 VCC.n4979 93.2412
R1292 VCC.n5461 VCC.n5460 93.2412
R1293 VCC.n5483 VCC.n5482 93.2412
R1294 VCC.n5484 VCC.n5483 93.2412
R1295 VCC.n5537 VCC.n4995 93.2412
R1296 VCC.n6020 VCC.n6016 93.2412
R1297 VCC.n6018 VCC.n5578 93.2412
R1298 VCC.n6054 VCC.n5578 93.2412
R1299 VCC.n6088 VCC.n6087 93.2412
R1300 VCC.n6568 VCC.n6567 93.2412
R1301 VCC.n6590 VCC.n6589 93.2412
R1302 VCC.n6591 VCC.n6590 93.2412
R1303 VCC.n6644 VCC.n6102 93.2412
R1304 VCC.n7127 VCC.n7123 93.2412
R1305 VCC.n7125 VCC.n6685 93.2412
R1306 VCC.n7161 VCC.n6685 93.2412
R1307 VCC.n7195 VCC.n7194 93.2412
R1308 VCC.n7675 VCC.n7674 93.2412
R1309 VCC.n7697 VCC.n7696 93.2412
R1310 VCC.n7698 VCC.n7697 93.2412
R1311 VCC.n7751 VCC.n7209 93.2412
R1312 VCC.n8234 VCC.n8230 93.2412
R1313 VCC.n8232 VCC.n7792 93.2412
R1314 VCC.n8268 VCC.n7792 93.2412
R1315 VCC.n8302 VCC.n8301 93.2412
R1316 VCC.n8595 VCC.n8594 93.2412
R1317 VCC.n8617 VCC.n8616 93.2412
R1318 VCC.n8618 VCC.n8617 93.2412
R1319 VCC.n8671 VCC.n8316 93.2412
R1320 VCC.n213 VCC.n194 92.5398
R1321 VCC.n333 VCC.n123 92.5398
R1322 VCC.n430 VCC.n79 92.5398
R1323 VCC.n765 VCC.n746 92.5398
R1324 VCC.n885 VCC.n675 92.5398
R1325 VCC.n982 VCC.n631 92.5398
R1326 VCC.n1442 VCC.n1232 92.5398
R1327 VCC.n1540 VCC.n1188 92.5398
R1328 VCC.n1323 VCC.n1304 92.5398
R1329 VCC.n1874 VCC.n1855 92.5398
R1330 VCC.n1994 VCC.n1784 92.5398
R1331 VCC.n2091 VCC.n1740 92.5398
R1332 VCC.n2551 VCC.n2341 92.5398
R1333 VCC.n2649 VCC.n2297 92.5398
R1334 VCC.n2432 VCC.n2413 92.5398
R1335 VCC.n2983 VCC.n2964 92.5398
R1336 VCC.n3103 VCC.n2893 92.5398
R1337 VCC.n3200 VCC.n2849 92.5398
R1338 VCC.n3660 VCC.n3450 92.5398
R1339 VCC.n3758 VCC.n3406 92.5398
R1340 VCC.n3541 VCC.n3522 92.5398
R1341 VCC.n4092 VCC.n4073 92.5398
R1342 VCC.n4212 VCC.n4002 92.5398
R1343 VCC.n4309 VCC.n3958 92.5398
R1344 VCC.n4769 VCC.n4559 92.5398
R1345 VCC.n4867 VCC.n4515 92.5398
R1346 VCC.n4650 VCC.n4631 92.5398
R1347 VCC.n5201 VCC.n5182 92.5398
R1348 VCC.n5321 VCC.n5111 92.5398
R1349 VCC.n5418 VCC.n5067 92.5398
R1350 VCC.n5877 VCC.n5667 92.5398
R1351 VCC.n5975 VCC.n5623 92.5398
R1352 VCC.n5758 VCC.n5739 92.5398
R1353 VCC.n6308 VCC.n6289 92.5398
R1354 VCC.n6428 VCC.n6218 92.5398
R1355 VCC.n6525 VCC.n6174 92.5398
R1356 VCC.n6984 VCC.n6774 92.5398
R1357 VCC.n7082 VCC.n6730 92.5398
R1358 VCC.n6865 VCC.n6846 92.5398
R1359 VCC.n7415 VCC.n7396 92.5398
R1360 VCC.n7535 VCC.n7325 92.5398
R1361 VCC.n7632 VCC.n7281 92.5398
R1362 VCC.n8091 VCC.n7881 92.5398
R1363 VCC.n8189 VCC.n7837 92.5398
R1364 VCC.n7972 VCC.n7953 92.5398
R1365 VCC.n8455 VCC.n8432 92.5398
R1366 VCC.n8552 VCC.n8388 92.5398
R1367 VCC.n265 VCC.n264 92.5005
R1368 VCC.n266 VCC.n265 92.5005
R1369 VCC.n385 VCC.n94 92.5005
R1370 VCC.n94 VCC.n93 92.5005
R1371 VCC.n817 VCC.n816 92.5005
R1372 VCC.n818 VCC.n817 92.5005
R1373 VCC.n937 VCC.n646 92.5005
R1374 VCC.n646 VCC.n645 92.5005
R1375 VCC.n1494 VCC.n1203 92.5005
R1376 VCC.n1203 VCC.n1202 92.5005
R1377 VCC.n1375 VCC.n1374 92.5005
R1378 VCC.n1376 VCC.n1375 92.5005
R1379 VCC.n1926 VCC.n1925 92.5005
R1380 VCC.n1927 VCC.n1926 92.5005
R1381 VCC.n2046 VCC.n1755 92.5005
R1382 VCC.n1755 VCC.n1754 92.5005
R1383 VCC.n2603 VCC.n2312 92.5005
R1384 VCC.n2312 VCC.n2311 92.5005
R1385 VCC.n2484 VCC.n2483 92.5005
R1386 VCC.n2485 VCC.n2484 92.5005
R1387 VCC.n3035 VCC.n3034 92.5005
R1388 VCC.n3036 VCC.n3035 92.5005
R1389 VCC.n3155 VCC.n2864 92.5005
R1390 VCC.n2864 VCC.n2863 92.5005
R1391 VCC.n3712 VCC.n3421 92.5005
R1392 VCC.n3421 VCC.n3420 92.5005
R1393 VCC.n3593 VCC.n3592 92.5005
R1394 VCC.n3594 VCC.n3593 92.5005
R1395 VCC.n4144 VCC.n4143 92.5005
R1396 VCC.n4145 VCC.n4144 92.5005
R1397 VCC.n4264 VCC.n3973 92.5005
R1398 VCC.n3973 VCC.n3972 92.5005
R1399 VCC.n4821 VCC.n4530 92.5005
R1400 VCC.n4530 VCC.n4529 92.5005
R1401 VCC.n4702 VCC.n4701 92.5005
R1402 VCC.n4703 VCC.n4702 92.5005
R1403 VCC.n5253 VCC.n5252 92.5005
R1404 VCC.n5254 VCC.n5253 92.5005
R1405 VCC.n5373 VCC.n5082 92.5005
R1406 VCC.n5082 VCC.n5081 92.5005
R1407 VCC.n5929 VCC.n5638 92.5005
R1408 VCC.n5638 VCC.n5637 92.5005
R1409 VCC.n5810 VCC.n5809 92.5005
R1410 VCC.n5811 VCC.n5810 92.5005
R1411 VCC.n6360 VCC.n6359 92.5005
R1412 VCC.n6361 VCC.n6360 92.5005
R1413 VCC.n6480 VCC.n6189 92.5005
R1414 VCC.n6189 VCC.n6188 92.5005
R1415 VCC.n7036 VCC.n6745 92.5005
R1416 VCC.n6745 VCC.n6744 92.5005
R1417 VCC.n6917 VCC.n6916 92.5005
R1418 VCC.n6918 VCC.n6917 92.5005
R1419 VCC.n7467 VCC.n7466 92.5005
R1420 VCC.n7468 VCC.n7467 92.5005
R1421 VCC.n7587 VCC.n7296 92.5005
R1422 VCC.n7296 VCC.n7295 92.5005
R1423 VCC.n8143 VCC.n7852 92.5005
R1424 VCC.n7852 VCC.n7851 92.5005
R1425 VCC.n8024 VCC.n8023 92.5005
R1426 VCC.n8025 VCC.n8024 92.5005
R1427 VCC.n8507 VCC.n8403 92.5005
R1428 VCC.n8403 VCC.n8402 92.5005
R1429 VCC.n211 VCC.t262 74.9043
R1430 VCC.n763 VCC.t305 74.9043
R1431 VCC.n1321 VCC.t4 74.9043
R1432 VCC.n1872 VCC.t208 74.9043
R1433 VCC.n2430 VCC.t226 74.9043
R1434 VCC.n2981 VCC.t185 74.9043
R1435 VCC.n3539 VCC.t287 74.9043
R1436 VCC.n4090 VCC.t73 74.9043
R1437 VCC.n4648 VCC.t56 74.9043
R1438 VCC.n5199 VCC.t140 74.9043
R1439 VCC.n5756 VCC.t53 74.9043
R1440 VCC.n6306 VCC.t59 74.9043
R1441 VCC.n6863 VCC.t41 74.9043
R1442 VCC.n7413 VCC.t12 74.9043
R1443 VCC.n7970 VCC.t78 74.9043
R1444 VCC.t248 VCC.n335 73.0774
R1445 VCC.t105 VCC.n887 73.0774
R1446 VCC.t138 VCC.n1444 73.0774
R1447 VCC.t50 VCC.n1996 73.0774
R1448 VCC.t195 VCC.n2553 73.0774
R1449 VCC.t292 VCC.n3105 73.0774
R1450 VCC.t178 VCC.n3662 73.0774
R1451 VCC.t202 VCC.n4214 73.0774
R1452 VCC.t159 VCC.n4771 73.0774
R1453 VCC.t233 VCC.n5323 73.0774
R1454 VCC.t191 VCC.n5879 73.0774
R1455 VCC.t15 VCC.n6430 73.0774
R1456 VCC.t156 VCC.n6986 73.0774
R1457 VCC.t279 VCC.n7537 73.0774
R1458 VCC.t215 VCC.n8093 73.0774
R1459 VCC.t152 VCC.n8457 73.0774
R1460 VCC.n293 VCC.t289 72.544
R1461 VCC.n845 VCC.t235 72.544
R1462 VCC.n1403 VCC.t149 72.544
R1463 VCC.n1954 VCC.t76 72.544
R1464 VCC.n2512 VCC.t32 72.544
R1465 VCC.n3063 VCC.t147 72.544
R1466 VCC.n3621 VCC.t311 72.544
R1467 VCC.n4172 VCC.t298 72.544
R1468 VCC.n4730 VCC.t175 72.544
R1469 VCC.n5281 VCC.t125 72.544
R1470 VCC.n5838 VCC.t259 72.544
R1471 VCC.n6388 VCC.t88 72.544
R1472 VCC.n6945 VCC.t82 72.544
R1473 VCC.n7495 VCC.t172 72.544
R1474 VCC.n8052 VCC.t206 72.544
R1475 VCC.t35 VCC.n525 70.3709
R1476 VCC.t284 VCC.n1077 70.3709
R1477 VCC.n1621 VCC.t134 70.3709
R1478 VCC.t2 VCC.n2186 70.3709
R1479 VCC.n2730 VCC.t45 70.3709
R1480 VCC.t198 VCC.n3295 70.3709
R1481 VCC.n3839 VCC.t274 70.3709
R1482 VCC.t99 VCC.n4404 70.3709
R1483 VCC.n4948 VCC.t264 70.3709
R1484 VCC.t116 VCC.n5513 70.3709
R1485 VCC.n6056 VCC.t8 70.3709
R1486 VCC.t237 VCC.n6620 70.3709
R1487 VCC.n7163 VCC.t85 70.3709
R1488 VCC.t308 VCC.n7727 70.3709
R1489 VCC.n8270 VCC.t39 70.3709
R1490 VCC.t294 VCC.n8647 70.3709
R1491 VCC.n470 VCC.t252 66.8524
R1492 VCC.n1022 VCC.t29 66.8524
R1493 VCC.t24 VCC.n1163 66.8524
R1494 VCC.n2131 VCC.t21 66.8524
R1495 VCC.t187 VCC.n2272 66.8524
R1496 VCC.n3240 VCC.t95 66.8524
R1497 VCC.t269 VCC.n3381 66.8524
R1498 VCC.n4349 VCC.t300 66.8524
R1499 VCC.t113 VCC.n4490 66.8524
R1500 VCC.n5458 VCC.t223 66.8524
R1501 VCC.t245 VCC.n5598 66.8524
R1502 VCC.n6565 VCC.t169 66.8524
R1503 VCC.t108 VCC.n6705 66.8524
R1504 VCC.n7672 VCC.t69 66.8524
R1505 VCC.t218 VCC.n7812 66.8524
R1506 VCC.n8592 VCC.t65 66.8524
R1507 VCC.n428 VCC.t102 65.7697
R1508 VCC.n980 VCC.t212 65.7697
R1509 VCC.n1538 VCC.t255 65.7697
R1510 VCC.n2089 VCC.t18 65.7697
R1511 VCC.n2647 VCC.t143 65.7697
R1512 VCC.n3198 VCC.t230 65.7697
R1513 VCC.n3756 VCC.t181 65.7697
R1514 VCC.n4307 VCC.t91 65.7697
R1515 VCC.n4865 VCC.t123 65.7697
R1516 VCC.n5416 VCC.t161 65.7697
R1517 VCC.n5973 VCC.t242 65.7697
R1518 VCC.n6523 VCC.t165 65.7697
R1519 VCC.n7080 VCC.t130 65.7697
R1520 VCC.n7630 VCC.t63 65.7697
R1521 VCC.n8187 VCC.t120 65.7697
R1522 VCC.n8550 VCC.t276 65.7697
R1523 VCC.n293 VCC.n292 50.4194
R1524 VCC.n845 VCC.n844 50.4194
R1525 VCC.n1403 VCC.n1402 50.4194
R1526 VCC.n1954 VCC.n1953 50.4194
R1527 VCC.n2512 VCC.n2511 50.4194
R1528 VCC.n3063 VCC.n3062 50.4194
R1529 VCC.n3621 VCC.n3620 50.4194
R1530 VCC.n4172 VCC.n4171 50.4194
R1531 VCC.n4730 VCC.n4729 50.4194
R1532 VCC.n5281 VCC.n5280 50.4194
R1533 VCC.n5838 VCC.n5837 50.4194
R1534 VCC.n6388 VCC.n6387 50.4194
R1535 VCC.n6945 VCC.n6944 50.4194
R1536 VCC.n7495 VCC.n7494 50.4194
R1537 VCC.n8052 VCC.n8051 50.4194
R1538 VCC.n212 VCC.n182 50.3505
R1539 VCC.n230 VCC.n179 50.3505
R1540 VCC.n288 VCC.n143 50.3505
R1541 VCC.n334 VCC.n119 50.3505
R1542 VCC.n359 VCC.n109 50.3505
R1543 VCC.n397 VCC.n83 50.3505
R1544 VCC.n429 VCC.n80 50.3505
R1545 VCC.n764 VCC.n734 50.3505
R1546 VCC.n782 VCC.n731 50.3505
R1547 VCC.n840 VCC.n695 50.3505
R1548 VCC.n886 VCC.n671 50.3505
R1549 VCC.n911 VCC.n661 50.3505
R1550 VCC.n949 VCC.n635 50.3505
R1551 VCC.n981 VCC.n632 50.3505
R1552 VCC.n1443 VCC.n1228 50.3505
R1553 VCC.n1468 VCC.n1218 50.3505
R1554 VCC.n1506 VCC.n1192 50.3505
R1555 VCC.n1539 VCC.n1189 50.3505
R1556 VCC.n1322 VCC.n1292 50.3505
R1557 VCC.n1340 VCC.n1289 50.3505
R1558 VCC.n1398 VCC.n1253 50.3505
R1559 VCC.n1873 VCC.n1843 50.3505
R1560 VCC.n1891 VCC.n1840 50.3505
R1561 VCC.n1949 VCC.n1804 50.3505
R1562 VCC.n1995 VCC.n1780 50.3505
R1563 VCC.n2020 VCC.n1770 50.3505
R1564 VCC.n2058 VCC.n1744 50.3505
R1565 VCC.n2090 VCC.n1741 50.3505
R1566 VCC.n2552 VCC.n2337 50.3505
R1567 VCC.n2577 VCC.n2327 50.3505
R1568 VCC.n2615 VCC.n2301 50.3505
R1569 VCC.n2648 VCC.n2298 50.3505
R1570 VCC.n2431 VCC.n2401 50.3505
R1571 VCC.n2449 VCC.n2398 50.3505
R1572 VCC.n2507 VCC.n2362 50.3505
R1573 VCC.n2982 VCC.n2952 50.3505
R1574 VCC.n3000 VCC.n2949 50.3505
R1575 VCC.n3058 VCC.n2913 50.3505
R1576 VCC.n3104 VCC.n2889 50.3505
R1577 VCC.n3129 VCC.n2879 50.3505
R1578 VCC.n3167 VCC.n2853 50.3505
R1579 VCC.n3199 VCC.n2850 50.3505
R1580 VCC.n3661 VCC.n3446 50.3505
R1581 VCC.n3686 VCC.n3436 50.3505
R1582 VCC.n3724 VCC.n3410 50.3505
R1583 VCC.n3757 VCC.n3407 50.3505
R1584 VCC.n3540 VCC.n3510 50.3505
R1585 VCC.n3558 VCC.n3507 50.3505
R1586 VCC.n3616 VCC.n3471 50.3505
R1587 VCC.n4091 VCC.n4061 50.3505
R1588 VCC.n4109 VCC.n4058 50.3505
R1589 VCC.n4167 VCC.n4022 50.3505
R1590 VCC.n4213 VCC.n3998 50.3505
R1591 VCC.n4238 VCC.n3988 50.3505
R1592 VCC.n4276 VCC.n3962 50.3505
R1593 VCC.n4308 VCC.n3959 50.3505
R1594 VCC.n4770 VCC.n4555 50.3505
R1595 VCC.n4795 VCC.n4545 50.3505
R1596 VCC.n4833 VCC.n4519 50.3505
R1597 VCC.n4866 VCC.n4516 50.3505
R1598 VCC.n4649 VCC.n4619 50.3505
R1599 VCC.n4667 VCC.n4616 50.3505
R1600 VCC.n4725 VCC.n4580 50.3505
R1601 VCC.n5200 VCC.n5170 50.3505
R1602 VCC.n5218 VCC.n5167 50.3505
R1603 VCC.n5276 VCC.n5131 50.3505
R1604 VCC.n5322 VCC.n5107 50.3505
R1605 VCC.n5347 VCC.n5097 50.3505
R1606 VCC.n5385 VCC.n5071 50.3505
R1607 VCC.n5417 VCC.n5068 50.3505
R1608 VCC.n5878 VCC.n5663 50.3505
R1609 VCC.n5903 VCC.n5653 50.3505
R1610 VCC.n5941 VCC.n5627 50.3505
R1611 VCC.n5974 VCC.n5624 50.3505
R1612 VCC.n5757 VCC.n5727 50.3505
R1613 VCC.n5775 VCC.n5724 50.3505
R1614 VCC.n5833 VCC.n5688 50.3505
R1615 VCC.n6307 VCC.n6277 50.3505
R1616 VCC.n6325 VCC.n6274 50.3505
R1617 VCC.n6383 VCC.n6238 50.3505
R1618 VCC.n6429 VCC.n6214 50.3505
R1619 VCC.n6454 VCC.n6204 50.3505
R1620 VCC.n6492 VCC.n6178 50.3505
R1621 VCC.n6524 VCC.n6175 50.3505
R1622 VCC.n6985 VCC.n6770 50.3505
R1623 VCC.n7010 VCC.n6760 50.3505
R1624 VCC.n7048 VCC.n6734 50.3505
R1625 VCC.n7081 VCC.n6731 50.3505
R1626 VCC.n6864 VCC.n6834 50.3505
R1627 VCC.n6882 VCC.n6831 50.3505
R1628 VCC.n6940 VCC.n6795 50.3505
R1629 VCC.n7414 VCC.n7384 50.3505
R1630 VCC.n7432 VCC.n7381 50.3505
R1631 VCC.n7490 VCC.n7345 50.3505
R1632 VCC.n7536 VCC.n7321 50.3505
R1633 VCC.n7561 VCC.n7311 50.3505
R1634 VCC.n7599 VCC.n7285 50.3505
R1635 VCC.n7631 VCC.n7282 50.3505
R1636 VCC.n8092 VCC.n7877 50.3505
R1637 VCC.n8117 VCC.n7867 50.3505
R1638 VCC.n8155 VCC.n7841 50.3505
R1639 VCC.n8188 VCC.n7838 50.3505
R1640 VCC.n7971 VCC.n7941 50.3505
R1641 VCC.n7989 VCC.n7938 50.3505
R1642 VCC.n8047 VCC.n7902 50.3505
R1643 VCC.n8456 VCC.n8428 50.3505
R1644 VCC.n8481 VCC.n8418 50.3505
R1645 VCC.n8519 VCC.n8392 50.3505
R1646 VCC.n8551 VCC.n8389 50.3505
R1647 VCC.n265 VCC.n154 49.4005
R1648 VCC.n265 VCC.n152 49.4005
R1649 VCC.n363 VCC.n94 49.4005
R1650 VCC.n393 VCC.n94 49.4005
R1651 VCC.n817 VCC.n706 49.4005
R1652 VCC.n817 VCC.n704 49.4005
R1653 VCC.n915 VCC.n646 49.4005
R1654 VCC.n945 VCC.n646 49.4005
R1655 VCC.n1472 VCC.n1203 49.4005
R1656 VCC.n1502 VCC.n1203 49.4005
R1657 VCC.n1375 VCC.n1264 49.4005
R1658 VCC.n1375 VCC.n1262 49.4005
R1659 VCC.n1926 VCC.n1815 49.4005
R1660 VCC.n1926 VCC.n1813 49.4005
R1661 VCC.n2024 VCC.n1755 49.4005
R1662 VCC.n2054 VCC.n1755 49.4005
R1663 VCC.n2581 VCC.n2312 49.4005
R1664 VCC.n2611 VCC.n2312 49.4005
R1665 VCC.n2484 VCC.n2373 49.4005
R1666 VCC.n2484 VCC.n2371 49.4005
R1667 VCC.n3035 VCC.n2924 49.4005
R1668 VCC.n3035 VCC.n2922 49.4005
R1669 VCC.n3133 VCC.n2864 49.4005
R1670 VCC.n3163 VCC.n2864 49.4005
R1671 VCC.n3690 VCC.n3421 49.4005
R1672 VCC.n3720 VCC.n3421 49.4005
R1673 VCC.n3593 VCC.n3482 49.4005
R1674 VCC.n3593 VCC.n3480 49.4005
R1675 VCC.n4144 VCC.n4033 49.4005
R1676 VCC.n4144 VCC.n4031 49.4005
R1677 VCC.n4242 VCC.n3973 49.4005
R1678 VCC.n4272 VCC.n3973 49.4005
R1679 VCC.n4799 VCC.n4530 49.4005
R1680 VCC.n4829 VCC.n4530 49.4005
R1681 VCC.n4702 VCC.n4591 49.4005
R1682 VCC.n4702 VCC.n4589 49.4005
R1683 VCC.n5253 VCC.n5142 49.4005
R1684 VCC.n5253 VCC.n5140 49.4005
R1685 VCC.n5351 VCC.n5082 49.4005
R1686 VCC.n5381 VCC.n5082 49.4005
R1687 VCC.n5907 VCC.n5638 49.4005
R1688 VCC.n5937 VCC.n5638 49.4005
R1689 VCC.n5810 VCC.n5699 49.4005
R1690 VCC.n5810 VCC.n5697 49.4005
R1691 VCC.n6360 VCC.n6249 49.4005
R1692 VCC.n6360 VCC.n6247 49.4005
R1693 VCC.n6458 VCC.n6189 49.4005
R1694 VCC.n6488 VCC.n6189 49.4005
R1695 VCC.n7014 VCC.n6745 49.4005
R1696 VCC.n7044 VCC.n6745 49.4005
R1697 VCC.n6917 VCC.n6806 49.4005
R1698 VCC.n6917 VCC.n6804 49.4005
R1699 VCC.n7467 VCC.n7356 49.4005
R1700 VCC.n7467 VCC.n7354 49.4005
R1701 VCC.n7565 VCC.n7296 49.4005
R1702 VCC.n7595 VCC.n7296 49.4005
R1703 VCC.n8121 VCC.n7852 49.4005
R1704 VCC.n8151 VCC.n7852 49.4005
R1705 VCC.n8024 VCC.n7913 49.4005
R1706 VCC.n8024 VCC.n7911 49.4005
R1707 VCC.n8485 VCC.n8403 49.4005
R1708 VCC.n8515 VCC.n8403 49.4005
R1709 VCC.n469 VCC.n56 43.1576
R1710 VCC.n474 VCC.n42 43.1576
R1711 VCC.n493 VCC.n40 43.1576
R1712 VCC.n497 VCC.n40 43.1576
R1713 VCC.n524 VCC.n21 43.1576
R1714 VCC.n546 VCC.n6 43.1576
R1715 VCC.n1021 VCC.n608 43.1576
R1716 VCC.n1026 VCC.n594 43.1576
R1717 VCC.n1045 VCC.n592 43.1576
R1718 VCC.n1049 VCC.n592 43.1576
R1719 VCC.n1076 VCC.n573 43.1576
R1720 VCC.n1100 VCC.n560 43.1576
R1721 VCC.n1530 VCC.n1164 43.1576
R1722 VCC.n1586 VCC.n1161 43.1576
R1723 VCC.n1582 VCC.n1144 43.1576
R1724 VCC.n1618 VCC.n1144 43.1576
R1725 VCC.n1622 VCC.n1115 43.1576
R1726 VCC.n1654 VCC.n1113 43.1576
R1727 VCC.n2130 VCC.n1717 43.1576
R1728 VCC.n2135 VCC.n1703 43.1576
R1729 VCC.n2154 VCC.n1701 43.1576
R1730 VCC.n2158 VCC.n1701 43.1576
R1731 VCC.n2185 VCC.n1682 43.1576
R1732 VCC.n2209 VCC.n1669 43.1576
R1733 VCC.n2639 VCC.n2273 43.1576
R1734 VCC.n2695 VCC.n2270 43.1576
R1735 VCC.n2691 VCC.n2253 43.1576
R1736 VCC.n2727 VCC.n2253 43.1576
R1737 VCC.n2731 VCC.n2224 43.1576
R1738 VCC.n2763 VCC.n2222 43.1576
R1739 VCC.n3239 VCC.n2826 43.1576
R1740 VCC.n3244 VCC.n2812 43.1576
R1741 VCC.n3263 VCC.n2810 43.1576
R1742 VCC.n3267 VCC.n2810 43.1576
R1743 VCC.n3294 VCC.n2791 43.1576
R1744 VCC.n3318 VCC.n2778 43.1576
R1745 VCC.n3748 VCC.n3382 43.1576
R1746 VCC.n3804 VCC.n3379 43.1576
R1747 VCC.n3800 VCC.n3362 43.1576
R1748 VCC.n3836 VCC.n3362 43.1576
R1749 VCC.n3840 VCC.n3333 43.1576
R1750 VCC.n3872 VCC.n3331 43.1576
R1751 VCC.n4348 VCC.n3935 43.1576
R1752 VCC.n4353 VCC.n3921 43.1576
R1753 VCC.n4372 VCC.n3919 43.1576
R1754 VCC.n4376 VCC.n3919 43.1576
R1755 VCC.n4403 VCC.n3900 43.1576
R1756 VCC.n4427 VCC.n3887 43.1576
R1757 VCC.n4857 VCC.n4491 43.1576
R1758 VCC.n4913 VCC.n4488 43.1576
R1759 VCC.n4909 VCC.n4471 43.1576
R1760 VCC.n4945 VCC.n4471 43.1576
R1761 VCC.n4949 VCC.n4442 43.1576
R1762 VCC.n4981 VCC.n4440 43.1576
R1763 VCC.n5457 VCC.n5044 43.1576
R1764 VCC.n5462 VCC.n5030 43.1576
R1765 VCC.n5481 VCC.n5028 43.1576
R1766 VCC.n5485 VCC.n5028 43.1576
R1767 VCC.n5512 VCC.n5009 43.1576
R1768 VCC.n5536 VCC.n4996 43.1576
R1769 VCC.n5965 VCC.n5599 43.1576
R1770 VCC.n6021 VCC.n5596 43.1576
R1771 VCC.n6017 VCC.n5579 43.1576
R1772 VCC.n6053 VCC.n5579 43.1576
R1773 VCC.n6057 VCC.n5550 43.1576
R1774 VCC.n6089 VCC.n5548 43.1576
R1775 VCC.n6564 VCC.n6151 43.1576
R1776 VCC.n6569 VCC.n6137 43.1576
R1777 VCC.n6588 VCC.n6135 43.1576
R1778 VCC.n6592 VCC.n6135 43.1576
R1779 VCC.n6619 VCC.n6116 43.1576
R1780 VCC.n6643 VCC.n6103 43.1576
R1781 VCC.n7072 VCC.n6706 43.1576
R1782 VCC.n7128 VCC.n6703 43.1576
R1783 VCC.n7124 VCC.n6686 43.1576
R1784 VCC.n7160 VCC.n6686 43.1576
R1785 VCC.n7164 VCC.n6657 43.1576
R1786 VCC.n7196 VCC.n6655 43.1576
R1787 VCC.n7671 VCC.n7258 43.1576
R1788 VCC.n7676 VCC.n7244 43.1576
R1789 VCC.n7695 VCC.n7242 43.1576
R1790 VCC.n7699 VCC.n7242 43.1576
R1791 VCC.n7726 VCC.n7223 43.1576
R1792 VCC.n7750 VCC.n7210 43.1576
R1793 VCC.n8179 VCC.n7813 43.1576
R1794 VCC.n8235 VCC.n7810 43.1576
R1795 VCC.n8231 VCC.n7793 43.1576
R1796 VCC.n8267 VCC.n7793 43.1576
R1797 VCC.n8271 VCC.n7764 43.1576
R1798 VCC.n8303 VCC.n7762 43.1576
R1799 VCC.n8591 VCC.n8365 43.1576
R1800 VCC.n8596 VCC.n8351 43.1576
R1801 VCC.n8615 VCC.n8349 43.1576
R1802 VCC.n8619 VCC.n8349 43.1576
R1803 VCC.n8646 VCC.n8330 43.1576
R1804 VCC.n8670 VCC.n8317 43.1576
R1805 VCC.n548 VCC.n547 36.8662
R1806 VCC.n1102 VCC.n1101 36.8662
R1807 VCC.n1653 VCC.n1111 36.8662
R1808 VCC.n2211 VCC.n2210 36.8662
R1809 VCC.n2762 VCC.n2220 36.8662
R1810 VCC.n3320 VCC.n3319 36.8662
R1811 VCC.n3871 VCC.n3329 36.8662
R1812 VCC.n4429 VCC.n4428 36.8662
R1813 VCC.n4980 VCC.n4438 36.8662
R1814 VCC.n5538 VCC.n5537 36.8662
R1815 VCC.n6088 VCC.n5546 36.8662
R1816 VCC.n6645 VCC.n6644 36.8662
R1817 VCC.n7195 VCC.n6653 36.8662
R1818 VCC.n7752 VCC.n7751 36.8662
R1819 VCC.n8302 VCC.n7760 36.8662
R1820 VCC.n8672 VCC.n8671 36.8662
R1821 VCC.n446 VCC.t103 35.5869
R1822 VCC.n998 VCC.t213 35.5869
R1823 VCC.n1556 VCC.t256 35.5869
R1824 VCC.n2107 VCC.t19 35.5869
R1825 VCC.n2665 VCC.t144 35.5869
R1826 VCC.n3216 VCC.t231 35.5869
R1827 VCC.n3774 VCC.t182 35.5869
R1828 VCC.n4325 VCC.t92 35.5869
R1829 VCC.n4883 VCC.t124 35.5869
R1830 VCC.n5434 VCC.t162 35.5869
R1831 VCC.n5991 VCC.t243 35.5869
R1832 VCC.n6541 VCC.t166 35.5869
R1833 VCC.n7098 VCC.t131 35.5869
R1834 VCC.n7648 VCC.t64 35.5869
R1835 VCC.n8205 VCC.t121 35.5869
R1836 VCC.n8568 VCC.t277 35.5869
R1837 VCC.n11 VCC.t36 34.994
R1838 VCC.n1091 VCC.t285 34.994
R1839 VCC.n1640 VCC.t135 34.994
R1840 VCC.n2200 VCC.t3 34.994
R1841 VCC.n2749 VCC.t46 34.994
R1842 VCC.n3309 VCC.t199 34.994
R1843 VCC.n3858 VCC.t275 34.994
R1844 VCC.n4418 VCC.t100 34.994
R1845 VCC.n4967 VCC.t265 34.994
R1846 VCC.n5527 VCC.t117 34.994
R1847 VCC.n6075 VCC.t9 34.994
R1848 VCC.n6634 VCC.t238 34.994
R1849 VCC.n7182 VCC.t86 34.994
R1850 VCC.n7741 VCC.t309 34.994
R1851 VCC.n8289 VCC.t40 34.994
R1852 VCC.n8661 VCC.t295 34.994
R1853 VCC.n52 VCC.t253 34.9892
R1854 VCC.n604 VCC.t30 34.9892
R1855 VCC.n1157 VCC.t25 34.9892
R1856 VCC.n1713 VCC.t22 34.9892
R1857 VCC.n2266 VCC.t188 34.9892
R1858 VCC.n2822 VCC.t96 34.9892
R1859 VCC.n3375 VCC.t270 34.9892
R1860 VCC.n3931 VCC.t301 34.9892
R1861 VCC.n4484 VCC.t114 34.9892
R1862 VCC.n5040 VCC.t224 34.9892
R1863 VCC.n5592 VCC.t246 34.9892
R1864 VCC.n6147 VCC.t170 34.9892
R1865 VCC.n6699 VCC.t109 34.9892
R1866 VCC.n7254 VCC.t70 34.9892
R1867 VCC.n7806 VCC.t219 34.9892
R1868 VCC.n8361 VCC.t66 34.9892
R1869 VCC.n311 VCC.t290 34.9619
R1870 VCC.n863 VCC.t236 34.9619
R1871 VCC.n1421 VCC.t150 34.9619
R1872 VCC.n1972 VCC.t77 34.9619
R1873 VCC.n2530 VCC.t33 34.9619
R1874 VCC.n3081 VCC.t148 34.9619
R1875 VCC.n3639 VCC.t312 34.9619
R1876 VCC.n4190 VCC.t299 34.9619
R1877 VCC.n4748 VCC.t176 34.9619
R1878 VCC.n5299 VCC.t126 34.9619
R1879 VCC.n5856 VCC.t260 34.9619
R1880 VCC.n6406 VCC.t89 34.9619
R1881 VCC.n6963 VCC.t83 34.9619
R1882 VCC.n7513 VCC.t173 34.9619
R1883 VCC.n8070 VCC.t207 34.9619
R1884 VCC.n112 VCC.t249 34.945
R1885 VCC.n664 VCC.t106 34.945
R1886 VCC.n1221 VCC.t139 34.945
R1887 VCC.n1773 VCC.t51 34.945
R1888 VCC.n2330 VCC.t196 34.945
R1889 VCC.n2882 VCC.t293 34.945
R1890 VCC.n3439 VCC.t179 34.945
R1891 VCC.n3991 VCC.t203 34.945
R1892 VCC.n4548 VCC.t160 34.945
R1893 VCC.n5100 VCC.t234 34.945
R1894 VCC.n5656 VCC.t192 34.945
R1895 VCC.n6207 VCC.t16 34.945
R1896 VCC.n6763 VCC.t157 34.945
R1897 VCC.n7314 VCC.t280 34.945
R1898 VCC.n7870 VCC.t216 34.945
R1899 VCC.n8421 VCC.t153 34.945
R1900 VCC.n237 VCC.t263 34.9423
R1901 VCC.n789 VCC.t306 34.9423
R1902 VCC.n1347 VCC.t5 34.9423
R1903 VCC.n1898 VCC.t209 34.9423
R1904 VCC.n2456 VCC.t227 34.9423
R1905 VCC.n3007 VCC.t186 34.9423
R1906 VCC.n3565 VCC.t288 34.9423
R1907 VCC.n4116 VCC.t74 34.9423
R1908 VCC.n4674 VCC.t57 34.9423
R1909 VCC.n5225 VCC.t141 34.9423
R1910 VCC.n5782 VCC.t54 34.9423
R1911 VCC.n6332 VCC.t60 34.9423
R1912 VCC.n6889 VCC.t42 34.9423
R1913 VCC.n7439 VCC.t13 34.9423
R1914 VCC.n7996 VCC.t79 34.9423
R1915 VCC.n291 VCC.t289 32.8851
R1916 VCC.n843 VCC.t235 32.8851
R1917 VCC.n1401 VCC.t149 32.8851
R1918 VCC.n1952 VCC.t76 32.8851
R1919 VCC.n2510 VCC.t32 32.8851
R1920 VCC.n3061 VCC.t147 32.8851
R1921 VCC.n3619 VCC.t311 32.8851
R1922 VCC.n4170 VCC.t298 32.8851
R1923 VCC.n4728 VCC.t175 32.8851
R1924 VCC.n5279 VCC.t125 32.8851
R1925 VCC.n5836 VCC.t259 32.8851
R1926 VCC.n6386 VCC.t88 32.8851
R1927 VCC.n6943 VCC.t82 32.8851
R1928 VCC.n7493 VCC.t172 32.8851
R1929 VCC.n8050 VCC.t206 32.8851
R1930 VCC.t102 VCC.n418 31.0582
R1931 VCC.t212 VCC.n970 31.0582
R1932 VCC.t255 VCC.n1527 31.0582
R1933 VCC.t18 VCC.n2079 31.0582
R1934 VCC.t143 VCC.n2636 31.0582
R1935 VCC.t230 VCC.n3188 31.0582
R1936 VCC.t181 VCC.n3745 31.0582
R1937 VCC.t91 VCC.n4297 31.0582
R1938 VCC.t123 VCC.n4854 31.0582
R1939 VCC.t161 VCC.n5406 31.0582
R1940 VCC.t242 VCC.n5962 31.0582
R1941 VCC.t165 VCC.n6513 31.0582
R1942 VCC.t130 VCC.n7069 31.0582
R1943 VCC.t63 VCC.n7620 31.0582
R1944 VCC.t120 VCC.n8176 31.0582
R1945 VCC.t276 VCC.n8540 31.0582
R1946 VCC.n228 VCC.n153 29.2313
R1947 VCC.n268 VCC.n267 29.2313
R1948 VCC.n362 VCC.n361 29.2313
R1949 VCC.n395 VCC.n394 29.2313
R1950 VCC.n780 VCC.n705 29.2313
R1951 VCC.n820 VCC.n819 29.2313
R1952 VCC.n914 VCC.n913 29.2313
R1953 VCC.n947 VCC.n946 29.2313
R1954 VCC.n1471 VCC.n1470 29.2313
R1955 VCC.n1504 VCC.n1503 29.2313
R1956 VCC.n1338 VCC.n1263 29.2313
R1957 VCC.n1378 VCC.n1377 29.2313
R1958 VCC.n1889 VCC.n1814 29.2313
R1959 VCC.n1929 VCC.n1928 29.2313
R1960 VCC.n2023 VCC.n2022 29.2313
R1961 VCC.n2056 VCC.n2055 29.2313
R1962 VCC.n2580 VCC.n2579 29.2313
R1963 VCC.n2613 VCC.n2612 29.2313
R1964 VCC.n2447 VCC.n2372 29.2313
R1965 VCC.n2487 VCC.n2486 29.2313
R1966 VCC.n2998 VCC.n2923 29.2313
R1967 VCC.n3038 VCC.n3037 29.2313
R1968 VCC.n3132 VCC.n3131 29.2313
R1969 VCC.n3165 VCC.n3164 29.2313
R1970 VCC.n3689 VCC.n3688 29.2313
R1971 VCC.n3722 VCC.n3721 29.2313
R1972 VCC.n3556 VCC.n3481 29.2313
R1973 VCC.n3596 VCC.n3595 29.2313
R1974 VCC.n4107 VCC.n4032 29.2313
R1975 VCC.n4147 VCC.n4146 29.2313
R1976 VCC.n4241 VCC.n4240 29.2313
R1977 VCC.n4274 VCC.n4273 29.2313
R1978 VCC.n4798 VCC.n4797 29.2313
R1979 VCC.n4831 VCC.n4830 29.2313
R1980 VCC.n4665 VCC.n4590 29.2313
R1981 VCC.n4705 VCC.n4704 29.2313
R1982 VCC.n5216 VCC.n5141 29.2313
R1983 VCC.n5256 VCC.n5255 29.2313
R1984 VCC.n5350 VCC.n5349 29.2313
R1985 VCC.n5383 VCC.n5382 29.2313
R1986 VCC.n5906 VCC.n5905 29.2313
R1987 VCC.n5939 VCC.n5938 29.2313
R1988 VCC.n5773 VCC.n5698 29.2313
R1989 VCC.n5813 VCC.n5812 29.2313
R1990 VCC.n6323 VCC.n6248 29.2313
R1991 VCC.n6363 VCC.n6362 29.2313
R1992 VCC.n6457 VCC.n6456 29.2313
R1993 VCC.n6490 VCC.n6489 29.2313
R1994 VCC.n7013 VCC.n7012 29.2313
R1995 VCC.n7046 VCC.n7045 29.2313
R1996 VCC.n6880 VCC.n6805 29.2313
R1997 VCC.n6920 VCC.n6919 29.2313
R1998 VCC.n7430 VCC.n7355 29.2313
R1999 VCC.n7470 VCC.n7469 29.2313
R2000 VCC.n7564 VCC.n7563 29.2313
R2001 VCC.n7597 VCC.n7596 29.2313
R2002 VCC.n8120 VCC.n8119 29.2313
R2003 VCC.n8153 VCC.n8152 29.2313
R2004 VCC.n7987 VCC.n7912 29.2313
R2005 VCC.n8027 VCC.n8026 29.2313
R2006 VCC.n8484 VCC.n8483 29.2313
R2007 VCC.n8517 VCC.n8516 29.2313
R2008 VCC.n419 VCC.t252 26.3894
R2009 VCC.n494 VCC.n41 26.3894
R2010 VCC.n496 VCC.n22 26.3894
R2011 VCC.n971 VCC.t29 26.3894
R2012 VCC.n1046 VCC.n593 26.3894
R2013 VCC.n1048 VCC.n574 26.3894
R2014 VCC.n1529 VCC.t24 26.3894
R2015 VCC.n1584 VCC.n1583 26.3894
R2016 VCC.n1620 VCC.n1619 26.3894
R2017 VCC.n2080 VCC.t21 26.3894
R2018 VCC.n2155 VCC.n1702 26.3894
R2019 VCC.n2157 VCC.n1683 26.3894
R2020 VCC.n2638 VCC.t187 26.3894
R2021 VCC.n2693 VCC.n2692 26.3894
R2022 VCC.n2729 VCC.n2728 26.3894
R2023 VCC.n3189 VCC.t95 26.3894
R2024 VCC.n3264 VCC.n2811 26.3894
R2025 VCC.n3266 VCC.n2792 26.3894
R2026 VCC.n3747 VCC.t269 26.3894
R2027 VCC.n3802 VCC.n3801 26.3894
R2028 VCC.n3838 VCC.n3837 26.3894
R2029 VCC.n4298 VCC.t300 26.3894
R2030 VCC.n4373 VCC.n3920 26.3894
R2031 VCC.n4375 VCC.n3901 26.3894
R2032 VCC.n4856 VCC.t113 26.3894
R2033 VCC.n4911 VCC.n4910 26.3894
R2034 VCC.n4947 VCC.n4946 26.3894
R2035 VCC.n5407 VCC.t223 26.3894
R2036 VCC.n5482 VCC.n5029 26.3894
R2037 VCC.n5484 VCC.n5010 26.3894
R2038 VCC.n5964 VCC.t245 26.3894
R2039 VCC.n6019 VCC.n6018 26.3894
R2040 VCC.n6055 VCC.n6054 26.3894
R2041 VCC.n6514 VCC.t169 26.3894
R2042 VCC.n6589 VCC.n6136 26.3894
R2043 VCC.n6591 VCC.n6117 26.3894
R2044 VCC.n7071 VCC.t108 26.3894
R2045 VCC.n7126 VCC.n7125 26.3894
R2046 VCC.n7162 VCC.n7161 26.3894
R2047 VCC.n7621 VCC.t69 26.3894
R2048 VCC.n7696 VCC.n7243 26.3894
R2049 VCC.n7698 VCC.n7224 26.3894
R2050 VCC.n8178 VCC.t218 26.3894
R2051 VCC.n8233 VCC.n8232 26.3894
R2052 VCC.n8269 VCC.n8268 26.3894
R2053 VCC.n8541 VCC.t65 26.3894
R2054 VCC.n8616 VCC.n8350 26.3894
R2055 VCC.n8618 VCC.n8331 26.3894
R2056 VCC.n227 VCC.n226 25.5774
R2057 VCC.n290 VCC.n289 25.5774
R2058 VCC.n337 VCC.n108 25.5774
R2059 VCC.n417 VCC.n82 25.5774
R2060 VCC.n779 VCC.n778 25.5774
R2061 VCC.n842 VCC.n841 25.5774
R2062 VCC.n889 VCC.n660 25.5774
R2063 VCC.n969 VCC.n634 25.5774
R2064 VCC.n1446 VCC.n1217 25.5774
R2065 VCC.n1526 VCC.n1191 25.5774
R2066 VCC.n1337 VCC.n1336 25.5774
R2067 VCC.n1400 VCC.n1399 25.5774
R2068 VCC.n1888 VCC.n1887 25.5774
R2069 VCC.n1951 VCC.n1950 25.5774
R2070 VCC.n1998 VCC.n1769 25.5774
R2071 VCC.n2078 VCC.n1743 25.5774
R2072 VCC.n2555 VCC.n2326 25.5774
R2073 VCC.n2635 VCC.n2300 25.5774
R2074 VCC.n2446 VCC.n2445 25.5774
R2075 VCC.n2509 VCC.n2508 25.5774
R2076 VCC.n2997 VCC.n2996 25.5774
R2077 VCC.n3060 VCC.n3059 25.5774
R2078 VCC.n3107 VCC.n2878 25.5774
R2079 VCC.n3187 VCC.n2852 25.5774
R2080 VCC.n3664 VCC.n3435 25.5774
R2081 VCC.n3744 VCC.n3409 25.5774
R2082 VCC.n3555 VCC.n3554 25.5774
R2083 VCC.n3618 VCC.n3617 25.5774
R2084 VCC.n4106 VCC.n4105 25.5774
R2085 VCC.n4169 VCC.n4168 25.5774
R2086 VCC.n4216 VCC.n3987 25.5774
R2087 VCC.n4296 VCC.n3961 25.5774
R2088 VCC.n4773 VCC.n4544 25.5774
R2089 VCC.n4853 VCC.n4518 25.5774
R2090 VCC.n4664 VCC.n4663 25.5774
R2091 VCC.n4727 VCC.n4726 25.5774
R2092 VCC.n5215 VCC.n5214 25.5774
R2093 VCC.n5278 VCC.n5277 25.5774
R2094 VCC.n5325 VCC.n5096 25.5774
R2095 VCC.n5405 VCC.n5070 25.5774
R2096 VCC.n5881 VCC.n5652 25.5774
R2097 VCC.n5961 VCC.n5626 25.5774
R2098 VCC.n5772 VCC.n5771 25.5774
R2099 VCC.n5835 VCC.n5834 25.5774
R2100 VCC.n6322 VCC.n6321 25.5774
R2101 VCC.n6385 VCC.n6384 25.5774
R2102 VCC.n6432 VCC.n6203 25.5774
R2103 VCC.n6512 VCC.n6177 25.5774
R2104 VCC.n6988 VCC.n6759 25.5774
R2105 VCC.n7068 VCC.n6733 25.5774
R2106 VCC.n6879 VCC.n6878 25.5774
R2107 VCC.n6942 VCC.n6941 25.5774
R2108 VCC.n7429 VCC.n7428 25.5774
R2109 VCC.n7492 VCC.n7491 25.5774
R2110 VCC.n7539 VCC.n7310 25.5774
R2111 VCC.n7619 VCC.n7284 25.5774
R2112 VCC.n8095 VCC.n7866 25.5774
R2113 VCC.n8175 VCC.n7840 25.5774
R2114 VCC.n7986 VCC.n7985 25.5774
R2115 VCC.n8049 VCC.n8048 25.5774
R2116 VCC.n8459 VCC.n8417 25.5774
R2117 VCC.n8539 VCC.n8391 25.5774
R2118 VCC.n336 VCC.t248 23.7505
R2119 VCC.n888 VCC.t105 23.7505
R2120 VCC.n1445 VCC.t138 23.7505
R2121 VCC.n1997 VCC.t50 23.7505
R2122 VCC.n2554 VCC.t195 23.7505
R2123 VCC.n3106 VCC.t292 23.7505
R2124 VCC.n3663 VCC.t178 23.7505
R2125 VCC.n4215 VCC.t202 23.7505
R2126 VCC.n4772 VCC.t159 23.7505
R2127 VCC.n5324 VCC.t233 23.7505
R2128 VCC.n5880 VCC.t191 23.7505
R2129 VCC.n6431 VCC.t15 23.7505
R2130 VCC.n6987 VCC.t156 23.7505
R2131 VCC.n7538 VCC.t279 23.7505
R2132 VCC.n8094 VCC.t215 23.7505
R2133 VCC.n8458 VCC.t152 23.7505
R2134 VCC.n473 VCC.n471 22.8709
R2135 VCC.n526 VCC.t35 22.8709
R2136 VCC.n527 VCC.n526 22.8709
R2137 VCC.n1025 VCC.n1023 22.8709
R2138 VCC.n1078 VCC.t284 22.8709
R2139 VCC.n1079 VCC.n1078 22.8709
R2140 VCC.n1581 VCC.n1580 22.8709
R2141 VCC.t134 VCC.n1114 22.8709
R2142 VCC.n1651 VCC.n1114 22.8709
R2143 VCC.n2134 VCC.n2132 22.8709
R2144 VCC.n2187 VCC.t2 22.8709
R2145 VCC.n2188 VCC.n2187 22.8709
R2146 VCC.n2690 VCC.n2689 22.8709
R2147 VCC.t45 VCC.n2223 22.8709
R2148 VCC.n2760 VCC.n2223 22.8709
R2149 VCC.n3243 VCC.n3241 22.8709
R2150 VCC.n3296 VCC.t198 22.8709
R2151 VCC.n3297 VCC.n3296 22.8709
R2152 VCC.n3799 VCC.n3798 22.8709
R2153 VCC.t274 VCC.n3332 22.8709
R2154 VCC.n3869 VCC.n3332 22.8709
R2155 VCC.n4352 VCC.n4350 22.8709
R2156 VCC.n4405 VCC.t99 22.8709
R2157 VCC.n4406 VCC.n4405 22.8709
R2158 VCC.n4908 VCC.n4907 22.8709
R2159 VCC.t264 VCC.n4441 22.8709
R2160 VCC.n4978 VCC.n4441 22.8709
R2161 VCC.n5461 VCC.n5459 22.8709
R2162 VCC.n5514 VCC.t116 22.8709
R2163 VCC.n5515 VCC.n5514 22.8709
R2164 VCC.n6016 VCC.n6015 22.8709
R2165 VCC.t8 VCC.n5549 22.8709
R2166 VCC.n6086 VCC.n5549 22.8709
R2167 VCC.n6568 VCC.n6566 22.8709
R2168 VCC.n6621 VCC.t237 22.8709
R2169 VCC.n6622 VCC.n6621 22.8709
R2170 VCC.n7123 VCC.n7122 22.8709
R2171 VCC.t85 VCC.n6656 22.8709
R2172 VCC.n7193 VCC.n6656 22.8709
R2173 VCC.n7675 VCC.n7673 22.8709
R2174 VCC.n7728 VCC.t308 22.8709
R2175 VCC.n7729 VCC.n7728 22.8709
R2176 VCC.n8230 VCC.n8229 22.8709
R2177 VCC.t39 VCC.n7763 22.8709
R2178 VCC.n8300 VCC.n7763 22.8709
R2179 VCC.n8595 VCC.n8593 22.8709
R2180 VCC.n8648 VCC.t294 22.8709
R2181 VCC.n8649 VCC.n8648 22.8709
R2182 VCC.n211 VCC.n210 21.9236
R2183 VCC.t262 VCC.n181 21.9236
R2184 VCC.n335 VCC.n120 21.9236
R2185 VCC.n428 VCC.n427 21.9236
R2186 VCC.n763 VCC.n762 21.9236
R2187 VCC.t305 VCC.n733 21.9236
R2188 VCC.n887 VCC.n672 21.9236
R2189 VCC.n980 VCC.n979 21.9236
R2190 VCC.n1444 VCC.n1229 21.9236
R2191 VCC.n1538 VCC.n1537 21.9236
R2192 VCC.n1321 VCC.n1320 21.9236
R2193 VCC.t4 VCC.n1291 21.9236
R2194 VCC.n1872 VCC.n1871 21.9236
R2195 VCC.t208 VCC.n1842 21.9236
R2196 VCC.n1996 VCC.n1781 21.9236
R2197 VCC.n2089 VCC.n2088 21.9236
R2198 VCC.n2553 VCC.n2338 21.9236
R2199 VCC.n2647 VCC.n2646 21.9236
R2200 VCC.n2430 VCC.n2429 21.9236
R2201 VCC.t226 VCC.n2400 21.9236
R2202 VCC.n2981 VCC.n2980 21.9236
R2203 VCC.t185 VCC.n2951 21.9236
R2204 VCC.n3105 VCC.n2890 21.9236
R2205 VCC.n3198 VCC.n3197 21.9236
R2206 VCC.n3662 VCC.n3447 21.9236
R2207 VCC.n3756 VCC.n3755 21.9236
R2208 VCC.n3539 VCC.n3538 21.9236
R2209 VCC.t287 VCC.n3509 21.9236
R2210 VCC.n4090 VCC.n4089 21.9236
R2211 VCC.t73 VCC.n4060 21.9236
R2212 VCC.n4214 VCC.n3999 21.9236
R2213 VCC.n4307 VCC.n4306 21.9236
R2214 VCC.n4771 VCC.n4556 21.9236
R2215 VCC.n4865 VCC.n4864 21.9236
R2216 VCC.n4648 VCC.n4647 21.9236
R2217 VCC.t56 VCC.n4618 21.9236
R2218 VCC.n5199 VCC.n5198 21.9236
R2219 VCC.t140 VCC.n5169 21.9236
R2220 VCC.n5323 VCC.n5108 21.9236
R2221 VCC.n5416 VCC.n5415 21.9236
R2222 VCC.n5879 VCC.n5664 21.9236
R2223 VCC.n5973 VCC.n5972 21.9236
R2224 VCC.n5756 VCC.n5755 21.9236
R2225 VCC.t53 VCC.n5726 21.9236
R2226 VCC.n6306 VCC.n6305 21.9236
R2227 VCC.t59 VCC.n6276 21.9236
R2228 VCC.n6430 VCC.n6215 21.9236
R2229 VCC.n6523 VCC.n6522 21.9236
R2230 VCC.n6986 VCC.n6771 21.9236
R2231 VCC.n7080 VCC.n7079 21.9236
R2232 VCC.n6863 VCC.n6862 21.9236
R2233 VCC.t41 VCC.n6833 21.9236
R2234 VCC.n7413 VCC.n7412 21.9236
R2235 VCC.t12 VCC.n7383 21.9236
R2236 VCC.n7537 VCC.n7322 21.9236
R2237 VCC.n7630 VCC.n7629 21.9236
R2238 VCC.n8093 VCC.n7878 21.9236
R2239 VCC.n8187 VCC.n8186 21.9236
R2240 VCC.n7970 VCC.n7969 21.9236
R2241 VCC.t78 VCC.n7940 21.9236
R2242 VCC.n8457 VCC.n8429 21.9236
R2243 VCC.n8550 VCC.n8549 21.9236
R2244 VCC.n420 VCC.n419 19.3524
R2245 VCC.n972 VCC.n971 19.3524
R2246 VCC.n1529 VCC.n1528 19.3524
R2247 VCC.n2081 VCC.n2080 19.3524
R2248 VCC.n2638 VCC.n2637 19.3524
R2249 VCC.n3190 VCC.n3189 19.3524
R2250 VCC.n3747 VCC.n3746 19.3524
R2251 VCC.n4299 VCC.n4298 19.3524
R2252 VCC.n4856 VCC.n4855 19.3524
R2253 VCC.n5408 VCC.n5407 19.3524
R2254 VCC.n5964 VCC.n5963 19.3524
R2255 VCC.n6515 VCC.n6514 19.3524
R2256 VCC.n7071 VCC.n7070 19.3524
R2257 VCC.n7622 VCC.n7621 19.3524
R2258 VCC.n8178 VCC.n8177 19.3524
R2259 VCC.n8542 VCC.n8541 19.3524
R2260 VCC.n180 VCC.n154 15.2005
R2261 VCC.n269 VCC.n152 15.2005
R2262 VCC.n363 VCC.n107 15.2005
R2263 VCC.n393 VCC.n92 15.2005
R2264 VCC.n732 VCC.n706 15.2005
R2265 VCC.n821 VCC.n704 15.2005
R2266 VCC.n915 VCC.n659 15.2005
R2267 VCC.n945 VCC.n644 15.2005
R2268 VCC.n1472 VCC.n1216 15.2005
R2269 VCC.n1502 VCC.n1201 15.2005
R2270 VCC.n1290 VCC.n1264 15.2005
R2271 VCC.n1379 VCC.n1262 15.2005
R2272 VCC.n1841 VCC.n1815 15.2005
R2273 VCC.n1930 VCC.n1813 15.2005
R2274 VCC.n2024 VCC.n1768 15.2005
R2275 VCC.n2054 VCC.n1753 15.2005
R2276 VCC.n2581 VCC.n2325 15.2005
R2277 VCC.n2611 VCC.n2310 15.2005
R2278 VCC.n2399 VCC.n2373 15.2005
R2279 VCC.n2488 VCC.n2371 15.2005
R2280 VCC.n2950 VCC.n2924 15.2005
R2281 VCC.n3039 VCC.n2922 15.2005
R2282 VCC.n3133 VCC.n2877 15.2005
R2283 VCC.n3163 VCC.n2862 15.2005
R2284 VCC.n3690 VCC.n3434 15.2005
R2285 VCC.n3720 VCC.n3419 15.2005
R2286 VCC.n3508 VCC.n3482 15.2005
R2287 VCC.n3597 VCC.n3480 15.2005
R2288 VCC.n4059 VCC.n4033 15.2005
R2289 VCC.n4148 VCC.n4031 15.2005
R2290 VCC.n4242 VCC.n3986 15.2005
R2291 VCC.n4272 VCC.n3971 15.2005
R2292 VCC.n4799 VCC.n4543 15.2005
R2293 VCC.n4829 VCC.n4528 15.2005
R2294 VCC.n4617 VCC.n4591 15.2005
R2295 VCC.n4706 VCC.n4589 15.2005
R2296 VCC.n5168 VCC.n5142 15.2005
R2297 VCC.n5257 VCC.n5140 15.2005
R2298 VCC.n5351 VCC.n5095 15.2005
R2299 VCC.n5381 VCC.n5080 15.2005
R2300 VCC.n5907 VCC.n5651 15.2005
R2301 VCC.n5937 VCC.n5636 15.2005
R2302 VCC.n5725 VCC.n5699 15.2005
R2303 VCC.n5814 VCC.n5697 15.2005
R2304 VCC.n6275 VCC.n6249 15.2005
R2305 VCC.n6364 VCC.n6247 15.2005
R2306 VCC.n6458 VCC.n6202 15.2005
R2307 VCC.n6488 VCC.n6187 15.2005
R2308 VCC.n7014 VCC.n6758 15.2005
R2309 VCC.n7044 VCC.n6743 15.2005
R2310 VCC.n6832 VCC.n6806 15.2005
R2311 VCC.n6921 VCC.n6804 15.2005
R2312 VCC.n7382 VCC.n7356 15.2005
R2313 VCC.n7471 VCC.n7354 15.2005
R2314 VCC.n7565 VCC.n7309 15.2005
R2315 VCC.n7595 VCC.n7294 15.2005
R2316 VCC.n8121 VCC.n7865 15.2005
R2317 VCC.n8151 VCC.n7850 15.2005
R2318 VCC.n7939 VCC.n7913 15.2005
R2319 VCC.n8028 VCC.n7911 15.2005
R2320 VCC.n8485 VCC.n8416 15.2005
R2321 VCC.n8515 VCC.n8401 15.2005
R2322 VCC.n225 VCC.n179 13.3005
R2323 VCC.n288 VCC.n140 13.3005
R2324 VCC.n338 VCC.n109 13.3005
R2325 VCC.n416 VCC.n83 13.3005
R2326 VCC.n777 VCC.n731 13.3005
R2327 VCC.n840 VCC.n692 13.3005
R2328 VCC.n890 VCC.n661 13.3005
R2329 VCC.n968 VCC.n635 13.3005
R2330 VCC.n1447 VCC.n1218 13.3005
R2331 VCC.n1525 VCC.n1192 13.3005
R2332 VCC.n1335 VCC.n1289 13.3005
R2333 VCC.n1398 VCC.n1250 13.3005
R2334 VCC.n1886 VCC.n1840 13.3005
R2335 VCC.n1949 VCC.n1801 13.3005
R2336 VCC.n1999 VCC.n1770 13.3005
R2337 VCC.n2077 VCC.n1744 13.3005
R2338 VCC.n2556 VCC.n2327 13.3005
R2339 VCC.n2634 VCC.n2301 13.3005
R2340 VCC.n2444 VCC.n2398 13.3005
R2341 VCC.n2507 VCC.n2359 13.3005
R2342 VCC.n2995 VCC.n2949 13.3005
R2343 VCC.n3058 VCC.n2910 13.3005
R2344 VCC.n3108 VCC.n2879 13.3005
R2345 VCC.n3186 VCC.n2853 13.3005
R2346 VCC.n3665 VCC.n3436 13.3005
R2347 VCC.n3743 VCC.n3410 13.3005
R2348 VCC.n3553 VCC.n3507 13.3005
R2349 VCC.n3616 VCC.n3468 13.3005
R2350 VCC.n4104 VCC.n4058 13.3005
R2351 VCC.n4167 VCC.n4019 13.3005
R2352 VCC.n4217 VCC.n3988 13.3005
R2353 VCC.n4295 VCC.n3962 13.3005
R2354 VCC.n4774 VCC.n4545 13.3005
R2355 VCC.n4852 VCC.n4519 13.3005
R2356 VCC.n4662 VCC.n4616 13.3005
R2357 VCC.n4725 VCC.n4577 13.3005
R2358 VCC.n5213 VCC.n5167 13.3005
R2359 VCC.n5276 VCC.n5128 13.3005
R2360 VCC.n5326 VCC.n5097 13.3005
R2361 VCC.n5404 VCC.n5071 13.3005
R2362 VCC.n5882 VCC.n5653 13.3005
R2363 VCC.n5960 VCC.n5627 13.3005
R2364 VCC.n5770 VCC.n5724 13.3005
R2365 VCC.n5833 VCC.n5685 13.3005
R2366 VCC.n6320 VCC.n6274 13.3005
R2367 VCC.n6383 VCC.n6235 13.3005
R2368 VCC.n6433 VCC.n6204 13.3005
R2369 VCC.n6511 VCC.n6178 13.3005
R2370 VCC.n6989 VCC.n6760 13.3005
R2371 VCC.n7067 VCC.n6734 13.3005
R2372 VCC.n6877 VCC.n6831 13.3005
R2373 VCC.n6940 VCC.n6792 13.3005
R2374 VCC.n7427 VCC.n7381 13.3005
R2375 VCC.n7490 VCC.n7342 13.3005
R2376 VCC.n7540 VCC.n7311 13.3005
R2377 VCC.n7618 VCC.n7285 13.3005
R2378 VCC.n8096 VCC.n7867 13.3005
R2379 VCC.n8174 VCC.n7841 13.3005
R2380 VCC.n7984 VCC.n7938 13.3005
R2381 VCC.n8047 VCC.n7899 13.3005
R2382 VCC.n8460 VCC.n8418 13.3005
R2383 VCC.n8538 VCC.n8392 13.3005
R2384 VCC.n493 VCC.n492 12.2148
R2385 VCC.n497 VCC.n23 12.2148
R2386 VCC.n1045 VCC.n1044 12.2148
R2387 VCC.n1049 VCC.n575 12.2148
R2388 VCC.n1582 VCC.n1162 12.2148
R2389 VCC.n1618 VCC.n1142 12.2148
R2390 VCC.n2154 VCC.n2153 12.2148
R2391 VCC.n2158 VCC.n1684 12.2148
R2392 VCC.n2691 VCC.n2271 12.2148
R2393 VCC.n2727 VCC.n2251 12.2148
R2394 VCC.n3263 VCC.n3262 12.2148
R2395 VCC.n3267 VCC.n2793 12.2148
R2396 VCC.n3800 VCC.n3380 12.2148
R2397 VCC.n3836 VCC.n3360 12.2148
R2398 VCC.n4372 VCC.n4371 12.2148
R2399 VCC.n4376 VCC.n3902 12.2148
R2400 VCC.n4909 VCC.n4489 12.2148
R2401 VCC.n4945 VCC.n4469 12.2148
R2402 VCC.n5481 VCC.n5480 12.2148
R2403 VCC.n5485 VCC.n5011 12.2148
R2404 VCC.n6017 VCC.n5597 12.2148
R2405 VCC.n6053 VCC.n5577 12.2148
R2406 VCC.n6588 VCC.n6587 12.2148
R2407 VCC.n6592 VCC.n6118 12.2148
R2408 VCC.n7124 VCC.n6704 12.2148
R2409 VCC.n7160 VCC.n6684 12.2148
R2410 VCC.n7695 VCC.n7694 12.2148
R2411 VCC.n7699 VCC.n7225 12.2148
R2412 VCC.n8231 VCC.n7811 12.2148
R2413 VCC.n8267 VCC.n7791 12.2148
R2414 VCC.n8615 VCC.n8614 12.2148
R2415 VCC.n8619 VCC.n8332 12.2148
R2416 VCC.n212 VCC.n208 11.4005
R2417 VCC.n334 VCC.n121 11.4005
R2418 VCC.n429 VCC.n81 11.4005
R2419 VCC.n764 VCC.n760 11.4005
R2420 VCC.n886 VCC.n673 11.4005
R2421 VCC.n981 VCC.n633 11.4005
R2422 VCC.n1443 VCC.n1230 11.4005
R2423 VCC.n1539 VCC.n1190 11.4005
R2424 VCC.n1322 VCC.n1318 11.4005
R2425 VCC.n1873 VCC.n1869 11.4005
R2426 VCC.n1995 VCC.n1782 11.4005
R2427 VCC.n2090 VCC.n1742 11.4005
R2428 VCC.n2552 VCC.n2339 11.4005
R2429 VCC.n2648 VCC.n2299 11.4005
R2430 VCC.n2431 VCC.n2427 11.4005
R2431 VCC.n2982 VCC.n2978 11.4005
R2432 VCC.n3104 VCC.n2891 11.4005
R2433 VCC.n3199 VCC.n2851 11.4005
R2434 VCC.n3661 VCC.n3448 11.4005
R2435 VCC.n3757 VCC.n3408 11.4005
R2436 VCC.n3540 VCC.n3536 11.4005
R2437 VCC.n4091 VCC.n4087 11.4005
R2438 VCC.n4213 VCC.n4000 11.4005
R2439 VCC.n4308 VCC.n3960 11.4005
R2440 VCC.n4770 VCC.n4557 11.4005
R2441 VCC.n4866 VCC.n4517 11.4005
R2442 VCC.n4649 VCC.n4645 11.4005
R2443 VCC.n5200 VCC.n5196 11.4005
R2444 VCC.n5322 VCC.n5109 11.4005
R2445 VCC.n5417 VCC.n5069 11.4005
R2446 VCC.n5878 VCC.n5665 11.4005
R2447 VCC.n5974 VCC.n5625 11.4005
R2448 VCC.n5757 VCC.n5753 11.4005
R2449 VCC.n6307 VCC.n6303 11.4005
R2450 VCC.n6429 VCC.n6216 11.4005
R2451 VCC.n6524 VCC.n6176 11.4005
R2452 VCC.n6985 VCC.n6772 11.4005
R2453 VCC.n7081 VCC.n6732 11.4005
R2454 VCC.n6864 VCC.n6860 11.4005
R2455 VCC.n7414 VCC.n7410 11.4005
R2456 VCC.n7536 VCC.n7323 11.4005
R2457 VCC.n7631 VCC.n7283 11.4005
R2458 VCC.n8092 VCC.n7879 11.4005
R2459 VCC.n8188 VCC.n7839 11.4005
R2460 VCC.n7971 VCC.n7967 11.4005
R2461 VCC.n8456 VCC.n8430 11.4005
R2462 VCC.n8551 VCC.n8390 11.4005
R2463 VCC.n474 VCC.n55 10.5862
R2464 VCC.n528 VCC.n21 10.5862
R2465 VCC.n1026 VCC.n607 10.5862
R2466 VCC.n1080 VCC.n573 10.5862
R2467 VCC.n1579 VCC.n1161 10.5862
R2468 VCC.n1650 VCC.n1115 10.5862
R2469 VCC.n2135 VCC.n1716 10.5862
R2470 VCC.n2189 VCC.n1682 10.5862
R2471 VCC.n2688 VCC.n2270 10.5862
R2472 VCC.n2759 VCC.n2224 10.5862
R2473 VCC.n3244 VCC.n2825 10.5862
R2474 VCC.n3298 VCC.n2791 10.5862
R2475 VCC.n3797 VCC.n3379 10.5862
R2476 VCC.n3868 VCC.n3333 10.5862
R2477 VCC.n4353 VCC.n3934 10.5862
R2478 VCC.n4407 VCC.n3900 10.5862
R2479 VCC.n4906 VCC.n4488 10.5862
R2480 VCC.n4977 VCC.n4442 10.5862
R2481 VCC.n5462 VCC.n5043 10.5862
R2482 VCC.n5516 VCC.n5009 10.5862
R2483 VCC.n6014 VCC.n5596 10.5862
R2484 VCC.n6085 VCC.n5550 10.5862
R2485 VCC.n6569 VCC.n6150 10.5862
R2486 VCC.n6623 VCC.n6116 10.5862
R2487 VCC.n7121 VCC.n6703 10.5862
R2488 VCC.n7192 VCC.n6657 10.5862
R2489 VCC.n7676 VCC.n7257 10.5862
R2490 VCC.n7730 VCC.n7223 10.5862
R2491 VCC.n8228 VCC.n7810 10.5862
R2492 VCC.n8299 VCC.n7764 10.5862
R2493 VCC.n8596 VCC.n8364 10.5862
R2494 VCC.n8650 VCC.n8330 10.5862
R2495 VCC.n425 VCC.n420 10.5561
R2496 VCC.n977 VCC.n972 10.5561
R2497 VCC.n1535 VCC.n1528 10.5561
R2498 VCC.n2086 VCC.n2081 10.5561
R2499 VCC.n2644 VCC.n2637 10.5561
R2500 VCC.n3195 VCC.n3190 10.5561
R2501 VCC.n3753 VCC.n3746 10.5561
R2502 VCC.n4304 VCC.n4299 10.5561
R2503 VCC.n4862 VCC.n4855 10.5561
R2504 VCC.n5413 VCC.n5408 10.5561
R2505 VCC.n5970 VCC.n5963 10.5561
R2506 VCC.n6520 VCC.n6515 10.5561
R2507 VCC.n7077 VCC.n7070 10.5561
R2508 VCC.n7627 VCC.n7622 10.5561
R2509 VCC.n8184 VCC.n8177 10.5561
R2510 VCC.n8547 VCC.n8542 10.5561
R2511 VCC.n549 VCC.n548 9.80483
R2512 VCC.n1103 VCC.n1102 9.80483
R2513 VCC.n1657 VCC.n1111 9.80483
R2514 VCC.n2212 VCC.n2211 9.80483
R2515 VCC.n2766 VCC.n2220 9.80483
R2516 VCC.n3321 VCC.n3320 9.80483
R2517 VCC.n3875 VCC.n3329 9.80483
R2518 VCC.n4430 VCC.n4429 9.80483
R2519 VCC.n4984 VCC.n4438 9.80483
R2520 VCC.n5539 VCC.n5538 9.80483
R2521 VCC.n6092 VCC.n5546 9.80483
R2522 VCC.n6646 VCC.n6645 9.80483
R2523 VCC.n7199 VCC.n6653 9.80483
R2524 VCC.n7753 VCC.n7752 9.80483
R2525 VCC.n8306 VCC.n7760 9.80483
R2526 VCC.n8673 VCC.n8672 9.80483
R2527 VCC.n424 VCC.n65 9.38146
R2528 VCC.n976 VCC.n617 9.38146
R2529 VCC.n2085 VCC.n1726 9.38146
R2530 VCC.n3194 VCC.n2835 9.38146
R2531 VCC.n4303 VCC.n3944 9.38146
R2532 VCC.n5412 VCC.n5053 9.38146
R2533 VCC.n6519 VCC.n6160 9.38146
R2534 VCC.n7626 VCC.n7267 9.38146
R2535 VCC.n8546 VCC.n8374 9.38146
R2536 VCC.n1534 VCC.n1174 9.38145
R2537 VCC.n2643 VCC.n2283 9.38145
R2538 VCC.n3752 VCC.n3392 9.38145
R2539 VCC.n4861 VCC.n4501 9.38145
R2540 VCC.n5969 VCC.n5609 9.38145
R2541 VCC.n7076 VCC.n6716 9.38145
R2542 VCC.n8183 VCC.n7823 9.38145
R2543 VCC.n233 VCC.n232 9.3005
R2544 VCC.n202 VCC.n201 9.3005
R2545 VCC.n298 VCC.n297 9.3005
R2546 VCC.n273 VCC.n272 9.3005
R2547 VCC.n161 VCC.n160 9.3005
R2548 VCC.n162 VCC.n156 9.3005
R2549 VCC.n151 VCC.n150 9.3005
R2550 VCC.n152 VCC.n151 9.3005
R2551 VCC.n267 VCC.n152 9.3005
R2552 VCC.n145 VCC.n144 9.3005
R2553 VCC.n287 VCC.n134 9.3005
R2554 VCC.n288 VCC.n287 9.3005
R2555 VCC.n289 VCC.n288 9.3005
R2556 VCC.n139 VCC.n137 9.3005
R2557 VCC.n295 VCC.n294 9.3005
R2558 VCC.n177 VCC.n176 9.3005
R2559 VCC.n214 VCC.n213 9.3005
R2560 VCC.n213 VCC.n212 9.3005
R2561 VCC.n212 VCC.n211 9.3005
R2562 VCC.n196 VCC.n195 9.3005
R2563 VCC.n223 VCC.n222 9.3005
R2564 VCC.n223 VCC.n179 9.3005
R2565 VCC.n227 VCC.n179 9.3005
R2566 VCC.n170 VCC.n169 9.3005
R2567 VCC.n169 VCC.n154 9.3005
R2568 VCC.n154 VCC.n153 9.3005
R2569 VCC.n248 VCC.n168 9.3005
R2570 VCC.n250 VCC.n249 9.3005
R2571 VCC.n357 VCC.n356 9.3005
R2572 VCC.n327 VCC.n326 9.3005
R2573 VCC.n433 VCC.n432 9.3005
R2574 VCC.n400 VCC.n399 9.3005
R2575 VCC.n389 VCC.n95 9.3005
R2576 VCC.n388 VCC.n387 9.3005
R2577 VCC.n85 VCC.n84 9.3005
R2578 VCC.n78 VCC.n76 9.3005
R2579 VCC.n111 VCC.n110 9.3005
R2580 VCC.n325 VCC.n320 9.3005
R2581 VCC.n365 VCC.n105 9.3005
R2582 VCC.n98 VCC.n97 9.3005
R2583 VCC.n392 VCC.n90 9.3005
R2584 VCC.n393 VCC.n392 9.3005
R2585 VCC.n394 VCC.n393 9.3005
R2586 VCC.n413 VCC.n73 9.3005
R2587 VCC.n413 VCC.n83 9.3005
R2588 VCC.n83 VCC.n82 9.3005
R2589 VCC.n430 VCC.n68 9.3005
R2590 VCC.n430 VCC.n429 9.3005
R2591 VCC.n429 VCC.n428 9.3005
R2592 VCC.n333 VCC.n332 9.3005
R2593 VCC.n334 VCC.n333 9.3005
R2594 VCC.n335 VCC.n334 9.3005
R2595 VCC.n342 VCC.n341 9.3005
R2596 VCC.n341 VCC.n109 9.3005
R2597 VCC.n109 VCC.n108 9.3005
R2598 VCC.n364 VCC.n104 9.3005
R2599 VCC.n364 VCC.n363 9.3005
R2600 VCC.n363 VCC.n362 9.3005
R2601 VCC.n477 VCC.n476 9.3005
R2602 VCC.n523 VCC.n522 9.3005
R2603 VCC.n524 VCC.n523 9.3005
R2604 VCC.n525 VCC.n524 9.3005
R2605 VCC.n8 VCC.n7 9.3005
R2606 VCC.n516 VCC.n515 9.3005
R2607 VCC.n544 VCC.n543 9.3005
R2608 VCC.n532 VCC.n531 9.3005
R2609 VCC.n531 VCC.n6 9.3005
R2610 VCC.n6 VCC.n5 9.3005
R2611 VCC.n490 VCC.n489 9.3005
R2612 VCC.n490 VCC.n42 9.3005
R2613 VCC.n472 VCC.n42 9.3005
R2614 VCC.n469 VCC.n468 9.3005
R2615 VCC.n470 VCC.n469 9.3005
R2616 VCC.n425 VCC.n424 9.3005
R2617 VCC.n785 VCC.n784 9.3005
R2618 VCC.n754 VCC.n753 9.3005
R2619 VCC.n850 VCC.n849 9.3005
R2620 VCC.n825 VCC.n824 9.3005
R2621 VCC.n713 VCC.n712 9.3005
R2622 VCC.n714 VCC.n708 9.3005
R2623 VCC.n703 VCC.n702 9.3005
R2624 VCC.n704 VCC.n703 9.3005
R2625 VCC.n819 VCC.n704 9.3005
R2626 VCC.n697 VCC.n696 9.3005
R2627 VCC.n839 VCC.n686 9.3005
R2628 VCC.n840 VCC.n839 9.3005
R2629 VCC.n841 VCC.n840 9.3005
R2630 VCC.n691 VCC.n689 9.3005
R2631 VCC.n847 VCC.n846 9.3005
R2632 VCC.n729 VCC.n728 9.3005
R2633 VCC.n766 VCC.n765 9.3005
R2634 VCC.n765 VCC.n764 9.3005
R2635 VCC.n764 VCC.n763 9.3005
R2636 VCC.n748 VCC.n747 9.3005
R2637 VCC.n775 VCC.n774 9.3005
R2638 VCC.n775 VCC.n731 9.3005
R2639 VCC.n779 VCC.n731 9.3005
R2640 VCC.n722 VCC.n721 9.3005
R2641 VCC.n721 VCC.n706 9.3005
R2642 VCC.n706 VCC.n705 9.3005
R2643 VCC.n800 VCC.n720 9.3005
R2644 VCC.n802 VCC.n801 9.3005
R2645 VCC.n909 VCC.n908 9.3005
R2646 VCC.n879 VCC.n878 9.3005
R2647 VCC.n985 VCC.n984 9.3005
R2648 VCC.n952 VCC.n951 9.3005
R2649 VCC.n941 VCC.n647 9.3005
R2650 VCC.n940 VCC.n939 9.3005
R2651 VCC.n637 VCC.n636 9.3005
R2652 VCC.n630 VCC.n628 9.3005
R2653 VCC.n663 VCC.n662 9.3005
R2654 VCC.n877 VCC.n872 9.3005
R2655 VCC.n917 VCC.n657 9.3005
R2656 VCC.n650 VCC.n649 9.3005
R2657 VCC.n944 VCC.n642 9.3005
R2658 VCC.n945 VCC.n944 9.3005
R2659 VCC.n946 VCC.n945 9.3005
R2660 VCC.n965 VCC.n625 9.3005
R2661 VCC.n965 VCC.n635 9.3005
R2662 VCC.n635 VCC.n634 9.3005
R2663 VCC.n982 VCC.n620 9.3005
R2664 VCC.n982 VCC.n981 9.3005
R2665 VCC.n981 VCC.n980 9.3005
R2666 VCC.n885 VCC.n884 9.3005
R2667 VCC.n886 VCC.n885 9.3005
R2668 VCC.n887 VCC.n886 9.3005
R2669 VCC.n894 VCC.n893 9.3005
R2670 VCC.n893 VCC.n661 9.3005
R2671 VCC.n661 VCC.n660 9.3005
R2672 VCC.n916 VCC.n656 9.3005
R2673 VCC.n916 VCC.n915 9.3005
R2674 VCC.n915 VCC.n914 9.3005
R2675 VCC.n1075 VCC.n1074 9.3005
R2676 VCC.n1076 VCC.n1075 9.3005
R2677 VCC.n1077 VCC.n1076 9.3005
R2678 VCC.n1021 VCC.n1020 9.3005
R2679 VCC.n1022 VCC.n1021 9.3005
R2680 VCC.n1029 VCC.n1028 9.3005
R2681 VCC.n1042 VCC.n1041 9.3005
R2682 VCC.n1042 VCC.n594 9.3005
R2683 VCC.n1024 VCC.n594 9.3005
R2684 VCC.n1068 VCC.n1067 9.3005
R2685 VCC.n1084 VCC.n1083 9.3005
R2686 VCC.n1083 VCC.n560 9.3005
R2687 VCC.n560 VCC.n559 9.3005
R2688 VCC.n562 VCC.n561 9.3005
R2689 VCC.n1098 VCC.n1097 9.3005
R2690 VCC.n977 VCC.n976 9.3005
R2691 VCC.n1140 VCC.n1139 9.3005
R2692 VCC.n1125 VCC.n1124 9.3005
R2693 VCC.n1123 VCC.n1122 9.3005
R2694 VCC.n1595 VCC.n1594 9.3005
R2695 VCC.n1588 VCC.n1587 9.3005
R2696 VCC.n1587 VCC.n1586 9.3005
R2697 VCC.n1586 VCC.n1585 9.3005
R2698 VCC.n1648 VCC.n1647 9.3005
R2699 VCC.n1648 VCC.n1113 9.3005
R2700 VCC.n1652 VCC.n1113 9.3005
R2701 VCC.n1624 VCC.n1623 9.3005
R2702 VCC.n1623 VCC.n1622 9.3005
R2703 VCC.n1622 VCC.n1621 9.3005
R2704 VCC.n1577 VCC.n1164 9.3005
R2705 VCC.n1164 VCC.n1163 9.3005
R2706 VCC.n1535 VCC.n1534 9.3005
R2707 VCC.n1543 VCC.n1542 9.3005
R2708 VCC.n1509 VCC.n1508 9.3005
R2709 VCC.n1498 VCC.n1204 9.3005
R2710 VCC.n1207 VCC.n1206 9.3005
R2711 VCC.n1451 VCC.n1450 9.3005
R2712 VCC.n1450 VCC.n1218 9.3005
R2713 VCC.n1218 VCC.n1217 9.3005
R2714 VCC.n1220 VCC.n1219 9.3005
R2715 VCC.n1466 VCC.n1465 9.3005
R2716 VCC.n1473 VCC.n1213 9.3005
R2717 VCC.n1473 VCC.n1472 9.3005
R2718 VCC.n1472 VCC.n1471 9.3005
R2719 VCC.n1474 VCC.n1214 9.3005
R2720 VCC.n1497 VCC.n1496 9.3005
R2721 VCC.n1501 VCC.n1199 9.3005
R2722 VCC.n1502 VCC.n1501 9.3005
R2723 VCC.n1503 VCC.n1502 9.3005
R2724 VCC.n1194 VCC.n1193 9.3005
R2725 VCC.n1522 VCC.n1182 9.3005
R2726 VCC.n1522 VCC.n1192 9.3005
R2727 VCC.n1192 VCC.n1191 9.3005
R2728 VCC.n1187 VCC.n1185 9.3005
R2729 VCC.n1540 VCC.n1177 9.3005
R2730 VCC.n1540 VCC.n1539 9.3005
R2731 VCC.n1539 VCC.n1538 9.3005
R2732 VCC.n1442 VCC.n1441 9.3005
R2733 VCC.n1443 VCC.n1442 9.3005
R2734 VCC.n1444 VCC.n1443 9.3005
R2735 VCC.n1434 VCC.n1430 9.3005
R2736 VCC.n1436 VCC.n1435 9.3005
R2737 VCC.n1408 VCC.n1407 9.3005
R2738 VCC.n1383 VCC.n1382 9.3005
R2739 VCC.n1271 VCC.n1270 9.3005
R2740 VCC.n1360 VCC.n1359 9.3005
R2741 VCC.n1333 VCC.n1332 9.3005
R2742 VCC.n1333 VCC.n1289 9.3005
R2743 VCC.n1337 VCC.n1289 9.3005
R2744 VCC.n1287 VCC.n1286 9.3005
R2745 VCC.n1343 VCC.n1342 9.3005
R2746 VCC.n1280 VCC.n1279 9.3005
R2747 VCC.n1279 VCC.n1264 9.3005
R2748 VCC.n1264 VCC.n1263 9.3005
R2749 VCC.n1358 VCC.n1278 9.3005
R2750 VCC.n1272 VCC.n1266 9.3005
R2751 VCC.n1261 VCC.n1260 9.3005
R2752 VCC.n1262 VCC.n1261 9.3005
R2753 VCC.n1377 VCC.n1262 9.3005
R2754 VCC.n1255 VCC.n1254 9.3005
R2755 VCC.n1397 VCC.n1244 9.3005
R2756 VCC.n1398 VCC.n1397 9.3005
R2757 VCC.n1399 VCC.n1398 9.3005
R2758 VCC.n1249 VCC.n1247 9.3005
R2759 VCC.n1405 VCC.n1404 9.3005
R2760 VCC.n1324 VCC.n1323 9.3005
R2761 VCC.n1323 VCC.n1322 9.3005
R2762 VCC.n1322 VCC.n1321 9.3005
R2763 VCC.n1306 VCC.n1305 9.3005
R2764 VCC.n1312 VCC.n1311 9.3005
R2765 VCC.n1894 VCC.n1893 9.3005
R2766 VCC.n1863 VCC.n1862 9.3005
R2767 VCC.n1959 VCC.n1958 9.3005
R2768 VCC.n1934 VCC.n1933 9.3005
R2769 VCC.n1822 VCC.n1821 9.3005
R2770 VCC.n1823 VCC.n1817 9.3005
R2771 VCC.n1812 VCC.n1811 9.3005
R2772 VCC.n1813 VCC.n1812 9.3005
R2773 VCC.n1928 VCC.n1813 9.3005
R2774 VCC.n1806 VCC.n1805 9.3005
R2775 VCC.n1948 VCC.n1795 9.3005
R2776 VCC.n1949 VCC.n1948 9.3005
R2777 VCC.n1950 VCC.n1949 9.3005
R2778 VCC.n1800 VCC.n1798 9.3005
R2779 VCC.n1956 VCC.n1955 9.3005
R2780 VCC.n1838 VCC.n1837 9.3005
R2781 VCC.n1875 VCC.n1874 9.3005
R2782 VCC.n1874 VCC.n1873 9.3005
R2783 VCC.n1873 VCC.n1872 9.3005
R2784 VCC.n1857 VCC.n1856 9.3005
R2785 VCC.n1884 VCC.n1883 9.3005
R2786 VCC.n1884 VCC.n1840 9.3005
R2787 VCC.n1888 VCC.n1840 9.3005
R2788 VCC.n1831 VCC.n1830 9.3005
R2789 VCC.n1830 VCC.n1815 9.3005
R2790 VCC.n1815 VCC.n1814 9.3005
R2791 VCC.n1909 VCC.n1829 9.3005
R2792 VCC.n1911 VCC.n1910 9.3005
R2793 VCC.n2018 VCC.n2017 9.3005
R2794 VCC.n1988 VCC.n1987 9.3005
R2795 VCC.n2094 VCC.n2093 9.3005
R2796 VCC.n2061 VCC.n2060 9.3005
R2797 VCC.n2050 VCC.n1756 9.3005
R2798 VCC.n2049 VCC.n2048 9.3005
R2799 VCC.n1746 VCC.n1745 9.3005
R2800 VCC.n1739 VCC.n1737 9.3005
R2801 VCC.n1772 VCC.n1771 9.3005
R2802 VCC.n1986 VCC.n1981 9.3005
R2803 VCC.n2026 VCC.n1766 9.3005
R2804 VCC.n1759 VCC.n1758 9.3005
R2805 VCC.n2053 VCC.n1751 9.3005
R2806 VCC.n2054 VCC.n2053 9.3005
R2807 VCC.n2055 VCC.n2054 9.3005
R2808 VCC.n2074 VCC.n1734 9.3005
R2809 VCC.n2074 VCC.n1744 9.3005
R2810 VCC.n1744 VCC.n1743 9.3005
R2811 VCC.n2091 VCC.n1729 9.3005
R2812 VCC.n2091 VCC.n2090 9.3005
R2813 VCC.n2090 VCC.n2089 9.3005
R2814 VCC.n1994 VCC.n1993 9.3005
R2815 VCC.n1995 VCC.n1994 9.3005
R2816 VCC.n1996 VCC.n1995 9.3005
R2817 VCC.n2003 VCC.n2002 9.3005
R2818 VCC.n2002 VCC.n1770 9.3005
R2819 VCC.n1770 VCC.n1769 9.3005
R2820 VCC.n2025 VCC.n1765 9.3005
R2821 VCC.n2025 VCC.n2024 9.3005
R2822 VCC.n2024 VCC.n2023 9.3005
R2823 VCC.n2184 VCC.n2183 9.3005
R2824 VCC.n2185 VCC.n2184 9.3005
R2825 VCC.n2186 VCC.n2185 9.3005
R2826 VCC.n2130 VCC.n2129 9.3005
R2827 VCC.n2131 VCC.n2130 9.3005
R2828 VCC.n2138 VCC.n2137 9.3005
R2829 VCC.n2151 VCC.n2150 9.3005
R2830 VCC.n2151 VCC.n1703 9.3005
R2831 VCC.n2133 VCC.n1703 9.3005
R2832 VCC.n2177 VCC.n2176 9.3005
R2833 VCC.n2193 VCC.n2192 9.3005
R2834 VCC.n2192 VCC.n1669 9.3005
R2835 VCC.n1669 VCC.n1668 9.3005
R2836 VCC.n1671 VCC.n1670 9.3005
R2837 VCC.n2207 VCC.n2206 9.3005
R2838 VCC.n2086 VCC.n2085 9.3005
R2839 VCC.n2249 VCC.n2248 9.3005
R2840 VCC.n2234 VCC.n2233 9.3005
R2841 VCC.n2232 VCC.n2231 9.3005
R2842 VCC.n2704 VCC.n2703 9.3005
R2843 VCC.n2697 VCC.n2696 9.3005
R2844 VCC.n2696 VCC.n2695 9.3005
R2845 VCC.n2695 VCC.n2694 9.3005
R2846 VCC.n2757 VCC.n2756 9.3005
R2847 VCC.n2757 VCC.n2222 9.3005
R2848 VCC.n2761 VCC.n2222 9.3005
R2849 VCC.n2733 VCC.n2732 9.3005
R2850 VCC.n2732 VCC.n2731 9.3005
R2851 VCC.n2731 VCC.n2730 9.3005
R2852 VCC.n2686 VCC.n2273 9.3005
R2853 VCC.n2273 VCC.n2272 9.3005
R2854 VCC.n2644 VCC.n2643 9.3005
R2855 VCC.n2652 VCC.n2651 9.3005
R2856 VCC.n2618 VCC.n2617 9.3005
R2857 VCC.n2607 VCC.n2313 9.3005
R2858 VCC.n2316 VCC.n2315 9.3005
R2859 VCC.n2560 VCC.n2559 9.3005
R2860 VCC.n2559 VCC.n2327 9.3005
R2861 VCC.n2327 VCC.n2326 9.3005
R2862 VCC.n2329 VCC.n2328 9.3005
R2863 VCC.n2575 VCC.n2574 9.3005
R2864 VCC.n2582 VCC.n2322 9.3005
R2865 VCC.n2582 VCC.n2581 9.3005
R2866 VCC.n2581 VCC.n2580 9.3005
R2867 VCC.n2583 VCC.n2323 9.3005
R2868 VCC.n2606 VCC.n2605 9.3005
R2869 VCC.n2610 VCC.n2308 9.3005
R2870 VCC.n2611 VCC.n2610 9.3005
R2871 VCC.n2612 VCC.n2611 9.3005
R2872 VCC.n2303 VCC.n2302 9.3005
R2873 VCC.n2631 VCC.n2291 9.3005
R2874 VCC.n2631 VCC.n2301 9.3005
R2875 VCC.n2301 VCC.n2300 9.3005
R2876 VCC.n2296 VCC.n2294 9.3005
R2877 VCC.n2649 VCC.n2286 9.3005
R2878 VCC.n2649 VCC.n2648 9.3005
R2879 VCC.n2648 VCC.n2647 9.3005
R2880 VCC.n2551 VCC.n2550 9.3005
R2881 VCC.n2552 VCC.n2551 9.3005
R2882 VCC.n2553 VCC.n2552 9.3005
R2883 VCC.n2543 VCC.n2539 9.3005
R2884 VCC.n2545 VCC.n2544 9.3005
R2885 VCC.n2517 VCC.n2516 9.3005
R2886 VCC.n2492 VCC.n2491 9.3005
R2887 VCC.n2380 VCC.n2379 9.3005
R2888 VCC.n2469 VCC.n2468 9.3005
R2889 VCC.n2442 VCC.n2441 9.3005
R2890 VCC.n2442 VCC.n2398 9.3005
R2891 VCC.n2446 VCC.n2398 9.3005
R2892 VCC.n2396 VCC.n2395 9.3005
R2893 VCC.n2452 VCC.n2451 9.3005
R2894 VCC.n2389 VCC.n2388 9.3005
R2895 VCC.n2388 VCC.n2373 9.3005
R2896 VCC.n2373 VCC.n2372 9.3005
R2897 VCC.n2467 VCC.n2387 9.3005
R2898 VCC.n2381 VCC.n2375 9.3005
R2899 VCC.n2370 VCC.n2369 9.3005
R2900 VCC.n2371 VCC.n2370 9.3005
R2901 VCC.n2486 VCC.n2371 9.3005
R2902 VCC.n2364 VCC.n2363 9.3005
R2903 VCC.n2506 VCC.n2353 9.3005
R2904 VCC.n2507 VCC.n2506 9.3005
R2905 VCC.n2508 VCC.n2507 9.3005
R2906 VCC.n2358 VCC.n2356 9.3005
R2907 VCC.n2514 VCC.n2513 9.3005
R2908 VCC.n2433 VCC.n2432 9.3005
R2909 VCC.n2432 VCC.n2431 9.3005
R2910 VCC.n2431 VCC.n2430 9.3005
R2911 VCC.n2415 VCC.n2414 9.3005
R2912 VCC.n2421 VCC.n2420 9.3005
R2913 VCC.n3003 VCC.n3002 9.3005
R2914 VCC.n2972 VCC.n2971 9.3005
R2915 VCC.n3068 VCC.n3067 9.3005
R2916 VCC.n3043 VCC.n3042 9.3005
R2917 VCC.n2931 VCC.n2930 9.3005
R2918 VCC.n2932 VCC.n2926 9.3005
R2919 VCC.n2921 VCC.n2920 9.3005
R2920 VCC.n2922 VCC.n2921 9.3005
R2921 VCC.n3037 VCC.n2922 9.3005
R2922 VCC.n2915 VCC.n2914 9.3005
R2923 VCC.n3057 VCC.n2904 9.3005
R2924 VCC.n3058 VCC.n3057 9.3005
R2925 VCC.n3059 VCC.n3058 9.3005
R2926 VCC.n2909 VCC.n2907 9.3005
R2927 VCC.n3065 VCC.n3064 9.3005
R2928 VCC.n2947 VCC.n2946 9.3005
R2929 VCC.n2984 VCC.n2983 9.3005
R2930 VCC.n2983 VCC.n2982 9.3005
R2931 VCC.n2982 VCC.n2981 9.3005
R2932 VCC.n2966 VCC.n2965 9.3005
R2933 VCC.n2993 VCC.n2992 9.3005
R2934 VCC.n2993 VCC.n2949 9.3005
R2935 VCC.n2997 VCC.n2949 9.3005
R2936 VCC.n2940 VCC.n2939 9.3005
R2937 VCC.n2939 VCC.n2924 9.3005
R2938 VCC.n2924 VCC.n2923 9.3005
R2939 VCC.n3018 VCC.n2938 9.3005
R2940 VCC.n3020 VCC.n3019 9.3005
R2941 VCC.n3127 VCC.n3126 9.3005
R2942 VCC.n3097 VCC.n3096 9.3005
R2943 VCC.n3203 VCC.n3202 9.3005
R2944 VCC.n3170 VCC.n3169 9.3005
R2945 VCC.n3159 VCC.n2865 9.3005
R2946 VCC.n3158 VCC.n3157 9.3005
R2947 VCC.n2855 VCC.n2854 9.3005
R2948 VCC.n2848 VCC.n2846 9.3005
R2949 VCC.n2881 VCC.n2880 9.3005
R2950 VCC.n3095 VCC.n3090 9.3005
R2951 VCC.n3135 VCC.n2875 9.3005
R2952 VCC.n2868 VCC.n2867 9.3005
R2953 VCC.n3162 VCC.n2860 9.3005
R2954 VCC.n3163 VCC.n3162 9.3005
R2955 VCC.n3164 VCC.n3163 9.3005
R2956 VCC.n3183 VCC.n2843 9.3005
R2957 VCC.n3183 VCC.n2853 9.3005
R2958 VCC.n2853 VCC.n2852 9.3005
R2959 VCC.n3200 VCC.n2838 9.3005
R2960 VCC.n3200 VCC.n3199 9.3005
R2961 VCC.n3199 VCC.n3198 9.3005
R2962 VCC.n3103 VCC.n3102 9.3005
R2963 VCC.n3104 VCC.n3103 9.3005
R2964 VCC.n3105 VCC.n3104 9.3005
R2965 VCC.n3112 VCC.n3111 9.3005
R2966 VCC.n3111 VCC.n2879 9.3005
R2967 VCC.n2879 VCC.n2878 9.3005
R2968 VCC.n3134 VCC.n2874 9.3005
R2969 VCC.n3134 VCC.n3133 9.3005
R2970 VCC.n3133 VCC.n3132 9.3005
R2971 VCC.n3293 VCC.n3292 9.3005
R2972 VCC.n3294 VCC.n3293 9.3005
R2973 VCC.n3295 VCC.n3294 9.3005
R2974 VCC.n3239 VCC.n3238 9.3005
R2975 VCC.n3240 VCC.n3239 9.3005
R2976 VCC.n3247 VCC.n3246 9.3005
R2977 VCC.n3260 VCC.n3259 9.3005
R2978 VCC.n3260 VCC.n2812 9.3005
R2979 VCC.n3242 VCC.n2812 9.3005
R2980 VCC.n3286 VCC.n3285 9.3005
R2981 VCC.n3302 VCC.n3301 9.3005
R2982 VCC.n3301 VCC.n2778 9.3005
R2983 VCC.n2778 VCC.n2777 9.3005
R2984 VCC.n2780 VCC.n2779 9.3005
R2985 VCC.n3316 VCC.n3315 9.3005
R2986 VCC.n3195 VCC.n3194 9.3005
R2987 VCC.n3358 VCC.n3357 9.3005
R2988 VCC.n3343 VCC.n3342 9.3005
R2989 VCC.n3341 VCC.n3340 9.3005
R2990 VCC.n3813 VCC.n3812 9.3005
R2991 VCC.n3806 VCC.n3805 9.3005
R2992 VCC.n3805 VCC.n3804 9.3005
R2993 VCC.n3804 VCC.n3803 9.3005
R2994 VCC.n3866 VCC.n3865 9.3005
R2995 VCC.n3866 VCC.n3331 9.3005
R2996 VCC.n3870 VCC.n3331 9.3005
R2997 VCC.n3842 VCC.n3841 9.3005
R2998 VCC.n3841 VCC.n3840 9.3005
R2999 VCC.n3840 VCC.n3839 9.3005
R3000 VCC.n3795 VCC.n3382 9.3005
R3001 VCC.n3382 VCC.n3381 9.3005
R3002 VCC.n3753 VCC.n3752 9.3005
R3003 VCC.n3761 VCC.n3760 9.3005
R3004 VCC.n3727 VCC.n3726 9.3005
R3005 VCC.n3716 VCC.n3422 9.3005
R3006 VCC.n3425 VCC.n3424 9.3005
R3007 VCC.n3669 VCC.n3668 9.3005
R3008 VCC.n3668 VCC.n3436 9.3005
R3009 VCC.n3436 VCC.n3435 9.3005
R3010 VCC.n3438 VCC.n3437 9.3005
R3011 VCC.n3684 VCC.n3683 9.3005
R3012 VCC.n3691 VCC.n3431 9.3005
R3013 VCC.n3691 VCC.n3690 9.3005
R3014 VCC.n3690 VCC.n3689 9.3005
R3015 VCC.n3692 VCC.n3432 9.3005
R3016 VCC.n3715 VCC.n3714 9.3005
R3017 VCC.n3719 VCC.n3417 9.3005
R3018 VCC.n3720 VCC.n3719 9.3005
R3019 VCC.n3721 VCC.n3720 9.3005
R3020 VCC.n3412 VCC.n3411 9.3005
R3021 VCC.n3740 VCC.n3400 9.3005
R3022 VCC.n3740 VCC.n3410 9.3005
R3023 VCC.n3410 VCC.n3409 9.3005
R3024 VCC.n3405 VCC.n3403 9.3005
R3025 VCC.n3758 VCC.n3395 9.3005
R3026 VCC.n3758 VCC.n3757 9.3005
R3027 VCC.n3757 VCC.n3756 9.3005
R3028 VCC.n3660 VCC.n3659 9.3005
R3029 VCC.n3661 VCC.n3660 9.3005
R3030 VCC.n3662 VCC.n3661 9.3005
R3031 VCC.n3652 VCC.n3648 9.3005
R3032 VCC.n3654 VCC.n3653 9.3005
R3033 VCC.n3626 VCC.n3625 9.3005
R3034 VCC.n3601 VCC.n3600 9.3005
R3035 VCC.n3489 VCC.n3488 9.3005
R3036 VCC.n3578 VCC.n3577 9.3005
R3037 VCC.n3551 VCC.n3550 9.3005
R3038 VCC.n3551 VCC.n3507 9.3005
R3039 VCC.n3555 VCC.n3507 9.3005
R3040 VCC.n3505 VCC.n3504 9.3005
R3041 VCC.n3561 VCC.n3560 9.3005
R3042 VCC.n3498 VCC.n3497 9.3005
R3043 VCC.n3497 VCC.n3482 9.3005
R3044 VCC.n3482 VCC.n3481 9.3005
R3045 VCC.n3576 VCC.n3496 9.3005
R3046 VCC.n3490 VCC.n3484 9.3005
R3047 VCC.n3479 VCC.n3478 9.3005
R3048 VCC.n3480 VCC.n3479 9.3005
R3049 VCC.n3595 VCC.n3480 9.3005
R3050 VCC.n3473 VCC.n3472 9.3005
R3051 VCC.n3615 VCC.n3462 9.3005
R3052 VCC.n3616 VCC.n3615 9.3005
R3053 VCC.n3617 VCC.n3616 9.3005
R3054 VCC.n3467 VCC.n3465 9.3005
R3055 VCC.n3623 VCC.n3622 9.3005
R3056 VCC.n3542 VCC.n3541 9.3005
R3057 VCC.n3541 VCC.n3540 9.3005
R3058 VCC.n3540 VCC.n3539 9.3005
R3059 VCC.n3524 VCC.n3523 9.3005
R3060 VCC.n3530 VCC.n3529 9.3005
R3061 VCC.n4112 VCC.n4111 9.3005
R3062 VCC.n4081 VCC.n4080 9.3005
R3063 VCC.n4177 VCC.n4176 9.3005
R3064 VCC.n4152 VCC.n4151 9.3005
R3065 VCC.n4040 VCC.n4039 9.3005
R3066 VCC.n4041 VCC.n4035 9.3005
R3067 VCC.n4030 VCC.n4029 9.3005
R3068 VCC.n4031 VCC.n4030 9.3005
R3069 VCC.n4146 VCC.n4031 9.3005
R3070 VCC.n4024 VCC.n4023 9.3005
R3071 VCC.n4166 VCC.n4013 9.3005
R3072 VCC.n4167 VCC.n4166 9.3005
R3073 VCC.n4168 VCC.n4167 9.3005
R3074 VCC.n4018 VCC.n4016 9.3005
R3075 VCC.n4174 VCC.n4173 9.3005
R3076 VCC.n4056 VCC.n4055 9.3005
R3077 VCC.n4093 VCC.n4092 9.3005
R3078 VCC.n4092 VCC.n4091 9.3005
R3079 VCC.n4091 VCC.n4090 9.3005
R3080 VCC.n4075 VCC.n4074 9.3005
R3081 VCC.n4102 VCC.n4101 9.3005
R3082 VCC.n4102 VCC.n4058 9.3005
R3083 VCC.n4106 VCC.n4058 9.3005
R3084 VCC.n4049 VCC.n4048 9.3005
R3085 VCC.n4048 VCC.n4033 9.3005
R3086 VCC.n4033 VCC.n4032 9.3005
R3087 VCC.n4127 VCC.n4047 9.3005
R3088 VCC.n4129 VCC.n4128 9.3005
R3089 VCC.n4236 VCC.n4235 9.3005
R3090 VCC.n4206 VCC.n4205 9.3005
R3091 VCC.n4312 VCC.n4311 9.3005
R3092 VCC.n4279 VCC.n4278 9.3005
R3093 VCC.n4268 VCC.n3974 9.3005
R3094 VCC.n4267 VCC.n4266 9.3005
R3095 VCC.n3964 VCC.n3963 9.3005
R3096 VCC.n3957 VCC.n3955 9.3005
R3097 VCC.n3990 VCC.n3989 9.3005
R3098 VCC.n4204 VCC.n4199 9.3005
R3099 VCC.n4244 VCC.n3984 9.3005
R3100 VCC.n3977 VCC.n3976 9.3005
R3101 VCC.n4271 VCC.n3969 9.3005
R3102 VCC.n4272 VCC.n4271 9.3005
R3103 VCC.n4273 VCC.n4272 9.3005
R3104 VCC.n4292 VCC.n3952 9.3005
R3105 VCC.n4292 VCC.n3962 9.3005
R3106 VCC.n3962 VCC.n3961 9.3005
R3107 VCC.n4309 VCC.n3947 9.3005
R3108 VCC.n4309 VCC.n4308 9.3005
R3109 VCC.n4308 VCC.n4307 9.3005
R3110 VCC.n4212 VCC.n4211 9.3005
R3111 VCC.n4213 VCC.n4212 9.3005
R3112 VCC.n4214 VCC.n4213 9.3005
R3113 VCC.n4221 VCC.n4220 9.3005
R3114 VCC.n4220 VCC.n3988 9.3005
R3115 VCC.n3988 VCC.n3987 9.3005
R3116 VCC.n4243 VCC.n3983 9.3005
R3117 VCC.n4243 VCC.n4242 9.3005
R3118 VCC.n4242 VCC.n4241 9.3005
R3119 VCC.n4402 VCC.n4401 9.3005
R3120 VCC.n4403 VCC.n4402 9.3005
R3121 VCC.n4404 VCC.n4403 9.3005
R3122 VCC.n4348 VCC.n4347 9.3005
R3123 VCC.n4349 VCC.n4348 9.3005
R3124 VCC.n4356 VCC.n4355 9.3005
R3125 VCC.n4369 VCC.n4368 9.3005
R3126 VCC.n4369 VCC.n3921 9.3005
R3127 VCC.n4351 VCC.n3921 9.3005
R3128 VCC.n4395 VCC.n4394 9.3005
R3129 VCC.n4411 VCC.n4410 9.3005
R3130 VCC.n4410 VCC.n3887 9.3005
R3131 VCC.n3887 VCC.n3886 9.3005
R3132 VCC.n3889 VCC.n3888 9.3005
R3133 VCC.n4425 VCC.n4424 9.3005
R3134 VCC.n4304 VCC.n4303 9.3005
R3135 VCC.n4467 VCC.n4466 9.3005
R3136 VCC.n4452 VCC.n4451 9.3005
R3137 VCC.n4450 VCC.n4449 9.3005
R3138 VCC.n4922 VCC.n4921 9.3005
R3139 VCC.n4915 VCC.n4914 9.3005
R3140 VCC.n4914 VCC.n4913 9.3005
R3141 VCC.n4913 VCC.n4912 9.3005
R3142 VCC.n4975 VCC.n4974 9.3005
R3143 VCC.n4975 VCC.n4440 9.3005
R3144 VCC.n4979 VCC.n4440 9.3005
R3145 VCC.n4951 VCC.n4950 9.3005
R3146 VCC.n4950 VCC.n4949 9.3005
R3147 VCC.n4949 VCC.n4948 9.3005
R3148 VCC.n4904 VCC.n4491 9.3005
R3149 VCC.n4491 VCC.n4490 9.3005
R3150 VCC.n4862 VCC.n4861 9.3005
R3151 VCC.n4870 VCC.n4869 9.3005
R3152 VCC.n4836 VCC.n4835 9.3005
R3153 VCC.n4825 VCC.n4531 9.3005
R3154 VCC.n4534 VCC.n4533 9.3005
R3155 VCC.n4778 VCC.n4777 9.3005
R3156 VCC.n4777 VCC.n4545 9.3005
R3157 VCC.n4545 VCC.n4544 9.3005
R3158 VCC.n4547 VCC.n4546 9.3005
R3159 VCC.n4793 VCC.n4792 9.3005
R3160 VCC.n4800 VCC.n4540 9.3005
R3161 VCC.n4800 VCC.n4799 9.3005
R3162 VCC.n4799 VCC.n4798 9.3005
R3163 VCC.n4801 VCC.n4541 9.3005
R3164 VCC.n4824 VCC.n4823 9.3005
R3165 VCC.n4828 VCC.n4526 9.3005
R3166 VCC.n4829 VCC.n4828 9.3005
R3167 VCC.n4830 VCC.n4829 9.3005
R3168 VCC.n4521 VCC.n4520 9.3005
R3169 VCC.n4849 VCC.n4509 9.3005
R3170 VCC.n4849 VCC.n4519 9.3005
R3171 VCC.n4519 VCC.n4518 9.3005
R3172 VCC.n4514 VCC.n4512 9.3005
R3173 VCC.n4867 VCC.n4504 9.3005
R3174 VCC.n4867 VCC.n4866 9.3005
R3175 VCC.n4866 VCC.n4865 9.3005
R3176 VCC.n4769 VCC.n4768 9.3005
R3177 VCC.n4770 VCC.n4769 9.3005
R3178 VCC.n4771 VCC.n4770 9.3005
R3179 VCC.n4761 VCC.n4757 9.3005
R3180 VCC.n4763 VCC.n4762 9.3005
R3181 VCC.n4735 VCC.n4734 9.3005
R3182 VCC.n4710 VCC.n4709 9.3005
R3183 VCC.n4598 VCC.n4597 9.3005
R3184 VCC.n4687 VCC.n4686 9.3005
R3185 VCC.n4660 VCC.n4659 9.3005
R3186 VCC.n4660 VCC.n4616 9.3005
R3187 VCC.n4664 VCC.n4616 9.3005
R3188 VCC.n4614 VCC.n4613 9.3005
R3189 VCC.n4670 VCC.n4669 9.3005
R3190 VCC.n4607 VCC.n4606 9.3005
R3191 VCC.n4606 VCC.n4591 9.3005
R3192 VCC.n4591 VCC.n4590 9.3005
R3193 VCC.n4685 VCC.n4605 9.3005
R3194 VCC.n4599 VCC.n4593 9.3005
R3195 VCC.n4588 VCC.n4587 9.3005
R3196 VCC.n4589 VCC.n4588 9.3005
R3197 VCC.n4704 VCC.n4589 9.3005
R3198 VCC.n4582 VCC.n4581 9.3005
R3199 VCC.n4724 VCC.n4571 9.3005
R3200 VCC.n4725 VCC.n4724 9.3005
R3201 VCC.n4726 VCC.n4725 9.3005
R3202 VCC.n4576 VCC.n4574 9.3005
R3203 VCC.n4732 VCC.n4731 9.3005
R3204 VCC.n4651 VCC.n4650 9.3005
R3205 VCC.n4650 VCC.n4649 9.3005
R3206 VCC.n4649 VCC.n4648 9.3005
R3207 VCC.n4633 VCC.n4632 9.3005
R3208 VCC.n4639 VCC.n4638 9.3005
R3209 VCC.n5221 VCC.n5220 9.3005
R3210 VCC.n5190 VCC.n5189 9.3005
R3211 VCC.n5286 VCC.n5285 9.3005
R3212 VCC.n5261 VCC.n5260 9.3005
R3213 VCC.n5149 VCC.n5148 9.3005
R3214 VCC.n5150 VCC.n5144 9.3005
R3215 VCC.n5139 VCC.n5138 9.3005
R3216 VCC.n5140 VCC.n5139 9.3005
R3217 VCC.n5255 VCC.n5140 9.3005
R3218 VCC.n5133 VCC.n5132 9.3005
R3219 VCC.n5275 VCC.n5122 9.3005
R3220 VCC.n5276 VCC.n5275 9.3005
R3221 VCC.n5277 VCC.n5276 9.3005
R3222 VCC.n5127 VCC.n5125 9.3005
R3223 VCC.n5283 VCC.n5282 9.3005
R3224 VCC.n5165 VCC.n5164 9.3005
R3225 VCC.n5202 VCC.n5201 9.3005
R3226 VCC.n5201 VCC.n5200 9.3005
R3227 VCC.n5200 VCC.n5199 9.3005
R3228 VCC.n5184 VCC.n5183 9.3005
R3229 VCC.n5211 VCC.n5210 9.3005
R3230 VCC.n5211 VCC.n5167 9.3005
R3231 VCC.n5215 VCC.n5167 9.3005
R3232 VCC.n5158 VCC.n5157 9.3005
R3233 VCC.n5157 VCC.n5142 9.3005
R3234 VCC.n5142 VCC.n5141 9.3005
R3235 VCC.n5236 VCC.n5156 9.3005
R3236 VCC.n5238 VCC.n5237 9.3005
R3237 VCC.n5345 VCC.n5344 9.3005
R3238 VCC.n5315 VCC.n5314 9.3005
R3239 VCC.n5421 VCC.n5420 9.3005
R3240 VCC.n5388 VCC.n5387 9.3005
R3241 VCC.n5377 VCC.n5083 9.3005
R3242 VCC.n5376 VCC.n5375 9.3005
R3243 VCC.n5073 VCC.n5072 9.3005
R3244 VCC.n5066 VCC.n5064 9.3005
R3245 VCC.n5099 VCC.n5098 9.3005
R3246 VCC.n5313 VCC.n5308 9.3005
R3247 VCC.n5353 VCC.n5093 9.3005
R3248 VCC.n5086 VCC.n5085 9.3005
R3249 VCC.n5380 VCC.n5078 9.3005
R3250 VCC.n5381 VCC.n5380 9.3005
R3251 VCC.n5382 VCC.n5381 9.3005
R3252 VCC.n5401 VCC.n5061 9.3005
R3253 VCC.n5401 VCC.n5071 9.3005
R3254 VCC.n5071 VCC.n5070 9.3005
R3255 VCC.n5418 VCC.n5056 9.3005
R3256 VCC.n5418 VCC.n5417 9.3005
R3257 VCC.n5417 VCC.n5416 9.3005
R3258 VCC.n5321 VCC.n5320 9.3005
R3259 VCC.n5322 VCC.n5321 9.3005
R3260 VCC.n5323 VCC.n5322 9.3005
R3261 VCC.n5330 VCC.n5329 9.3005
R3262 VCC.n5329 VCC.n5097 9.3005
R3263 VCC.n5097 VCC.n5096 9.3005
R3264 VCC.n5352 VCC.n5092 9.3005
R3265 VCC.n5352 VCC.n5351 9.3005
R3266 VCC.n5351 VCC.n5350 9.3005
R3267 VCC.n5511 VCC.n5510 9.3005
R3268 VCC.n5512 VCC.n5511 9.3005
R3269 VCC.n5513 VCC.n5512 9.3005
R3270 VCC.n5457 VCC.n5456 9.3005
R3271 VCC.n5458 VCC.n5457 9.3005
R3272 VCC.n5465 VCC.n5464 9.3005
R3273 VCC.n5478 VCC.n5477 9.3005
R3274 VCC.n5478 VCC.n5030 9.3005
R3275 VCC.n5460 VCC.n5030 9.3005
R3276 VCC.n5504 VCC.n5503 9.3005
R3277 VCC.n5520 VCC.n5519 9.3005
R3278 VCC.n5519 VCC.n4996 9.3005
R3279 VCC.n4996 VCC.n4995 9.3005
R3280 VCC.n4998 VCC.n4997 9.3005
R3281 VCC.n5534 VCC.n5533 9.3005
R3282 VCC.n5413 VCC.n5412 9.3005
R3283 VCC.n5575 VCC.n5574 9.3005
R3284 VCC.n5560 VCC.n5559 9.3005
R3285 VCC.n5558 VCC.n5557 9.3005
R3286 VCC.n6030 VCC.n6029 9.3005
R3287 VCC.n6023 VCC.n6022 9.3005
R3288 VCC.n6022 VCC.n6021 9.3005
R3289 VCC.n6021 VCC.n6020 9.3005
R3290 VCC.n6083 VCC.n6082 9.3005
R3291 VCC.n6083 VCC.n5548 9.3005
R3292 VCC.n6087 VCC.n5548 9.3005
R3293 VCC.n6059 VCC.n6058 9.3005
R3294 VCC.n6058 VCC.n6057 9.3005
R3295 VCC.n6057 VCC.n6056 9.3005
R3296 VCC.n6012 VCC.n5599 9.3005
R3297 VCC.n5599 VCC.n5598 9.3005
R3298 VCC.n5970 VCC.n5969 9.3005
R3299 VCC.n5978 VCC.n5977 9.3005
R3300 VCC.n5944 VCC.n5943 9.3005
R3301 VCC.n5933 VCC.n5639 9.3005
R3302 VCC.n5642 VCC.n5641 9.3005
R3303 VCC.n5886 VCC.n5885 9.3005
R3304 VCC.n5885 VCC.n5653 9.3005
R3305 VCC.n5653 VCC.n5652 9.3005
R3306 VCC.n5655 VCC.n5654 9.3005
R3307 VCC.n5901 VCC.n5900 9.3005
R3308 VCC.n5908 VCC.n5648 9.3005
R3309 VCC.n5908 VCC.n5907 9.3005
R3310 VCC.n5907 VCC.n5906 9.3005
R3311 VCC.n5909 VCC.n5649 9.3005
R3312 VCC.n5932 VCC.n5931 9.3005
R3313 VCC.n5936 VCC.n5634 9.3005
R3314 VCC.n5937 VCC.n5936 9.3005
R3315 VCC.n5938 VCC.n5937 9.3005
R3316 VCC.n5629 VCC.n5628 9.3005
R3317 VCC.n5957 VCC.n5617 9.3005
R3318 VCC.n5957 VCC.n5627 9.3005
R3319 VCC.n5627 VCC.n5626 9.3005
R3320 VCC.n5622 VCC.n5620 9.3005
R3321 VCC.n5975 VCC.n5612 9.3005
R3322 VCC.n5975 VCC.n5974 9.3005
R3323 VCC.n5974 VCC.n5973 9.3005
R3324 VCC.n5877 VCC.n5876 9.3005
R3325 VCC.n5878 VCC.n5877 9.3005
R3326 VCC.n5879 VCC.n5878 9.3005
R3327 VCC.n5869 VCC.n5865 9.3005
R3328 VCC.n5871 VCC.n5870 9.3005
R3329 VCC.n5843 VCC.n5842 9.3005
R3330 VCC.n5818 VCC.n5817 9.3005
R3331 VCC.n5706 VCC.n5705 9.3005
R3332 VCC.n5795 VCC.n5794 9.3005
R3333 VCC.n5768 VCC.n5767 9.3005
R3334 VCC.n5768 VCC.n5724 9.3005
R3335 VCC.n5772 VCC.n5724 9.3005
R3336 VCC.n5722 VCC.n5721 9.3005
R3337 VCC.n5778 VCC.n5777 9.3005
R3338 VCC.n5715 VCC.n5714 9.3005
R3339 VCC.n5714 VCC.n5699 9.3005
R3340 VCC.n5699 VCC.n5698 9.3005
R3341 VCC.n5793 VCC.n5713 9.3005
R3342 VCC.n5707 VCC.n5701 9.3005
R3343 VCC.n5696 VCC.n5695 9.3005
R3344 VCC.n5697 VCC.n5696 9.3005
R3345 VCC.n5812 VCC.n5697 9.3005
R3346 VCC.n5690 VCC.n5689 9.3005
R3347 VCC.n5832 VCC.n5679 9.3005
R3348 VCC.n5833 VCC.n5832 9.3005
R3349 VCC.n5834 VCC.n5833 9.3005
R3350 VCC.n5684 VCC.n5682 9.3005
R3351 VCC.n5840 VCC.n5839 9.3005
R3352 VCC.n5759 VCC.n5758 9.3005
R3353 VCC.n5758 VCC.n5757 9.3005
R3354 VCC.n5757 VCC.n5756 9.3005
R3355 VCC.n5741 VCC.n5740 9.3005
R3356 VCC.n5747 VCC.n5746 9.3005
R3357 VCC.n6328 VCC.n6327 9.3005
R3358 VCC.n6297 VCC.n6296 9.3005
R3359 VCC.n6393 VCC.n6392 9.3005
R3360 VCC.n6368 VCC.n6367 9.3005
R3361 VCC.n6256 VCC.n6255 9.3005
R3362 VCC.n6257 VCC.n6251 9.3005
R3363 VCC.n6246 VCC.n6245 9.3005
R3364 VCC.n6247 VCC.n6246 9.3005
R3365 VCC.n6362 VCC.n6247 9.3005
R3366 VCC.n6240 VCC.n6239 9.3005
R3367 VCC.n6382 VCC.n6229 9.3005
R3368 VCC.n6383 VCC.n6382 9.3005
R3369 VCC.n6384 VCC.n6383 9.3005
R3370 VCC.n6234 VCC.n6232 9.3005
R3371 VCC.n6390 VCC.n6389 9.3005
R3372 VCC.n6272 VCC.n6271 9.3005
R3373 VCC.n6309 VCC.n6308 9.3005
R3374 VCC.n6308 VCC.n6307 9.3005
R3375 VCC.n6307 VCC.n6306 9.3005
R3376 VCC.n6291 VCC.n6290 9.3005
R3377 VCC.n6318 VCC.n6317 9.3005
R3378 VCC.n6318 VCC.n6274 9.3005
R3379 VCC.n6322 VCC.n6274 9.3005
R3380 VCC.n6265 VCC.n6264 9.3005
R3381 VCC.n6264 VCC.n6249 9.3005
R3382 VCC.n6249 VCC.n6248 9.3005
R3383 VCC.n6343 VCC.n6263 9.3005
R3384 VCC.n6345 VCC.n6344 9.3005
R3385 VCC.n6452 VCC.n6451 9.3005
R3386 VCC.n6422 VCC.n6421 9.3005
R3387 VCC.n6528 VCC.n6527 9.3005
R3388 VCC.n6495 VCC.n6494 9.3005
R3389 VCC.n6484 VCC.n6190 9.3005
R3390 VCC.n6483 VCC.n6482 9.3005
R3391 VCC.n6180 VCC.n6179 9.3005
R3392 VCC.n6173 VCC.n6171 9.3005
R3393 VCC.n6206 VCC.n6205 9.3005
R3394 VCC.n6420 VCC.n6415 9.3005
R3395 VCC.n6460 VCC.n6200 9.3005
R3396 VCC.n6193 VCC.n6192 9.3005
R3397 VCC.n6487 VCC.n6185 9.3005
R3398 VCC.n6488 VCC.n6487 9.3005
R3399 VCC.n6489 VCC.n6488 9.3005
R3400 VCC.n6508 VCC.n6168 9.3005
R3401 VCC.n6508 VCC.n6178 9.3005
R3402 VCC.n6178 VCC.n6177 9.3005
R3403 VCC.n6525 VCC.n6163 9.3005
R3404 VCC.n6525 VCC.n6524 9.3005
R3405 VCC.n6524 VCC.n6523 9.3005
R3406 VCC.n6428 VCC.n6427 9.3005
R3407 VCC.n6429 VCC.n6428 9.3005
R3408 VCC.n6430 VCC.n6429 9.3005
R3409 VCC.n6437 VCC.n6436 9.3005
R3410 VCC.n6436 VCC.n6204 9.3005
R3411 VCC.n6204 VCC.n6203 9.3005
R3412 VCC.n6459 VCC.n6199 9.3005
R3413 VCC.n6459 VCC.n6458 9.3005
R3414 VCC.n6458 VCC.n6457 9.3005
R3415 VCC.n6618 VCC.n6617 9.3005
R3416 VCC.n6619 VCC.n6618 9.3005
R3417 VCC.n6620 VCC.n6619 9.3005
R3418 VCC.n6564 VCC.n6563 9.3005
R3419 VCC.n6565 VCC.n6564 9.3005
R3420 VCC.n6572 VCC.n6571 9.3005
R3421 VCC.n6585 VCC.n6584 9.3005
R3422 VCC.n6585 VCC.n6137 9.3005
R3423 VCC.n6567 VCC.n6137 9.3005
R3424 VCC.n6611 VCC.n6610 9.3005
R3425 VCC.n6627 VCC.n6626 9.3005
R3426 VCC.n6626 VCC.n6103 9.3005
R3427 VCC.n6103 VCC.n6102 9.3005
R3428 VCC.n6105 VCC.n6104 9.3005
R3429 VCC.n6641 VCC.n6640 9.3005
R3430 VCC.n6520 VCC.n6519 9.3005
R3431 VCC.n6682 VCC.n6681 9.3005
R3432 VCC.n6667 VCC.n6666 9.3005
R3433 VCC.n6665 VCC.n6664 9.3005
R3434 VCC.n7137 VCC.n7136 9.3005
R3435 VCC.n7130 VCC.n7129 9.3005
R3436 VCC.n7129 VCC.n7128 9.3005
R3437 VCC.n7128 VCC.n7127 9.3005
R3438 VCC.n7190 VCC.n7189 9.3005
R3439 VCC.n7190 VCC.n6655 9.3005
R3440 VCC.n7194 VCC.n6655 9.3005
R3441 VCC.n7166 VCC.n7165 9.3005
R3442 VCC.n7165 VCC.n7164 9.3005
R3443 VCC.n7164 VCC.n7163 9.3005
R3444 VCC.n7119 VCC.n6706 9.3005
R3445 VCC.n6706 VCC.n6705 9.3005
R3446 VCC.n7077 VCC.n7076 9.3005
R3447 VCC.n7085 VCC.n7084 9.3005
R3448 VCC.n7051 VCC.n7050 9.3005
R3449 VCC.n7040 VCC.n6746 9.3005
R3450 VCC.n6749 VCC.n6748 9.3005
R3451 VCC.n6993 VCC.n6992 9.3005
R3452 VCC.n6992 VCC.n6760 9.3005
R3453 VCC.n6760 VCC.n6759 9.3005
R3454 VCC.n6762 VCC.n6761 9.3005
R3455 VCC.n7008 VCC.n7007 9.3005
R3456 VCC.n7015 VCC.n6755 9.3005
R3457 VCC.n7015 VCC.n7014 9.3005
R3458 VCC.n7014 VCC.n7013 9.3005
R3459 VCC.n7016 VCC.n6756 9.3005
R3460 VCC.n7039 VCC.n7038 9.3005
R3461 VCC.n7043 VCC.n6741 9.3005
R3462 VCC.n7044 VCC.n7043 9.3005
R3463 VCC.n7045 VCC.n7044 9.3005
R3464 VCC.n6736 VCC.n6735 9.3005
R3465 VCC.n7064 VCC.n6724 9.3005
R3466 VCC.n7064 VCC.n6734 9.3005
R3467 VCC.n6734 VCC.n6733 9.3005
R3468 VCC.n6729 VCC.n6727 9.3005
R3469 VCC.n7082 VCC.n6719 9.3005
R3470 VCC.n7082 VCC.n7081 9.3005
R3471 VCC.n7081 VCC.n7080 9.3005
R3472 VCC.n6984 VCC.n6983 9.3005
R3473 VCC.n6985 VCC.n6984 9.3005
R3474 VCC.n6986 VCC.n6985 9.3005
R3475 VCC.n6976 VCC.n6972 9.3005
R3476 VCC.n6978 VCC.n6977 9.3005
R3477 VCC.n6950 VCC.n6949 9.3005
R3478 VCC.n6925 VCC.n6924 9.3005
R3479 VCC.n6813 VCC.n6812 9.3005
R3480 VCC.n6902 VCC.n6901 9.3005
R3481 VCC.n6875 VCC.n6874 9.3005
R3482 VCC.n6875 VCC.n6831 9.3005
R3483 VCC.n6879 VCC.n6831 9.3005
R3484 VCC.n6829 VCC.n6828 9.3005
R3485 VCC.n6885 VCC.n6884 9.3005
R3486 VCC.n6822 VCC.n6821 9.3005
R3487 VCC.n6821 VCC.n6806 9.3005
R3488 VCC.n6806 VCC.n6805 9.3005
R3489 VCC.n6900 VCC.n6820 9.3005
R3490 VCC.n6814 VCC.n6808 9.3005
R3491 VCC.n6803 VCC.n6802 9.3005
R3492 VCC.n6804 VCC.n6803 9.3005
R3493 VCC.n6919 VCC.n6804 9.3005
R3494 VCC.n6797 VCC.n6796 9.3005
R3495 VCC.n6939 VCC.n6786 9.3005
R3496 VCC.n6940 VCC.n6939 9.3005
R3497 VCC.n6941 VCC.n6940 9.3005
R3498 VCC.n6791 VCC.n6789 9.3005
R3499 VCC.n6947 VCC.n6946 9.3005
R3500 VCC.n6866 VCC.n6865 9.3005
R3501 VCC.n6865 VCC.n6864 9.3005
R3502 VCC.n6864 VCC.n6863 9.3005
R3503 VCC.n6848 VCC.n6847 9.3005
R3504 VCC.n6854 VCC.n6853 9.3005
R3505 VCC.n7435 VCC.n7434 9.3005
R3506 VCC.n7404 VCC.n7403 9.3005
R3507 VCC.n7500 VCC.n7499 9.3005
R3508 VCC.n7475 VCC.n7474 9.3005
R3509 VCC.n7363 VCC.n7362 9.3005
R3510 VCC.n7364 VCC.n7358 9.3005
R3511 VCC.n7353 VCC.n7352 9.3005
R3512 VCC.n7354 VCC.n7353 9.3005
R3513 VCC.n7469 VCC.n7354 9.3005
R3514 VCC.n7347 VCC.n7346 9.3005
R3515 VCC.n7489 VCC.n7336 9.3005
R3516 VCC.n7490 VCC.n7489 9.3005
R3517 VCC.n7491 VCC.n7490 9.3005
R3518 VCC.n7341 VCC.n7339 9.3005
R3519 VCC.n7497 VCC.n7496 9.3005
R3520 VCC.n7379 VCC.n7378 9.3005
R3521 VCC.n7416 VCC.n7415 9.3005
R3522 VCC.n7415 VCC.n7414 9.3005
R3523 VCC.n7414 VCC.n7413 9.3005
R3524 VCC.n7398 VCC.n7397 9.3005
R3525 VCC.n7425 VCC.n7424 9.3005
R3526 VCC.n7425 VCC.n7381 9.3005
R3527 VCC.n7429 VCC.n7381 9.3005
R3528 VCC.n7372 VCC.n7371 9.3005
R3529 VCC.n7371 VCC.n7356 9.3005
R3530 VCC.n7356 VCC.n7355 9.3005
R3531 VCC.n7450 VCC.n7370 9.3005
R3532 VCC.n7452 VCC.n7451 9.3005
R3533 VCC.n7559 VCC.n7558 9.3005
R3534 VCC.n7529 VCC.n7528 9.3005
R3535 VCC.n7635 VCC.n7634 9.3005
R3536 VCC.n7602 VCC.n7601 9.3005
R3537 VCC.n7591 VCC.n7297 9.3005
R3538 VCC.n7590 VCC.n7589 9.3005
R3539 VCC.n7287 VCC.n7286 9.3005
R3540 VCC.n7280 VCC.n7278 9.3005
R3541 VCC.n7313 VCC.n7312 9.3005
R3542 VCC.n7527 VCC.n7522 9.3005
R3543 VCC.n7567 VCC.n7307 9.3005
R3544 VCC.n7300 VCC.n7299 9.3005
R3545 VCC.n7594 VCC.n7292 9.3005
R3546 VCC.n7595 VCC.n7594 9.3005
R3547 VCC.n7596 VCC.n7595 9.3005
R3548 VCC.n7615 VCC.n7275 9.3005
R3549 VCC.n7615 VCC.n7285 9.3005
R3550 VCC.n7285 VCC.n7284 9.3005
R3551 VCC.n7632 VCC.n7270 9.3005
R3552 VCC.n7632 VCC.n7631 9.3005
R3553 VCC.n7631 VCC.n7630 9.3005
R3554 VCC.n7535 VCC.n7534 9.3005
R3555 VCC.n7536 VCC.n7535 9.3005
R3556 VCC.n7537 VCC.n7536 9.3005
R3557 VCC.n7544 VCC.n7543 9.3005
R3558 VCC.n7543 VCC.n7311 9.3005
R3559 VCC.n7311 VCC.n7310 9.3005
R3560 VCC.n7566 VCC.n7306 9.3005
R3561 VCC.n7566 VCC.n7565 9.3005
R3562 VCC.n7565 VCC.n7564 9.3005
R3563 VCC.n7725 VCC.n7724 9.3005
R3564 VCC.n7726 VCC.n7725 9.3005
R3565 VCC.n7727 VCC.n7726 9.3005
R3566 VCC.n7671 VCC.n7670 9.3005
R3567 VCC.n7672 VCC.n7671 9.3005
R3568 VCC.n7679 VCC.n7678 9.3005
R3569 VCC.n7692 VCC.n7691 9.3005
R3570 VCC.n7692 VCC.n7244 9.3005
R3571 VCC.n7674 VCC.n7244 9.3005
R3572 VCC.n7718 VCC.n7717 9.3005
R3573 VCC.n7734 VCC.n7733 9.3005
R3574 VCC.n7733 VCC.n7210 9.3005
R3575 VCC.n7210 VCC.n7209 9.3005
R3576 VCC.n7212 VCC.n7211 9.3005
R3577 VCC.n7748 VCC.n7747 9.3005
R3578 VCC.n7627 VCC.n7626 9.3005
R3579 VCC.n7789 VCC.n7788 9.3005
R3580 VCC.n7774 VCC.n7773 9.3005
R3581 VCC.n7772 VCC.n7771 9.3005
R3582 VCC.n8244 VCC.n8243 9.3005
R3583 VCC.n8237 VCC.n8236 9.3005
R3584 VCC.n8236 VCC.n8235 9.3005
R3585 VCC.n8235 VCC.n8234 9.3005
R3586 VCC.n8297 VCC.n8296 9.3005
R3587 VCC.n8297 VCC.n7762 9.3005
R3588 VCC.n8301 VCC.n7762 9.3005
R3589 VCC.n8273 VCC.n8272 9.3005
R3590 VCC.n8272 VCC.n8271 9.3005
R3591 VCC.n8271 VCC.n8270 9.3005
R3592 VCC.n8226 VCC.n7813 9.3005
R3593 VCC.n7813 VCC.n7812 9.3005
R3594 VCC.n8184 VCC.n8183 9.3005
R3595 VCC.n8192 VCC.n8191 9.3005
R3596 VCC.n8158 VCC.n8157 9.3005
R3597 VCC.n8147 VCC.n7853 9.3005
R3598 VCC.n7856 VCC.n7855 9.3005
R3599 VCC.n8100 VCC.n8099 9.3005
R3600 VCC.n8099 VCC.n7867 9.3005
R3601 VCC.n7867 VCC.n7866 9.3005
R3602 VCC.n7869 VCC.n7868 9.3005
R3603 VCC.n8115 VCC.n8114 9.3005
R3604 VCC.n8122 VCC.n7862 9.3005
R3605 VCC.n8122 VCC.n8121 9.3005
R3606 VCC.n8121 VCC.n8120 9.3005
R3607 VCC.n8123 VCC.n7863 9.3005
R3608 VCC.n8146 VCC.n8145 9.3005
R3609 VCC.n8150 VCC.n7848 9.3005
R3610 VCC.n8151 VCC.n8150 9.3005
R3611 VCC.n8152 VCC.n8151 9.3005
R3612 VCC.n7843 VCC.n7842 9.3005
R3613 VCC.n8171 VCC.n7831 9.3005
R3614 VCC.n8171 VCC.n7841 9.3005
R3615 VCC.n7841 VCC.n7840 9.3005
R3616 VCC.n7836 VCC.n7834 9.3005
R3617 VCC.n8189 VCC.n7826 9.3005
R3618 VCC.n8189 VCC.n8188 9.3005
R3619 VCC.n8188 VCC.n8187 9.3005
R3620 VCC.n8091 VCC.n8090 9.3005
R3621 VCC.n8092 VCC.n8091 9.3005
R3622 VCC.n8093 VCC.n8092 9.3005
R3623 VCC.n8083 VCC.n8079 9.3005
R3624 VCC.n8085 VCC.n8084 9.3005
R3625 VCC.n8057 VCC.n8056 9.3005
R3626 VCC.n8032 VCC.n8031 9.3005
R3627 VCC.n7920 VCC.n7919 9.3005
R3628 VCC.n8009 VCC.n8008 9.3005
R3629 VCC.n7982 VCC.n7981 9.3005
R3630 VCC.n7982 VCC.n7938 9.3005
R3631 VCC.n7986 VCC.n7938 9.3005
R3632 VCC.n7936 VCC.n7935 9.3005
R3633 VCC.n7992 VCC.n7991 9.3005
R3634 VCC.n7929 VCC.n7928 9.3005
R3635 VCC.n7928 VCC.n7913 9.3005
R3636 VCC.n7913 VCC.n7912 9.3005
R3637 VCC.n8007 VCC.n7927 9.3005
R3638 VCC.n7921 VCC.n7915 9.3005
R3639 VCC.n7910 VCC.n7909 9.3005
R3640 VCC.n7911 VCC.n7910 9.3005
R3641 VCC.n8026 VCC.n7911 9.3005
R3642 VCC.n7904 VCC.n7903 9.3005
R3643 VCC.n8046 VCC.n7893 9.3005
R3644 VCC.n8047 VCC.n8046 9.3005
R3645 VCC.n8048 VCC.n8047 9.3005
R3646 VCC.n7898 VCC.n7896 9.3005
R3647 VCC.n8054 VCC.n8053 9.3005
R3648 VCC.n7973 VCC.n7972 9.3005
R3649 VCC.n7972 VCC.n7971 9.3005
R3650 VCC.n7971 VCC.n7970 9.3005
R3651 VCC.n7955 VCC.n7954 9.3005
R3652 VCC.n7961 VCC.n7960 9.3005
R3653 VCC.n8479 VCC.n8478 9.3005
R3654 VCC.n8449 VCC.n8448 9.3005
R3655 VCC.n8555 VCC.n8554 9.3005
R3656 VCC.n8522 VCC.n8521 9.3005
R3657 VCC.n8511 VCC.n8404 9.3005
R3658 VCC.n8510 VCC.n8509 9.3005
R3659 VCC.n8394 VCC.n8393 9.3005
R3660 VCC.n8387 VCC.n8385 9.3005
R3661 VCC.n8420 VCC.n8419 9.3005
R3662 VCC.n8447 VCC.n8442 9.3005
R3663 VCC.n8487 VCC.n8414 9.3005
R3664 VCC.n8407 VCC.n8406 9.3005
R3665 VCC.n8514 VCC.n8399 9.3005
R3666 VCC.n8515 VCC.n8514 9.3005
R3667 VCC.n8516 VCC.n8515 9.3005
R3668 VCC.n8535 VCC.n8382 9.3005
R3669 VCC.n8535 VCC.n8392 9.3005
R3670 VCC.n8392 VCC.n8391 9.3005
R3671 VCC.n8552 VCC.n8377 9.3005
R3672 VCC.n8552 VCC.n8551 9.3005
R3673 VCC.n8551 VCC.n8550 9.3005
R3674 VCC.n8455 VCC.n8454 9.3005
R3675 VCC.n8456 VCC.n8455 9.3005
R3676 VCC.n8457 VCC.n8456 9.3005
R3677 VCC.n8464 VCC.n8463 9.3005
R3678 VCC.n8463 VCC.n8418 9.3005
R3679 VCC.n8418 VCC.n8417 9.3005
R3680 VCC.n8486 VCC.n8413 9.3005
R3681 VCC.n8486 VCC.n8485 9.3005
R3682 VCC.n8485 VCC.n8484 9.3005
R3683 VCC.n8645 VCC.n8644 9.3005
R3684 VCC.n8646 VCC.n8645 9.3005
R3685 VCC.n8647 VCC.n8646 9.3005
R3686 VCC.n8591 VCC.n8590 9.3005
R3687 VCC.n8592 VCC.n8591 9.3005
R3688 VCC.n8599 VCC.n8598 9.3005
R3689 VCC.n8612 VCC.n8611 9.3005
R3690 VCC.n8612 VCC.n8351 9.3005
R3691 VCC.n8594 VCC.n8351 9.3005
R3692 VCC.n8638 VCC.n8637 9.3005
R3693 VCC.n8654 VCC.n8653 9.3005
R3694 VCC.n8653 VCC.n8317 9.3005
R3695 VCC.n8317 VCC.n8316 9.3005
R3696 VCC.n8319 VCC.n8318 9.3005
R3697 VCC.n8668 VCC.n8667 9.3005
R3698 VCC.n8547 VCC.n8546 9.3005
R3699 VCC.n210 VCC.n209 9.13511
R3700 VCC.n122 VCC.n120 9.13511
R3701 VCC.n427 VCC.n426 9.13511
R3702 VCC.n762 VCC.n761 9.13511
R3703 VCC.n674 VCC.n672 9.13511
R3704 VCC.n979 VCC.n978 9.13511
R3705 VCC.n1231 VCC.n1229 9.13511
R3706 VCC.n1537 VCC.n1536 9.13511
R3707 VCC.n1320 VCC.n1319 9.13511
R3708 VCC.n1871 VCC.n1870 9.13511
R3709 VCC.n1783 VCC.n1781 9.13511
R3710 VCC.n2088 VCC.n2087 9.13511
R3711 VCC.n2340 VCC.n2338 9.13511
R3712 VCC.n2646 VCC.n2645 9.13511
R3713 VCC.n2429 VCC.n2428 9.13511
R3714 VCC.n2980 VCC.n2979 9.13511
R3715 VCC.n2892 VCC.n2890 9.13511
R3716 VCC.n3197 VCC.n3196 9.13511
R3717 VCC.n3449 VCC.n3447 9.13511
R3718 VCC.n3755 VCC.n3754 9.13511
R3719 VCC.n3538 VCC.n3537 9.13511
R3720 VCC.n4089 VCC.n4088 9.13511
R3721 VCC.n4001 VCC.n3999 9.13511
R3722 VCC.n4306 VCC.n4305 9.13511
R3723 VCC.n4558 VCC.n4556 9.13511
R3724 VCC.n4864 VCC.n4863 9.13511
R3725 VCC.n4647 VCC.n4646 9.13511
R3726 VCC.n5198 VCC.n5197 9.13511
R3727 VCC.n5110 VCC.n5108 9.13511
R3728 VCC.n5415 VCC.n5414 9.13511
R3729 VCC.n5666 VCC.n5664 9.13511
R3730 VCC.n5972 VCC.n5971 9.13511
R3731 VCC.n5755 VCC.n5754 9.13511
R3732 VCC.n6305 VCC.n6304 9.13511
R3733 VCC.n6217 VCC.n6215 9.13511
R3734 VCC.n6522 VCC.n6521 9.13511
R3735 VCC.n6773 VCC.n6771 9.13511
R3736 VCC.n7079 VCC.n7078 9.13511
R3737 VCC.n6862 VCC.n6861 9.13511
R3738 VCC.n7412 VCC.n7411 9.13511
R3739 VCC.n7324 VCC.n7322 9.13511
R3740 VCC.n7629 VCC.n7628 9.13511
R3741 VCC.n7880 VCC.n7878 9.13511
R3742 VCC.n8186 VCC.n8185 9.13511
R3743 VCC.n7969 VCC.n7968 9.13511
R3744 VCC.n8431 VCC.n8429 9.13511
R3745 VCC.n8549 VCC.n8548 9.13511
R3746 VCC.n423 VCC.n56 8.95764
R3747 VCC.n546 VCC.n4 8.95764
R3748 VCC.n975 VCC.n608 8.95764
R3749 VCC.n1100 VCC.n558 8.95764
R3750 VCC.n1533 VCC.n1530 8.95764
R3751 VCC.n1655 VCC.n1654 8.95764
R3752 VCC.n2084 VCC.n1717 8.95764
R3753 VCC.n2209 VCC.n1667 8.95764
R3754 VCC.n2642 VCC.n2639 8.95764
R3755 VCC.n2764 VCC.n2763 8.95764
R3756 VCC.n3193 VCC.n2826 8.95764
R3757 VCC.n3318 VCC.n2776 8.95764
R3758 VCC.n3751 VCC.n3748 8.95764
R3759 VCC.n3873 VCC.n3872 8.95764
R3760 VCC.n4302 VCC.n3935 8.95764
R3761 VCC.n4427 VCC.n3885 8.95764
R3762 VCC.n4860 VCC.n4857 8.95764
R3763 VCC.n4982 VCC.n4981 8.95764
R3764 VCC.n5411 VCC.n5044 8.95764
R3765 VCC.n5536 VCC.n4994 8.95764
R3766 VCC.n5968 VCC.n5965 8.95764
R3767 VCC.n6090 VCC.n6089 8.95764
R3768 VCC.n6518 VCC.n6151 8.95764
R3769 VCC.n6643 VCC.n6101 8.95764
R3770 VCC.n7075 VCC.n7072 8.95764
R3771 VCC.n7197 VCC.n7196 8.95764
R3772 VCC.n7625 VCC.n7258 8.95764
R3773 VCC.n7750 VCC.n7208 8.95764
R3774 VCC.n8182 VCC.n8179 8.95764
R3775 VCC.n8304 VCC.n8303 8.95764
R3776 VCC.n8545 VCC.n8365 8.95764
R3777 VCC.n8670 VCC.n8315 8.95764
R3778 VCC.n499 VCC.n40 8.85536
R3779 VCC.n495 VCC.n40 8.85536
R3780 VCC.n1051 VCC.n592 8.85536
R3781 VCC.n1047 VCC.n592 8.85536
R3782 VCC.n1616 VCC.n1144 8.85536
R3783 VCC.n1144 VCC.n1143 8.85536
R3784 VCC.n2160 VCC.n1701 8.85536
R3785 VCC.n2156 VCC.n1701 8.85536
R3786 VCC.n2725 VCC.n2253 8.85536
R3787 VCC.n2253 VCC.n2252 8.85536
R3788 VCC.n3269 VCC.n2810 8.85536
R3789 VCC.n3265 VCC.n2810 8.85536
R3790 VCC.n3834 VCC.n3362 8.85536
R3791 VCC.n3362 VCC.n3361 8.85536
R3792 VCC.n4378 VCC.n3919 8.85536
R3793 VCC.n4374 VCC.n3919 8.85536
R3794 VCC.n4943 VCC.n4471 8.85536
R3795 VCC.n4471 VCC.n4470 8.85536
R3796 VCC.n5487 VCC.n5028 8.85536
R3797 VCC.n5483 VCC.n5028 8.85536
R3798 VCC.n6051 VCC.n5579 8.85536
R3799 VCC.n5579 VCC.n5578 8.85536
R3800 VCC.n6594 VCC.n6135 8.85536
R3801 VCC.n6590 VCC.n6135 8.85536
R3802 VCC.n7158 VCC.n6686 8.85536
R3803 VCC.n6686 VCC.n6685 8.85536
R3804 VCC.n7701 VCC.n7242 8.85536
R3805 VCC.n7697 VCC.n7242 8.85536
R3806 VCC.n8265 VCC.n7793 8.85536
R3807 VCC.n7793 VCC.n7792 8.85536
R3808 VCC.n8621 VCC.n8349 8.85536
R3809 VCC.n8617 VCC.n8349 8.85536
R3810 VCC.n295 VCC.n293 8.47776
R3811 VCC.n847 VCC.n845 8.47776
R3812 VCC.n1405 VCC.n1403 8.47776
R3813 VCC.n1956 VCC.n1954 8.47776
R3814 VCC.n2514 VCC.n2512 8.47776
R3815 VCC.n3065 VCC.n3063 8.47776
R3816 VCC.n3623 VCC.n3621 8.47776
R3817 VCC.n4174 VCC.n4172 8.47776
R3818 VCC.n4732 VCC.n4730 8.47776
R3819 VCC.n5283 VCC.n5281 8.47776
R3820 VCC.n5840 VCC.n5838 8.47776
R3821 VCC.n6390 VCC.n6388 8.47776
R3822 VCC.n6947 VCC.n6945 8.47776
R3823 VCC.n7497 VCC.n7495 8.47776
R3824 VCC.n8054 VCC.n8052 8.47776
R3825 VCC.n471 VCC.n470 7.03754
R3826 VCC.n527 VCC.n5 7.03754
R3827 VCC.n1023 VCC.n1022 7.03754
R3828 VCC.n1079 VCC.n559 7.03754
R3829 VCC.n1580 VCC.n1163 7.03754
R3830 VCC.n1652 VCC.n1651 7.03754
R3831 VCC.n2132 VCC.n2131 7.03754
R3832 VCC.n2188 VCC.n1668 7.03754
R3833 VCC.n2689 VCC.n2272 7.03754
R3834 VCC.n2761 VCC.n2760 7.03754
R3835 VCC.n3241 VCC.n3240 7.03754
R3836 VCC.n3297 VCC.n2777 7.03754
R3837 VCC.n3798 VCC.n3381 7.03754
R3838 VCC.n3870 VCC.n3869 7.03754
R3839 VCC.n4350 VCC.n4349 7.03754
R3840 VCC.n4406 VCC.n3886 7.03754
R3841 VCC.n4907 VCC.n4490 7.03754
R3842 VCC.n4979 VCC.n4978 7.03754
R3843 VCC.n5459 VCC.n5458 7.03754
R3844 VCC.n5515 VCC.n4995 7.03754
R3845 VCC.n6015 VCC.n5598 7.03754
R3846 VCC.n6087 VCC.n6086 7.03754
R3847 VCC.n6566 VCC.n6565 7.03754
R3848 VCC.n6622 VCC.n6102 7.03754
R3849 VCC.n7122 VCC.n6705 7.03754
R3850 VCC.n7194 VCC.n7193 7.03754
R3851 VCC.n7673 VCC.n7672 7.03754
R3852 VCC.n7729 VCC.n7209 7.03754
R3853 VCC.n8229 VCC.n7812 7.03754
R3854 VCC.n8301 VCC.n8300 7.03754
R3855 VCC.n8593 VCC.n8592 7.03754
R3856 VCC.n8649 VCC.n8316 7.03754
R3857 VCC.n226 VCC.n181 5.48127
R3858 VCC.n291 VCC.n290 5.48127
R3859 VCC.n337 VCC.n336 5.48127
R3860 VCC.n418 VCC.n417 5.48127
R3861 VCC.n778 VCC.n733 5.48127
R3862 VCC.n843 VCC.n842 5.48127
R3863 VCC.n889 VCC.n888 5.48127
R3864 VCC.n970 VCC.n969 5.48127
R3865 VCC.n1446 VCC.n1445 5.48127
R3866 VCC.n1527 VCC.n1526 5.48127
R3867 VCC.n1336 VCC.n1291 5.48127
R3868 VCC.n1401 VCC.n1400 5.48127
R3869 VCC.n1887 VCC.n1842 5.48127
R3870 VCC.n1952 VCC.n1951 5.48127
R3871 VCC.n1998 VCC.n1997 5.48127
R3872 VCC.n2079 VCC.n2078 5.48127
R3873 VCC.n2555 VCC.n2554 5.48127
R3874 VCC.n2636 VCC.n2635 5.48127
R3875 VCC.n2445 VCC.n2400 5.48127
R3876 VCC.n2510 VCC.n2509 5.48127
R3877 VCC.n2996 VCC.n2951 5.48127
R3878 VCC.n3061 VCC.n3060 5.48127
R3879 VCC.n3107 VCC.n3106 5.48127
R3880 VCC.n3188 VCC.n3187 5.48127
R3881 VCC.n3664 VCC.n3663 5.48127
R3882 VCC.n3745 VCC.n3744 5.48127
R3883 VCC.n3554 VCC.n3509 5.48127
R3884 VCC.n3619 VCC.n3618 5.48127
R3885 VCC.n4105 VCC.n4060 5.48127
R3886 VCC.n4170 VCC.n4169 5.48127
R3887 VCC.n4216 VCC.n4215 5.48127
R3888 VCC.n4297 VCC.n4296 5.48127
R3889 VCC.n4773 VCC.n4772 5.48127
R3890 VCC.n4854 VCC.n4853 5.48127
R3891 VCC.n4663 VCC.n4618 5.48127
R3892 VCC.n4728 VCC.n4727 5.48127
R3893 VCC.n5214 VCC.n5169 5.48127
R3894 VCC.n5279 VCC.n5278 5.48127
R3895 VCC.n5325 VCC.n5324 5.48127
R3896 VCC.n5406 VCC.n5405 5.48127
R3897 VCC.n5881 VCC.n5880 5.48127
R3898 VCC.n5962 VCC.n5961 5.48127
R3899 VCC.n5771 VCC.n5726 5.48127
R3900 VCC.n5836 VCC.n5835 5.48127
R3901 VCC.n6321 VCC.n6276 5.48127
R3902 VCC.n6386 VCC.n6385 5.48127
R3903 VCC.n6432 VCC.n6431 5.48127
R3904 VCC.n6513 VCC.n6512 5.48127
R3905 VCC.n6988 VCC.n6987 5.48127
R3906 VCC.n7069 VCC.n7068 5.48127
R3907 VCC.n6878 VCC.n6833 5.48127
R3908 VCC.n6943 VCC.n6942 5.48127
R3909 VCC.n7428 VCC.n7383 5.48127
R3910 VCC.n7493 VCC.n7492 5.48127
R3911 VCC.n7539 VCC.n7538 5.48127
R3912 VCC.n7620 VCC.n7619 5.48127
R3913 VCC.n8095 VCC.n8094 5.48127
R3914 VCC.n8176 VCC.n8175 5.48127
R3915 VCC.n7985 VCC.n7940 5.48127
R3916 VCC.n8050 VCC.n8049 5.48127
R3917 VCC.n8459 VCC.n8458 5.48127
R3918 VCC.n8540 VCC.n8539 5.48127
R3919 VCC.n424 VCC.n423 4.88621
R3920 VCC.n976 VCC.n975 4.88621
R3921 VCC.n1534 VCC.n1533 4.88621
R3922 VCC.n2085 VCC.n2084 4.88621
R3923 VCC.n2643 VCC.n2642 4.88621
R3924 VCC.n3194 VCC.n3193 4.88621
R3925 VCC.n3752 VCC.n3751 4.88621
R3926 VCC.n4303 VCC.n4302 4.88621
R3927 VCC.n4861 VCC.n4860 4.88621
R3928 VCC.n5412 VCC.n5411 4.88621
R3929 VCC.n5969 VCC.n5968 4.88621
R3930 VCC.n6519 VCC.n6518 4.88621
R3931 VCC.n7076 VCC.n7075 4.88621
R3932 VCC.n7626 VCC.n7625 4.88621
R3933 VCC.n8183 VCC.n8182 4.88621
R3934 VCC.n8546 VCC.n8545 4.88621
R3935 VCC.n499 VCC.n39 4.84621
R3936 VCC.n499 VCC.n498 4.84621
R3937 VCC.n1051 VCC.n591 4.84621
R3938 VCC.n1051 VCC.n1050 4.84621
R3939 VCC.n1616 VCC.n1145 4.84621
R3940 VCC.n1617 VCC.n1616 4.84621
R3941 VCC.n2160 VCC.n1700 4.84621
R3942 VCC.n2160 VCC.n2159 4.84621
R3943 VCC.n2725 VCC.n2254 4.84621
R3944 VCC.n2726 VCC.n2725 4.84621
R3945 VCC.n3269 VCC.n2809 4.84621
R3946 VCC.n3269 VCC.n3268 4.84621
R3947 VCC.n3834 VCC.n3363 4.84621
R3948 VCC.n3835 VCC.n3834 4.84621
R3949 VCC.n4378 VCC.n3918 4.84621
R3950 VCC.n4378 VCC.n4377 4.84621
R3951 VCC.n4943 VCC.n4472 4.84621
R3952 VCC.n4944 VCC.n4943 4.84621
R3953 VCC.n5487 VCC.n5027 4.84621
R3954 VCC.n5487 VCC.n5486 4.84621
R3955 VCC.n6051 VCC.n5580 4.84621
R3956 VCC.n6052 VCC.n6051 4.84621
R3957 VCC.n6594 VCC.n6134 4.84621
R3958 VCC.n6594 VCC.n6593 4.84621
R3959 VCC.n7158 VCC.n6687 4.84621
R3960 VCC.n7159 VCC.n7158 4.84621
R3961 VCC.n7701 VCC.n7241 4.84621
R3962 VCC.n7701 VCC.n7700 4.84621
R3963 VCC.n8265 VCC.n7794 4.84621
R3964 VCC.n8266 VCC.n8265 4.84621
R3965 VCC.n8621 VCC.n8348 4.84621
R3966 VCC.n8621 VCC.n8620 4.84621
R3967 VCC.n452 VCC.n57 4.6505
R3968 VCC.n1004 VCC.n609 4.6505
R3969 VCC.n1562 VCC.n1165 4.6505
R3970 VCC.n2113 VCC.n1718 4.6505
R3971 VCC.n2671 VCC.n2274 4.6505
R3972 VCC.n3222 VCC.n2827 4.6505
R3973 VCC.n3780 VCC.n3383 4.6505
R3974 VCC.n4331 VCC.n3936 4.6505
R3975 VCC.n4889 VCC.n4492 4.6505
R3976 VCC.n5440 VCC.n5045 4.6505
R3977 VCC.n5997 VCC.n5600 4.6505
R3978 VCC.n6547 VCC.n6152 4.6505
R3979 VCC.n7104 VCC.n6707 4.6505
R3980 VCC.n7654 VCC.n7259 4.6505
R3981 VCC.n8211 VCC.n7814 4.6505
R3982 VCC.n8574 VCC.n8366 4.6505
R3983 VCC.n215 VCC.n192 4.51211
R3984 VCC.n767 VCC.n744 4.51211
R3985 VCC.n1325 VCC.n1302 4.51211
R3986 VCC.n1876 VCC.n1853 4.51211
R3987 VCC.n2434 VCC.n2411 4.51211
R3988 VCC.n2985 VCC.n2962 4.51211
R3989 VCC.n3543 VCC.n3520 4.51211
R3990 VCC.n4094 VCC.n4071 4.51211
R3991 VCC.n4652 VCC.n4629 4.51211
R3992 VCC.n5203 VCC.n5180 4.51211
R3993 VCC.n5760 VCC.n5737 4.51211
R3994 VCC.n6310 VCC.n6287 4.51211
R3995 VCC.n6867 VCC.n6844 4.51211
R3996 VCC.n7417 VCC.n7394 4.51211
R3997 VCC.n7974 VCC.n7951 4.51211
R3998 VCC.n314 VCC.n125 4.51121
R3999 VCC.n866 VCC.n677 4.51121
R4000 VCC.n1424 VCC.n1234 4.51121
R4001 VCC.n1975 VCC.n1786 4.51121
R4002 VCC.n2533 VCC.n2343 4.51121
R4003 VCC.n3084 VCC.n2895 4.51121
R4004 VCC.n3642 VCC.n3452 4.51121
R4005 VCC.n4193 VCC.n4004 4.51121
R4006 VCC.n4751 VCC.n4561 4.51121
R4007 VCC.n5302 VCC.n5113 4.51121
R4008 VCC.n5859 VCC.n5669 4.51121
R4009 VCC.n6409 VCC.n6220 4.51121
R4010 VCC.n6966 VCC.n6776 4.51121
R4011 VCC.n7516 VCC.n7327 4.51121
R4012 VCC.n8073 VCC.n7883 4.51121
R4013 VCC.n8436 VCC.n8434 4.51121
R4014 VCC.n301 VCC.n135 4.5005
R4015 VCC.n300 VCC.n299 4.5005
R4016 VCC.n204 VCC.n203 4.5005
R4017 VCC.n200 VCC.n197 4.5005
R4018 VCC.n236 VCC.n175 4.5005
R4019 VCC.n246 VCC.n245 4.5005
R4020 VCC.n247 VCC.n246 4.5005
R4021 VCC.n199 VCC.n198 4.5005
R4022 VCC.n221 VCC.n174 4.5005
R4023 VCC.n221 VCC.n184 4.5005
R4024 VCC.n206 VCC.n205 4.5005
R4025 VCC.n207 VCC.n206 4.5005
R4026 VCC.n251 VCC.n166 4.5005
R4027 VCC.n251 VCC.n155 4.5005
R4028 VCC.n312 VCC.n311 4.5005
R4029 VCC.n276 VCC.n275 4.5005
R4030 VCC.n274 VCC.n146 4.5005
R4031 VCC.n254 VCC.n167 4.5005
R4032 VCC.n262 VCC.n261 4.5005
R4033 VCC.n263 VCC.n262 4.5005
R4034 VCC.n158 VCC.n148 4.5005
R4035 VCC.n159 VCC.n158 4.5005
R4036 VCC.n284 VCC.n283 4.5005
R4037 VCC.n285 VCC.n284 4.5005
R4038 VCC.n303 VCC.n302 4.5005
R4039 VCC.n138 VCC.n136 4.5005
R4040 VCC.n296 VCC.n138 4.5005
R4041 VCC.n239 VCC.n238 4.5005
R4042 VCC.n436 VCC.n74 4.5005
R4043 VCC.n435 VCC.n434 4.5005
R4044 VCC.n329 VCC.n328 4.5005
R4045 VCC.n324 VCC.n321 4.5005
R4046 VCC.n353 VCC.n352 4.5005
R4047 VCC.n323 VCC.n322 4.5005
R4048 VCC.n447 VCC.n446 4.5005
R4049 VCC.n403 VCC.n402 4.5005
R4050 VCC.n401 VCC.n86 4.5005
R4051 VCC.n438 VCC.n437 4.5005
R4052 VCC.n355 VCC.n354 4.5005
R4053 VCC.n368 VCC.n367 4.5005
R4054 VCC.n367 VCC.n366 4.5005
R4055 VCC.n117 VCC.n113 4.5005
R4056 VCC.n340 VCC.n117 4.5005
R4057 VCC.n331 VCC.n330 4.5005
R4058 VCC.n331 VCC.n124 4.5005
R4059 VCC.n383 VCC.n382 4.5005
R4060 VCC.n384 VCC.n383 4.5005
R4061 VCC.n375 VCC.n96 4.5005
R4062 VCC.n386 VCC.n96 4.5005
R4063 VCC.n390 VCC.n88 4.5005
R4064 VCC.n391 VCC.n390 4.5005
R4065 VCC.n411 VCC.n410 4.5005
R4066 VCC.n412 VCC.n411 4.5005
R4067 VCC.n77 VCC.n75 4.5005
R4068 VCC.n431 VCC.n77 4.5005
R4069 VCC.n540 VCC.n9 4.5005
R4070 VCC.n542 VCC.n541 4.5005
R4071 VCC.n519 VCC.n27 4.5005
R4072 VCC.n53 VCC.n51 4.5005
R4073 VCC.n60 VCC.n58 4.5005
R4074 VCC.n451 VCC.n450 4.5005
R4075 VCC.n456 VCC.n455 4.5005
R4076 VCC.n462 VCC.n50 4.5005
R4077 VCC.n48 VCC.n47 4.5005
R4078 VCC.n518 VCC.n517 4.5005
R4079 VCC.n509 VCC.n31 4.5005
R4080 VCC.n521 VCC.n520 4.5005
R4081 VCC.n521 VCC.n25 4.5005
R4082 VCC.n29 VCC.n16 4.5005
R4083 VCC.n17 VCC.n10 4.5005
R4084 VCC.n19 VCC.n18 4.5005
R4085 VCC.n530 VCC.n19 4.5005
R4086 VCC.n508 VCC.n507 4.5005
R4087 VCC.n38 VCC.n36 4.5005
R4088 VCC.n46 VCC.n44 4.5005
R4089 VCC.n44 VCC.n43 4.5005
R4090 VCC.n479 VCC.n478 4.5005
R4091 VCC.n467 VCC.n466 4.5005
R4092 VCC.n454 VCC.n453 4.5005
R4093 VCC.n551 VCC.n550 4.5005
R4094 VCC.n853 VCC.n687 4.5005
R4095 VCC.n852 VCC.n851 4.5005
R4096 VCC.n756 VCC.n755 4.5005
R4097 VCC.n752 VCC.n749 4.5005
R4098 VCC.n788 VCC.n727 4.5005
R4099 VCC.n798 VCC.n797 4.5005
R4100 VCC.n799 VCC.n798 4.5005
R4101 VCC.n751 VCC.n750 4.5005
R4102 VCC.n773 VCC.n726 4.5005
R4103 VCC.n773 VCC.n736 4.5005
R4104 VCC.n758 VCC.n757 4.5005
R4105 VCC.n759 VCC.n758 4.5005
R4106 VCC.n803 VCC.n718 4.5005
R4107 VCC.n803 VCC.n707 4.5005
R4108 VCC.n864 VCC.n863 4.5005
R4109 VCC.n828 VCC.n827 4.5005
R4110 VCC.n826 VCC.n698 4.5005
R4111 VCC.n806 VCC.n719 4.5005
R4112 VCC.n814 VCC.n813 4.5005
R4113 VCC.n815 VCC.n814 4.5005
R4114 VCC.n710 VCC.n700 4.5005
R4115 VCC.n711 VCC.n710 4.5005
R4116 VCC.n836 VCC.n835 4.5005
R4117 VCC.n837 VCC.n836 4.5005
R4118 VCC.n855 VCC.n854 4.5005
R4119 VCC.n690 VCC.n688 4.5005
R4120 VCC.n848 VCC.n690 4.5005
R4121 VCC.n791 VCC.n790 4.5005
R4122 VCC.n988 VCC.n626 4.5005
R4123 VCC.n987 VCC.n986 4.5005
R4124 VCC.n881 VCC.n880 4.5005
R4125 VCC.n876 VCC.n873 4.5005
R4126 VCC.n905 VCC.n904 4.5005
R4127 VCC.n875 VCC.n874 4.5005
R4128 VCC.n999 VCC.n998 4.5005
R4129 VCC.n955 VCC.n954 4.5005
R4130 VCC.n953 VCC.n638 4.5005
R4131 VCC.n990 VCC.n989 4.5005
R4132 VCC.n907 VCC.n906 4.5005
R4133 VCC.n920 VCC.n919 4.5005
R4134 VCC.n919 VCC.n918 4.5005
R4135 VCC.n669 VCC.n665 4.5005
R4136 VCC.n892 VCC.n669 4.5005
R4137 VCC.n883 VCC.n882 4.5005
R4138 VCC.n883 VCC.n676 4.5005
R4139 VCC.n935 VCC.n934 4.5005
R4140 VCC.n936 VCC.n935 4.5005
R4141 VCC.n927 VCC.n648 4.5005
R4142 VCC.n938 VCC.n648 4.5005
R4143 VCC.n942 VCC.n640 4.5005
R4144 VCC.n943 VCC.n942 4.5005
R4145 VCC.n963 VCC.n962 4.5005
R4146 VCC.n964 VCC.n963 4.5005
R4147 VCC.n629 VCC.n627 4.5005
R4148 VCC.n983 VCC.n629 4.5005
R4149 VCC.n569 VCC.n564 4.5005
R4150 VCC.n1096 VCC.n1095 4.5005
R4151 VCC.n1006 VCC.n1005 4.5005
R4152 VCC.n612 VCC.n610 4.5005
R4153 VCC.n1031 VCC.n1030 4.5005
R4154 VCC.n598 VCC.n596 4.5005
R4155 VCC.n596 VCC.n595 4.5005
R4156 VCC.n600 VCC.n599 4.5005
R4157 VCC.n1014 VCC.n602 4.5005
R4158 VCC.n1019 VCC.n1018 4.5005
R4159 VCC.n1003 VCC.n1002 4.5005
R4160 VCC.n1008 VCC.n1007 4.5005
R4161 VCC.n571 VCC.n570 4.5005
R4162 VCC.n1082 VCC.n571 4.5005
R4163 VCC.n1070 VCC.n1069 4.5005
R4164 VCC.n581 VCC.n568 4.5005
R4165 VCC.n1060 VCC.n1059 4.5005
R4166 VCC.n590 VCC.n588 4.5005
R4167 VCC.n1061 VCC.n583 4.5005
R4168 VCC.n1071 VCC.n579 4.5005
R4169 VCC.n1073 VCC.n1072 4.5005
R4170 VCC.n1073 VCC.n577 4.5005
R4171 VCC.n1094 VCC.n563 4.5005
R4172 VCC.n1105 VCC.n1104 4.5005
R4173 VCC.n605 VCC.n603 4.5005
R4174 VCC.n1564 VCC.n1166 4.5005
R4175 VCC.n1567 VCC.n1566 4.5005
R4176 VCC.n1641 VCC.n1121 4.5005
R4177 VCC.n1643 VCC.n1642 4.5005
R4178 VCC.n1138 VCC.n1137 4.5005
R4179 VCC.n1158 VCC.n1156 4.5005
R4180 VCC.n1168 VCC.n1155 4.5005
R4181 VCC.n1597 VCC.n1596 4.5005
R4182 VCC.n1606 VCC.n1605 4.5005
R4183 VCC.n1149 VCC.n1148 4.5005
R4184 VCC.n1129 VCC.n1128 4.5005
R4185 VCC.n1632 VCC.n1631 4.5005
R4186 VCC.n1644 VCC.n1119 4.5005
R4187 VCC.n1133 VCC.n1131 4.5005
R4188 VCC.n1604 VCC.n1603 4.5005
R4189 VCC.n1565 VCC.n1563 4.5005
R4190 VCC.n1561 VCC.n1560 4.5005
R4191 VCC.n1576 VCC.n1167 4.5005
R4192 VCC.n1646 VCC.n1645 4.5005
R4193 VCC.n1646 VCC.n1117 4.5005
R4194 VCC.n1136 VCC.n1134 4.5005
R4195 VCC.n1141 VCC.n1134 4.5005
R4196 VCC.n1592 VCC.n1591 4.5005
R4197 VCC.n1593 VCC.n1592 4.5005
R4198 VCC.n1659 VCC.n1658 4.5005
R4199 VCC.n1546 VCC.n1183 4.5005
R4200 VCC.n1545 VCC.n1544 4.5005
R4201 VCC.n1510 VCC.n1195 4.5005
R4202 VCC.n1464 VCC.n1463 4.5005
R4203 VCC.n1438 VCC.n1437 4.5005
R4204 VCC.n1433 VCC.n1429 4.5005
R4205 VCC.n1439 VCC.n1235 4.5005
R4206 VCC.n1235 VCC.n1233 4.5005
R4207 VCC.n1557 VCC.n1556 4.5005
R4208 VCC.n1512 VCC.n1511 4.5005
R4209 VCC.n1432 VCC.n1431 4.5005
R4210 VCC.n1226 VCC.n1222 4.5005
R4211 VCC.n1449 VCC.n1226 4.5005
R4212 VCC.n1462 VCC.n1461 4.5005
R4213 VCC.n1477 VCC.n1476 4.5005
R4214 VCC.n1476 VCC.n1475 4.5005
R4215 VCC.n1492 VCC.n1491 4.5005
R4216 VCC.n1493 VCC.n1492 4.5005
R4217 VCC.n1484 VCC.n1205 4.5005
R4218 VCC.n1495 VCC.n1205 4.5005
R4219 VCC.n1499 VCC.n1197 4.5005
R4220 VCC.n1500 VCC.n1499 4.5005
R4221 VCC.n1520 VCC.n1519 4.5005
R4222 VCC.n1521 VCC.n1520 4.5005
R4223 VCC.n1548 VCC.n1547 4.5005
R4224 VCC.n1186 VCC.n1184 4.5005
R4225 VCC.n1541 VCC.n1186 4.5005
R4226 VCC.n1411 VCC.n1245 4.5005
R4227 VCC.n1410 VCC.n1409 4.5005
R4228 VCC.n1384 VCC.n1256 4.5005
R4229 VCC.n1349 VCC.n1348 4.5005
R4230 VCC.n1314 VCC.n1313 4.5005
R4231 VCC.n1310 VCC.n1307 4.5005
R4232 VCC.n1316 VCC.n1315 4.5005
R4233 VCC.n1317 VCC.n1316 4.5005
R4234 VCC.n1422 VCC.n1421 4.5005
R4235 VCC.n1386 VCC.n1385 4.5005
R4236 VCC.n1309 VCC.n1308 4.5005
R4237 VCC.n1331 VCC.n1284 4.5005
R4238 VCC.n1331 VCC.n1294 4.5005
R4239 VCC.n1346 VCC.n1285 4.5005
R4240 VCC.n1356 VCC.n1355 4.5005
R4241 VCC.n1357 VCC.n1356 4.5005
R4242 VCC.n1361 VCC.n1276 4.5005
R4243 VCC.n1361 VCC.n1265 4.5005
R4244 VCC.n1364 VCC.n1277 4.5005
R4245 VCC.n1372 VCC.n1371 4.5005
R4246 VCC.n1373 VCC.n1372 4.5005
R4247 VCC.n1268 VCC.n1258 4.5005
R4248 VCC.n1269 VCC.n1268 4.5005
R4249 VCC.n1394 VCC.n1393 4.5005
R4250 VCC.n1395 VCC.n1394 4.5005
R4251 VCC.n1413 VCC.n1412 4.5005
R4252 VCC.n1248 VCC.n1246 4.5005
R4253 VCC.n1406 VCC.n1248 4.5005
R4254 VCC.n1962 VCC.n1796 4.5005
R4255 VCC.n1961 VCC.n1960 4.5005
R4256 VCC.n1865 VCC.n1864 4.5005
R4257 VCC.n1861 VCC.n1858 4.5005
R4258 VCC.n1897 VCC.n1836 4.5005
R4259 VCC.n1907 VCC.n1906 4.5005
R4260 VCC.n1908 VCC.n1907 4.5005
R4261 VCC.n1860 VCC.n1859 4.5005
R4262 VCC.n1882 VCC.n1835 4.5005
R4263 VCC.n1882 VCC.n1845 4.5005
R4264 VCC.n1867 VCC.n1866 4.5005
R4265 VCC.n1868 VCC.n1867 4.5005
R4266 VCC.n1912 VCC.n1827 4.5005
R4267 VCC.n1912 VCC.n1816 4.5005
R4268 VCC.n1973 VCC.n1972 4.5005
R4269 VCC.n1937 VCC.n1936 4.5005
R4270 VCC.n1935 VCC.n1807 4.5005
R4271 VCC.n1915 VCC.n1828 4.5005
R4272 VCC.n1923 VCC.n1922 4.5005
R4273 VCC.n1924 VCC.n1923 4.5005
R4274 VCC.n1819 VCC.n1809 4.5005
R4275 VCC.n1820 VCC.n1819 4.5005
R4276 VCC.n1945 VCC.n1944 4.5005
R4277 VCC.n1946 VCC.n1945 4.5005
R4278 VCC.n1964 VCC.n1963 4.5005
R4279 VCC.n1799 VCC.n1797 4.5005
R4280 VCC.n1957 VCC.n1799 4.5005
R4281 VCC.n1900 VCC.n1899 4.5005
R4282 VCC.n2097 VCC.n1735 4.5005
R4283 VCC.n2096 VCC.n2095 4.5005
R4284 VCC.n1990 VCC.n1989 4.5005
R4285 VCC.n1985 VCC.n1982 4.5005
R4286 VCC.n2014 VCC.n2013 4.5005
R4287 VCC.n1984 VCC.n1983 4.5005
R4288 VCC.n2108 VCC.n2107 4.5005
R4289 VCC.n2064 VCC.n2063 4.5005
R4290 VCC.n2062 VCC.n1747 4.5005
R4291 VCC.n2099 VCC.n2098 4.5005
R4292 VCC.n2016 VCC.n2015 4.5005
R4293 VCC.n2029 VCC.n2028 4.5005
R4294 VCC.n2028 VCC.n2027 4.5005
R4295 VCC.n1778 VCC.n1774 4.5005
R4296 VCC.n2001 VCC.n1778 4.5005
R4297 VCC.n1992 VCC.n1991 4.5005
R4298 VCC.n1992 VCC.n1785 4.5005
R4299 VCC.n2044 VCC.n2043 4.5005
R4300 VCC.n2045 VCC.n2044 4.5005
R4301 VCC.n2036 VCC.n1757 4.5005
R4302 VCC.n2047 VCC.n1757 4.5005
R4303 VCC.n2051 VCC.n1749 4.5005
R4304 VCC.n2052 VCC.n2051 4.5005
R4305 VCC.n2072 VCC.n2071 4.5005
R4306 VCC.n2073 VCC.n2072 4.5005
R4307 VCC.n1738 VCC.n1736 4.5005
R4308 VCC.n2092 VCC.n1738 4.5005
R4309 VCC.n1678 VCC.n1673 4.5005
R4310 VCC.n2205 VCC.n2204 4.5005
R4311 VCC.n2115 VCC.n2114 4.5005
R4312 VCC.n1721 VCC.n1719 4.5005
R4313 VCC.n2140 VCC.n2139 4.5005
R4314 VCC.n1707 VCC.n1705 4.5005
R4315 VCC.n1705 VCC.n1704 4.5005
R4316 VCC.n1709 VCC.n1708 4.5005
R4317 VCC.n2123 VCC.n1711 4.5005
R4318 VCC.n2128 VCC.n2127 4.5005
R4319 VCC.n2112 VCC.n2111 4.5005
R4320 VCC.n2117 VCC.n2116 4.5005
R4321 VCC.n1680 VCC.n1679 4.5005
R4322 VCC.n2191 VCC.n1680 4.5005
R4323 VCC.n2179 VCC.n2178 4.5005
R4324 VCC.n1690 VCC.n1677 4.5005
R4325 VCC.n2169 VCC.n2168 4.5005
R4326 VCC.n1699 VCC.n1697 4.5005
R4327 VCC.n2170 VCC.n1692 4.5005
R4328 VCC.n2180 VCC.n1688 4.5005
R4329 VCC.n2182 VCC.n2181 4.5005
R4330 VCC.n2182 VCC.n1686 4.5005
R4331 VCC.n2203 VCC.n1672 4.5005
R4332 VCC.n2214 VCC.n2213 4.5005
R4333 VCC.n1714 VCC.n1712 4.5005
R4334 VCC.n2673 VCC.n2275 4.5005
R4335 VCC.n2676 VCC.n2675 4.5005
R4336 VCC.n2750 VCC.n2230 4.5005
R4337 VCC.n2752 VCC.n2751 4.5005
R4338 VCC.n2247 VCC.n2246 4.5005
R4339 VCC.n2267 VCC.n2265 4.5005
R4340 VCC.n2277 VCC.n2264 4.5005
R4341 VCC.n2706 VCC.n2705 4.5005
R4342 VCC.n2715 VCC.n2714 4.5005
R4343 VCC.n2258 VCC.n2257 4.5005
R4344 VCC.n2238 VCC.n2237 4.5005
R4345 VCC.n2741 VCC.n2740 4.5005
R4346 VCC.n2753 VCC.n2228 4.5005
R4347 VCC.n2242 VCC.n2240 4.5005
R4348 VCC.n2713 VCC.n2712 4.5005
R4349 VCC.n2674 VCC.n2672 4.5005
R4350 VCC.n2670 VCC.n2669 4.5005
R4351 VCC.n2685 VCC.n2276 4.5005
R4352 VCC.n2755 VCC.n2754 4.5005
R4353 VCC.n2755 VCC.n2226 4.5005
R4354 VCC.n2245 VCC.n2243 4.5005
R4355 VCC.n2250 VCC.n2243 4.5005
R4356 VCC.n2701 VCC.n2700 4.5005
R4357 VCC.n2702 VCC.n2701 4.5005
R4358 VCC.n2768 VCC.n2767 4.5005
R4359 VCC.n2655 VCC.n2292 4.5005
R4360 VCC.n2654 VCC.n2653 4.5005
R4361 VCC.n2619 VCC.n2304 4.5005
R4362 VCC.n2573 VCC.n2572 4.5005
R4363 VCC.n2547 VCC.n2546 4.5005
R4364 VCC.n2542 VCC.n2538 4.5005
R4365 VCC.n2548 VCC.n2344 4.5005
R4366 VCC.n2344 VCC.n2342 4.5005
R4367 VCC.n2666 VCC.n2665 4.5005
R4368 VCC.n2621 VCC.n2620 4.5005
R4369 VCC.n2541 VCC.n2540 4.5005
R4370 VCC.n2335 VCC.n2331 4.5005
R4371 VCC.n2558 VCC.n2335 4.5005
R4372 VCC.n2571 VCC.n2570 4.5005
R4373 VCC.n2586 VCC.n2585 4.5005
R4374 VCC.n2585 VCC.n2584 4.5005
R4375 VCC.n2601 VCC.n2600 4.5005
R4376 VCC.n2602 VCC.n2601 4.5005
R4377 VCC.n2593 VCC.n2314 4.5005
R4378 VCC.n2604 VCC.n2314 4.5005
R4379 VCC.n2608 VCC.n2306 4.5005
R4380 VCC.n2609 VCC.n2608 4.5005
R4381 VCC.n2629 VCC.n2628 4.5005
R4382 VCC.n2630 VCC.n2629 4.5005
R4383 VCC.n2657 VCC.n2656 4.5005
R4384 VCC.n2295 VCC.n2293 4.5005
R4385 VCC.n2650 VCC.n2295 4.5005
R4386 VCC.n2520 VCC.n2354 4.5005
R4387 VCC.n2519 VCC.n2518 4.5005
R4388 VCC.n2493 VCC.n2365 4.5005
R4389 VCC.n2458 VCC.n2457 4.5005
R4390 VCC.n2423 VCC.n2422 4.5005
R4391 VCC.n2419 VCC.n2416 4.5005
R4392 VCC.n2425 VCC.n2424 4.5005
R4393 VCC.n2426 VCC.n2425 4.5005
R4394 VCC.n2531 VCC.n2530 4.5005
R4395 VCC.n2495 VCC.n2494 4.5005
R4396 VCC.n2418 VCC.n2417 4.5005
R4397 VCC.n2440 VCC.n2393 4.5005
R4398 VCC.n2440 VCC.n2403 4.5005
R4399 VCC.n2455 VCC.n2394 4.5005
R4400 VCC.n2465 VCC.n2464 4.5005
R4401 VCC.n2466 VCC.n2465 4.5005
R4402 VCC.n2470 VCC.n2385 4.5005
R4403 VCC.n2470 VCC.n2374 4.5005
R4404 VCC.n2473 VCC.n2386 4.5005
R4405 VCC.n2481 VCC.n2480 4.5005
R4406 VCC.n2482 VCC.n2481 4.5005
R4407 VCC.n2377 VCC.n2367 4.5005
R4408 VCC.n2378 VCC.n2377 4.5005
R4409 VCC.n2503 VCC.n2502 4.5005
R4410 VCC.n2504 VCC.n2503 4.5005
R4411 VCC.n2522 VCC.n2521 4.5005
R4412 VCC.n2357 VCC.n2355 4.5005
R4413 VCC.n2515 VCC.n2357 4.5005
R4414 VCC.n3071 VCC.n2905 4.5005
R4415 VCC.n3070 VCC.n3069 4.5005
R4416 VCC.n2974 VCC.n2973 4.5005
R4417 VCC.n2970 VCC.n2967 4.5005
R4418 VCC.n3006 VCC.n2945 4.5005
R4419 VCC.n3016 VCC.n3015 4.5005
R4420 VCC.n3017 VCC.n3016 4.5005
R4421 VCC.n2969 VCC.n2968 4.5005
R4422 VCC.n2991 VCC.n2944 4.5005
R4423 VCC.n2991 VCC.n2954 4.5005
R4424 VCC.n2976 VCC.n2975 4.5005
R4425 VCC.n2977 VCC.n2976 4.5005
R4426 VCC.n3021 VCC.n2936 4.5005
R4427 VCC.n3021 VCC.n2925 4.5005
R4428 VCC.n3082 VCC.n3081 4.5005
R4429 VCC.n3046 VCC.n3045 4.5005
R4430 VCC.n3044 VCC.n2916 4.5005
R4431 VCC.n3024 VCC.n2937 4.5005
R4432 VCC.n3032 VCC.n3031 4.5005
R4433 VCC.n3033 VCC.n3032 4.5005
R4434 VCC.n2928 VCC.n2918 4.5005
R4435 VCC.n2929 VCC.n2928 4.5005
R4436 VCC.n3054 VCC.n3053 4.5005
R4437 VCC.n3055 VCC.n3054 4.5005
R4438 VCC.n3073 VCC.n3072 4.5005
R4439 VCC.n2908 VCC.n2906 4.5005
R4440 VCC.n3066 VCC.n2908 4.5005
R4441 VCC.n3009 VCC.n3008 4.5005
R4442 VCC.n3206 VCC.n2844 4.5005
R4443 VCC.n3205 VCC.n3204 4.5005
R4444 VCC.n3099 VCC.n3098 4.5005
R4445 VCC.n3094 VCC.n3091 4.5005
R4446 VCC.n3123 VCC.n3122 4.5005
R4447 VCC.n3093 VCC.n3092 4.5005
R4448 VCC.n3217 VCC.n3216 4.5005
R4449 VCC.n3173 VCC.n3172 4.5005
R4450 VCC.n3171 VCC.n2856 4.5005
R4451 VCC.n3208 VCC.n3207 4.5005
R4452 VCC.n3125 VCC.n3124 4.5005
R4453 VCC.n3138 VCC.n3137 4.5005
R4454 VCC.n3137 VCC.n3136 4.5005
R4455 VCC.n2887 VCC.n2883 4.5005
R4456 VCC.n3110 VCC.n2887 4.5005
R4457 VCC.n3101 VCC.n3100 4.5005
R4458 VCC.n3101 VCC.n2894 4.5005
R4459 VCC.n3153 VCC.n3152 4.5005
R4460 VCC.n3154 VCC.n3153 4.5005
R4461 VCC.n3145 VCC.n2866 4.5005
R4462 VCC.n3156 VCC.n2866 4.5005
R4463 VCC.n3160 VCC.n2858 4.5005
R4464 VCC.n3161 VCC.n3160 4.5005
R4465 VCC.n3181 VCC.n3180 4.5005
R4466 VCC.n3182 VCC.n3181 4.5005
R4467 VCC.n2847 VCC.n2845 4.5005
R4468 VCC.n3201 VCC.n2847 4.5005
R4469 VCC.n2787 VCC.n2782 4.5005
R4470 VCC.n3314 VCC.n3313 4.5005
R4471 VCC.n3224 VCC.n3223 4.5005
R4472 VCC.n2830 VCC.n2828 4.5005
R4473 VCC.n3249 VCC.n3248 4.5005
R4474 VCC.n2816 VCC.n2814 4.5005
R4475 VCC.n2814 VCC.n2813 4.5005
R4476 VCC.n2818 VCC.n2817 4.5005
R4477 VCC.n3232 VCC.n2820 4.5005
R4478 VCC.n3237 VCC.n3236 4.5005
R4479 VCC.n3221 VCC.n3220 4.5005
R4480 VCC.n3226 VCC.n3225 4.5005
R4481 VCC.n2789 VCC.n2788 4.5005
R4482 VCC.n3300 VCC.n2789 4.5005
R4483 VCC.n3288 VCC.n3287 4.5005
R4484 VCC.n2799 VCC.n2786 4.5005
R4485 VCC.n3278 VCC.n3277 4.5005
R4486 VCC.n2808 VCC.n2806 4.5005
R4487 VCC.n3279 VCC.n2801 4.5005
R4488 VCC.n3289 VCC.n2797 4.5005
R4489 VCC.n3291 VCC.n3290 4.5005
R4490 VCC.n3291 VCC.n2795 4.5005
R4491 VCC.n3312 VCC.n2781 4.5005
R4492 VCC.n3323 VCC.n3322 4.5005
R4493 VCC.n2823 VCC.n2821 4.5005
R4494 VCC.n3782 VCC.n3384 4.5005
R4495 VCC.n3785 VCC.n3784 4.5005
R4496 VCC.n3859 VCC.n3339 4.5005
R4497 VCC.n3861 VCC.n3860 4.5005
R4498 VCC.n3356 VCC.n3355 4.5005
R4499 VCC.n3376 VCC.n3374 4.5005
R4500 VCC.n3386 VCC.n3373 4.5005
R4501 VCC.n3815 VCC.n3814 4.5005
R4502 VCC.n3824 VCC.n3823 4.5005
R4503 VCC.n3367 VCC.n3366 4.5005
R4504 VCC.n3347 VCC.n3346 4.5005
R4505 VCC.n3850 VCC.n3849 4.5005
R4506 VCC.n3862 VCC.n3337 4.5005
R4507 VCC.n3351 VCC.n3349 4.5005
R4508 VCC.n3822 VCC.n3821 4.5005
R4509 VCC.n3783 VCC.n3781 4.5005
R4510 VCC.n3779 VCC.n3778 4.5005
R4511 VCC.n3794 VCC.n3385 4.5005
R4512 VCC.n3864 VCC.n3863 4.5005
R4513 VCC.n3864 VCC.n3335 4.5005
R4514 VCC.n3354 VCC.n3352 4.5005
R4515 VCC.n3359 VCC.n3352 4.5005
R4516 VCC.n3810 VCC.n3809 4.5005
R4517 VCC.n3811 VCC.n3810 4.5005
R4518 VCC.n3877 VCC.n3876 4.5005
R4519 VCC.n3764 VCC.n3401 4.5005
R4520 VCC.n3763 VCC.n3762 4.5005
R4521 VCC.n3728 VCC.n3413 4.5005
R4522 VCC.n3682 VCC.n3681 4.5005
R4523 VCC.n3656 VCC.n3655 4.5005
R4524 VCC.n3651 VCC.n3647 4.5005
R4525 VCC.n3657 VCC.n3453 4.5005
R4526 VCC.n3453 VCC.n3451 4.5005
R4527 VCC.n3775 VCC.n3774 4.5005
R4528 VCC.n3730 VCC.n3729 4.5005
R4529 VCC.n3650 VCC.n3649 4.5005
R4530 VCC.n3444 VCC.n3440 4.5005
R4531 VCC.n3667 VCC.n3444 4.5005
R4532 VCC.n3680 VCC.n3679 4.5005
R4533 VCC.n3695 VCC.n3694 4.5005
R4534 VCC.n3694 VCC.n3693 4.5005
R4535 VCC.n3710 VCC.n3709 4.5005
R4536 VCC.n3711 VCC.n3710 4.5005
R4537 VCC.n3702 VCC.n3423 4.5005
R4538 VCC.n3713 VCC.n3423 4.5005
R4539 VCC.n3717 VCC.n3415 4.5005
R4540 VCC.n3718 VCC.n3717 4.5005
R4541 VCC.n3738 VCC.n3737 4.5005
R4542 VCC.n3739 VCC.n3738 4.5005
R4543 VCC.n3766 VCC.n3765 4.5005
R4544 VCC.n3404 VCC.n3402 4.5005
R4545 VCC.n3759 VCC.n3404 4.5005
R4546 VCC.n3629 VCC.n3463 4.5005
R4547 VCC.n3628 VCC.n3627 4.5005
R4548 VCC.n3602 VCC.n3474 4.5005
R4549 VCC.n3567 VCC.n3566 4.5005
R4550 VCC.n3532 VCC.n3531 4.5005
R4551 VCC.n3528 VCC.n3525 4.5005
R4552 VCC.n3534 VCC.n3533 4.5005
R4553 VCC.n3535 VCC.n3534 4.5005
R4554 VCC.n3640 VCC.n3639 4.5005
R4555 VCC.n3604 VCC.n3603 4.5005
R4556 VCC.n3527 VCC.n3526 4.5005
R4557 VCC.n3549 VCC.n3502 4.5005
R4558 VCC.n3549 VCC.n3512 4.5005
R4559 VCC.n3564 VCC.n3503 4.5005
R4560 VCC.n3574 VCC.n3573 4.5005
R4561 VCC.n3575 VCC.n3574 4.5005
R4562 VCC.n3579 VCC.n3494 4.5005
R4563 VCC.n3579 VCC.n3483 4.5005
R4564 VCC.n3582 VCC.n3495 4.5005
R4565 VCC.n3590 VCC.n3589 4.5005
R4566 VCC.n3591 VCC.n3590 4.5005
R4567 VCC.n3486 VCC.n3476 4.5005
R4568 VCC.n3487 VCC.n3486 4.5005
R4569 VCC.n3612 VCC.n3611 4.5005
R4570 VCC.n3613 VCC.n3612 4.5005
R4571 VCC.n3631 VCC.n3630 4.5005
R4572 VCC.n3466 VCC.n3464 4.5005
R4573 VCC.n3624 VCC.n3466 4.5005
R4574 VCC.n4180 VCC.n4014 4.5005
R4575 VCC.n4179 VCC.n4178 4.5005
R4576 VCC.n4083 VCC.n4082 4.5005
R4577 VCC.n4079 VCC.n4076 4.5005
R4578 VCC.n4115 VCC.n4054 4.5005
R4579 VCC.n4125 VCC.n4124 4.5005
R4580 VCC.n4126 VCC.n4125 4.5005
R4581 VCC.n4078 VCC.n4077 4.5005
R4582 VCC.n4100 VCC.n4053 4.5005
R4583 VCC.n4100 VCC.n4063 4.5005
R4584 VCC.n4085 VCC.n4084 4.5005
R4585 VCC.n4086 VCC.n4085 4.5005
R4586 VCC.n4130 VCC.n4045 4.5005
R4587 VCC.n4130 VCC.n4034 4.5005
R4588 VCC.n4191 VCC.n4190 4.5005
R4589 VCC.n4155 VCC.n4154 4.5005
R4590 VCC.n4153 VCC.n4025 4.5005
R4591 VCC.n4133 VCC.n4046 4.5005
R4592 VCC.n4141 VCC.n4140 4.5005
R4593 VCC.n4142 VCC.n4141 4.5005
R4594 VCC.n4037 VCC.n4027 4.5005
R4595 VCC.n4038 VCC.n4037 4.5005
R4596 VCC.n4163 VCC.n4162 4.5005
R4597 VCC.n4164 VCC.n4163 4.5005
R4598 VCC.n4182 VCC.n4181 4.5005
R4599 VCC.n4017 VCC.n4015 4.5005
R4600 VCC.n4175 VCC.n4017 4.5005
R4601 VCC.n4118 VCC.n4117 4.5005
R4602 VCC.n4315 VCC.n3953 4.5005
R4603 VCC.n4314 VCC.n4313 4.5005
R4604 VCC.n4208 VCC.n4207 4.5005
R4605 VCC.n4203 VCC.n4200 4.5005
R4606 VCC.n4232 VCC.n4231 4.5005
R4607 VCC.n4202 VCC.n4201 4.5005
R4608 VCC.n4326 VCC.n4325 4.5005
R4609 VCC.n4282 VCC.n4281 4.5005
R4610 VCC.n4280 VCC.n3965 4.5005
R4611 VCC.n4317 VCC.n4316 4.5005
R4612 VCC.n4234 VCC.n4233 4.5005
R4613 VCC.n4247 VCC.n4246 4.5005
R4614 VCC.n4246 VCC.n4245 4.5005
R4615 VCC.n3996 VCC.n3992 4.5005
R4616 VCC.n4219 VCC.n3996 4.5005
R4617 VCC.n4210 VCC.n4209 4.5005
R4618 VCC.n4210 VCC.n4003 4.5005
R4619 VCC.n4262 VCC.n4261 4.5005
R4620 VCC.n4263 VCC.n4262 4.5005
R4621 VCC.n4254 VCC.n3975 4.5005
R4622 VCC.n4265 VCC.n3975 4.5005
R4623 VCC.n4269 VCC.n3967 4.5005
R4624 VCC.n4270 VCC.n4269 4.5005
R4625 VCC.n4290 VCC.n4289 4.5005
R4626 VCC.n4291 VCC.n4290 4.5005
R4627 VCC.n3956 VCC.n3954 4.5005
R4628 VCC.n4310 VCC.n3956 4.5005
R4629 VCC.n3896 VCC.n3891 4.5005
R4630 VCC.n4423 VCC.n4422 4.5005
R4631 VCC.n4333 VCC.n4332 4.5005
R4632 VCC.n3939 VCC.n3937 4.5005
R4633 VCC.n4358 VCC.n4357 4.5005
R4634 VCC.n3925 VCC.n3923 4.5005
R4635 VCC.n3923 VCC.n3922 4.5005
R4636 VCC.n3927 VCC.n3926 4.5005
R4637 VCC.n4341 VCC.n3929 4.5005
R4638 VCC.n4346 VCC.n4345 4.5005
R4639 VCC.n4330 VCC.n4329 4.5005
R4640 VCC.n4335 VCC.n4334 4.5005
R4641 VCC.n3898 VCC.n3897 4.5005
R4642 VCC.n4409 VCC.n3898 4.5005
R4643 VCC.n4397 VCC.n4396 4.5005
R4644 VCC.n3908 VCC.n3895 4.5005
R4645 VCC.n4387 VCC.n4386 4.5005
R4646 VCC.n3917 VCC.n3915 4.5005
R4647 VCC.n4388 VCC.n3910 4.5005
R4648 VCC.n4398 VCC.n3906 4.5005
R4649 VCC.n4400 VCC.n4399 4.5005
R4650 VCC.n4400 VCC.n3904 4.5005
R4651 VCC.n4421 VCC.n3890 4.5005
R4652 VCC.n4432 VCC.n4431 4.5005
R4653 VCC.n3932 VCC.n3930 4.5005
R4654 VCC.n4891 VCC.n4493 4.5005
R4655 VCC.n4894 VCC.n4893 4.5005
R4656 VCC.n4968 VCC.n4448 4.5005
R4657 VCC.n4970 VCC.n4969 4.5005
R4658 VCC.n4465 VCC.n4464 4.5005
R4659 VCC.n4485 VCC.n4483 4.5005
R4660 VCC.n4495 VCC.n4482 4.5005
R4661 VCC.n4924 VCC.n4923 4.5005
R4662 VCC.n4933 VCC.n4932 4.5005
R4663 VCC.n4476 VCC.n4475 4.5005
R4664 VCC.n4456 VCC.n4455 4.5005
R4665 VCC.n4959 VCC.n4958 4.5005
R4666 VCC.n4971 VCC.n4446 4.5005
R4667 VCC.n4460 VCC.n4458 4.5005
R4668 VCC.n4931 VCC.n4930 4.5005
R4669 VCC.n4892 VCC.n4890 4.5005
R4670 VCC.n4888 VCC.n4887 4.5005
R4671 VCC.n4903 VCC.n4494 4.5005
R4672 VCC.n4973 VCC.n4972 4.5005
R4673 VCC.n4973 VCC.n4444 4.5005
R4674 VCC.n4463 VCC.n4461 4.5005
R4675 VCC.n4468 VCC.n4461 4.5005
R4676 VCC.n4919 VCC.n4918 4.5005
R4677 VCC.n4920 VCC.n4919 4.5005
R4678 VCC.n4986 VCC.n4985 4.5005
R4679 VCC.n4873 VCC.n4510 4.5005
R4680 VCC.n4872 VCC.n4871 4.5005
R4681 VCC.n4837 VCC.n4522 4.5005
R4682 VCC.n4791 VCC.n4790 4.5005
R4683 VCC.n4765 VCC.n4764 4.5005
R4684 VCC.n4760 VCC.n4756 4.5005
R4685 VCC.n4766 VCC.n4562 4.5005
R4686 VCC.n4562 VCC.n4560 4.5005
R4687 VCC.n4884 VCC.n4883 4.5005
R4688 VCC.n4839 VCC.n4838 4.5005
R4689 VCC.n4759 VCC.n4758 4.5005
R4690 VCC.n4553 VCC.n4549 4.5005
R4691 VCC.n4776 VCC.n4553 4.5005
R4692 VCC.n4789 VCC.n4788 4.5005
R4693 VCC.n4804 VCC.n4803 4.5005
R4694 VCC.n4803 VCC.n4802 4.5005
R4695 VCC.n4819 VCC.n4818 4.5005
R4696 VCC.n4820 VCC.n4819 4.5005
R4697 VCC.n4811 VCC.n4532 4.5005
R4698 VCC.n4822 VCC.n4532 4.5005
R4699 VCC.n4826 VCC.n4524 4.5005
R4700 VCC.n4827 VCC.n4826 4.5005
R4701 VCC.n4847 VCC.n4846 4.5005
R4702 VCC.n4848 VCC.n4847 4.5005
R4703 VCC.n4875 VCC.n4874 4.5005
R4704 VCC.n4513 VCC.n4511 4.5005
R4705 VCC.n4868 VCC.n4513 4.5005
R4706 VCC.n4738 VCC.n4572 4.5005
R4707 VCC.n4737 VCC.n4736 4.5005
R4708 VCC.n4711 VCC.n4583 4.5005
R4709 VCC.n4676 VCC.n4675 4.5005
R4710 VCC.n4641 VCC.n4640 4.5005
R4711 VCC.n4637 VCC.n4634 4.5005
R4712 VCC.n4643 VCC.n4642 4.5005
R4713 VCC.n4644 VCC.n4643 4.5005
R4714 VCC.n4749 VCC.n4748 4.5005
R4715 VCC.n4713 VCC.n4712 4.5005
R4716 VCC.n4636 VCC.n4635 4.5005
R4717 VCC.n4658 VCC.n4611 4.5005
R4718 VCC.n4658 VCC.n4621 4.5005
R4719 VCC.n4673 VCC.n4612 4.5005
R4720 VCC.n4683 VCC.n4682 4.5005
R4721 VCC.n4684 VCC.n4683 4.5005
R4722 VCC.n4688 VCC.n4603 4.5005
R4723 VCC.n4688 VCC.n4592 4.5005
R4724 VCC.n4691 VCC.n4604 4.5005
R4725 VCC.n4699 VCC.n4698 4.5005
R4726 VCC.n4700 VCC.n4699 4.5005
R4727 VCC.n4595 VCC.n4585 4.5005
R4728 VCC.n4596 VCC.n4595 4.5005
R4729 VCC.n4721 VCC.n4720 4.5005
R4730 VCC.n4722 VCC.n4721 4.5005
R4731 VCC.n4740 VCC.n4739 4.5005
R4732 VCC.n4575 VCC.n4573 4.5005
R4733 VCC.n4733 VCC.n4575 4.5005
R4734 VCC.n5289 VCC.n5123 4.5005
R4735 VCC.n5288 VCC.n5287 4.5005
R4736 VCC.n5192 VCC.n5191 4.5005
R4737 VCC.n5188 VCC.n5185 4.5005
R4738 VCC.n5224 VCC.n5163 4.5005
R4739 VCC.n5234 VCC.n5233 4.5005
R4740 VCC.n5235 VCC.n5234 4.5005
R4741 VCC.n5187 VCC.n5186 4.5005
R4742 VCC.n5209 VCC.n5162 4.5005
R4743 VCC.n5209 VCC.n5172 4.5005
R4744 VCC.n5194 VCC.n5193 4.5005
R4745 VCC.n5195 VCC.n5194 4.5005
R4746 VCC.n5239 VCC.n5154 4.5005
R4747 VCC.n5239 VCC.n5143 4.5005
R4748 VCC.n5300 VCC.n5299 4.5005
R4749 VCC.n5264 VCC.n5263 4.5005
R4750 VCC.n5262 VCC.n5134 4.5005
R4751 VCC.n5242 VCC.n5155 4.5005
R4752 VCC.n5250 VCC.n5249 4.5005
R4753 VCC.n5251 VCC.n5250 4.5005
R4754 VCC.n5146 VCC.n5136 4.5005
R4755 VCC.n5147 VCC.n5146 4.5005
R4756 VCC.n5272 VCC.n5271 4.5005
R4757 VCC.n5273 VCC.n5272 4.5005
R4758 VCC.n5291 VCC.n5290 4.5005
R4759 VCC.n5126 VCC.n5124 4.5005
R4760 VCC.n5284 VCC.n5126 4.5005
R4761 VCC.n5227 VCC.n5226 4.5005
R4762 VCC.n5424 VCC.n5062 4.5005
R4763 VCC.n5423 VCC.n5422 4.5005
R4764 VCC.n5317 VCC.n5316 4.5005
R4765 VCC.n5312 VCC.n5309 4.5005
R4766 VCC.n5341 VCC.n5340 4.5005
R4767 VCC.n5311 VCC.n5310 4.5005
R4768 VCC.n5435 VCC.n5434 4.5005
R4769 VCC.n5391 VCC.n5390 4.5005
R4770 VCC.n5389 VCC.n5074 4.5005
R4771 VCC.n5426 VCC.n5425 4.5005
R4772 VCC.n5343 VCC.n5342 4.5005
R4773 VCC.n5356 VCC.n5355 4.5005
R4774 VCC.n5355 VCC.n5354 4.5005
R4775 VCC.n5105 VCC.n5101 4.5005
R4776 VCC.n5328 VCC.n5105 4.5005
R4777 VCC.n5319 VCC.n5318 4.5005
R4778 VCC.n5319 VCC.n5112 4.5005
R4779 VCC.n5371 VCC.n5370 4.5005
R4780 VCC.n5372 VCC.n5371 4.5005
R4781 VCC.n5363 VCC.n5084 4.5005
R4782 VCC.n5374 VCC.n5084 4.5005
R4783 VCC.n5378 VCC.n5076 4.5005
R4784 VCC.n5379 VCC.n5378 4.5005
R4785 VCC.n5399 VCC.n5398 4.5005
R4786 VCC.n5400 VCC.n5399 4.5005
R4787 VCC.n5065 VCC.n5063 4.5005
R4788 VCC.n5419 VCC.n5065 4.5005
R4789 VCC.n5005 VCC.n5000 4.5005
R4790 VCC.n5532 VCC.n5531 4.5005
R4791 VCC.n5442 VCC.n5441 4.5005
R4792 VCC.n5048 VCC.n5046 4.5005
R4793 VCC.n5467 VCC.n5466 4.5005
R4794 VCC.n5034 VCC.n5032 4.5005
R4795 VCC.n5032 VCC.n5031 4.5005
R4796 VCC.n5036 VCC.n5035 4.5005
R4797 VCC.n5450 VCC.n5038 4.5005
R4798 VCC.n5455 VCC.n5454 4.5005
R4799 VCC.n5439 VCC.n5438 4.5005
R4800 VCC.n5444 VCC.n5443 4.5005
R4801 VCC.n5007 VCC.n5006 4.5005
R4802 VCC.n5518 VCC.n5007 4.5005
R4803 VCC.n5506 VCC.n5505 4.5005
R4804 VCC.n5017 VCC.n5004 4.5005
R4805 VCC.n5496 VCC.n5495 4.5005
R4806 VCC.n5026 VCC.n5024 4.5005
R4807 VCC.n5497 VCC.n5019 4.5005
R4808 VCC.n5507 VCC.n5015 4.5005
R4809 VCC.n5509 VCC.n5508 4.5005
R4810 VCC.n5509 VCC.n5013 4.5005
R4811 VCC.n5530 VCC.n4999 4.5005
R4812 VCC.n5541 VCC.n5540 4.5005
R4813 VCC.n5041 VCC.n5039 4.5005
R4814 VCC.n5999 VCC.n5601 4.5005
R4815 VCC.n6002 VCC.n6001 4.5005
R4816 VCC.n6076 VCC.n5556 4.5005
R4817 VCC.n6078 VCC.n6077 4.5005
R4818 VCC.n5573 VCC.n5572 4.5005
R4819 VCC.n5593 VCC.n5591 4.5005
R4820 VCC.n5603 VCC.n5590 4.5005
R4821 VCC.n6032 VCC.n6031 4.5005
R4822 VCC.n6041 VCC.n6040 4.5005
R4823 VCC.n5584 VCC.n5583 4.5005
R4824 VCC.n5564 VCC.n5563 4.5005
R4825 VCC.n6067 VCC.n6066 4.5005
R4826 VCC.n6079 VCC.n5554 4.5005
R4827 VCC.n5568 VCC.n5566 4.5005
R4828 VCC.n6039 VCC.n6038 4.5005
R4829 VCC.n6000 VCC.n5998 4.5005
R4830 VCC.n5996 VCC.n5995 4.5005
R4831 VCC.n6011 VCC.n5602 4.5005
R4832 VCC.n6081 VCC.n6080 4.5005
R4833 VCC.n6081 VCC.n5552 4.5005
R4834 VCC.n5571 VCC.n5569 4.5005
R4835 VCC.n5576 VCC.n5569 4.5005
R4836 VCC.n6027 VCC.n6026 4.5005
R4837 VCC.n6028 VCC.n6027 4.5005
R4838 VCC.n6094 VCC.n6093 4.5005
R4839 VCC.n5981 VCC.n5618 4.5005
R4840 VCC.n5980 VCC.n5979 4.5005
R4841 VCC.n5945 VCC.n5630 4.5005
R4842 VCC.n5899 VCC.n5898 4.5005
R4843 VCC.n5873 VCC.n5872 4.5005
R4844 VCC.n5868 VCC.n5864 4.5005
R4845 VCC.n5874 VCC.n5670 4.5005
R4846 VCC.n5670 VCC.n5668 4.5005
R4847 VCC.n5992 VCC.n5991 4.5005
R4848 VCC.n5947 VCC.n5946 4.5005
R4849 VCC.n5867 VCC.n5866 4.5005
R4850 VCC.n5661 VCC.n5657 4.5005
R4851 VCC.n5884 VCC.n5661 4.5005
R4852 VCC.n5897 VCC.n5896 4.5005
R4853 VCC.n5912 VCC.n5911 4.5005
R4854 VCC.n5911 VCC.n5910 4.5005
R4855 VCC.n5927 VCC.n5926 4.5005
R4856 VCC.n5928 VCC.n5927 4.5005
R4857 VCC.n5919 VCC.n5640 4.5005
R4858 VCC.n5930 VCC.n5640 4.5005
R4859 VCC.n5934 VCC.n5632 4.5005
R4860 VCC.n5935 VCC.n5934 4.5005
R4861 VCC.n5955 VCC.n5954 4.5005
R4862 VCC.n5956 VCC.n5955 4.5005
R4863 VCC.n5983 VCC.n5982 4.5005
R4864 VCC.n5621 VCC.n5619 4.5005
R4865 VCC.n5976 VCC.n5621 4.5005
R4866 VCC.n5846 VCC.n5680 4.5005
R4867 VCC.n5845 VCC.n5844 4.5005
R4868 VCC.n5819 VCC.n5691 4.5005
R4869 VCC.n5784 VCC.n5783 4.5005
R4870 VCC.n5749 VCC.n5748 4.5005
R4871 VCC.n5745 VCC.n5742 4.5005
R4872 VCC.n5751 VCC.n5750 4.5005
R4873 VCC.n5752 VCC.n5751 4.5005
R4874 VCC.n5857 VCC.n5856 4.5005
R4875 VCC.n5821 VCC.n5820 4.5005
R4876 VCC.n5744 VCC.n5743 4.5005
R4877 VCC.n5766 VCC.n5719 4.5005
R4878 VCC.n5766 VCC.n5729 4.5005
R4879 VCC.n5781 VCC.n5720 4.5005
R4880 VCC.n5791 VCC.n5790 4.5005
R4881 VCC.n5792 VCC.n5791 4.5005
R4882 VCC.n5796 VCC.n5711 4.5005
R4883 VCC.n5796 VCC.n5700 4.5005
R4884 VCC.n5799 VCC.n5712 4.5005
R4885 VCC.n5807 VCC.n5806 4.5005
R4886 VCC.n5808 VCC.n5807 4.5005
R4887 VCC.n5703 VCC.n5693 4.5005
R4888 VCC.n5704 VCC.n5703 4.5005
R4889 VCC.n5829 VCC.n5828 4.5005
R4890 VCC.n5830 VCC.n5829 4.5005
R4891 VCC.n5848 VCC.n5847 4.5005
R4892 VCC.n5683 VCC.n5681 4.5005
R4893 VCC.n5841 VCC.n5683 4.5005
R4894 VCC.n6396 VCC.n6230 4.5005
R4895 VCC.n6395 VCC.n6394 4.5005
R4896 VCC.n6299 VCC.n6298 4.5005
R4897 VCC.n6295 VCC.n6292 4.5005
R4898 VCC.n6331 VCC.n6270 4.5005
R4899 VCC.n6341 VCC.n6340 4.5005
R4900 VCC.n6342 VCC.n6341 4.5005
R4901 VCC.n6294 VCC.n6293 4.5005
R4902 VCC.n6316 VCC.n6269 4.5005
R4903 VCC.n6316 VCC.n6279 4.5005
R4904 VCC.n6301 VCC.n6300 4.5005
R4905 VCC.n6302 VCC.n6301 4.5005
R4906 VCC.n6346 VCC.n6261 4.5005
R4907 VCC.n6346 VCC.n6250 4.5005
R4908 VCC.n6407 VCC.n6406 4.5005
R4909 VCC.n6371 VCC.n6370 4.5005
R4910 VCC.n6369 VCC.n6241 4.5005
R4911 VCC.n6349 VCC.n6262 4.5005
R4912 VCC.n6357 VCC.n6356 4.5005
R4913 VCC.n6358 VCC.n6357 4.5005
R4914 VCC.n6253 VCC.n6243 4.5005
R4915 VCC.n6254 VCC.n6253 4.5005
R4916 VCC.n6379 VCC.n6378 4.5005
R4917 VCC.n6380 VCC.n6379 4.5005
R4918 VCC.n6398 VCC.n6397 4.5005
R4919 VCC.n6233 VCC.n6231 4.5005
R4920 VCC.n6391 VCC.n6233 4.5005
R4921 VCC.n6334 VCC.n6333 4.5005
R4922 VCC.n6531 VCC.n6169 4.5005
R4923 VCC.n6530 VCC.n6529 4.5005
R4924 VCC.n6424 VCC.n6423 4.5005
R4925 VCC.n6419 VCC.n6416 4.5005
R4926 VCC.n6448 VCC.n6447 4.5005
R4927 VCC.n6418 VCC.n6417 4.5005
R4928 VCC.n6542 VCC.n6541 4.5005
R4929 VCC.n6498 VCC.n6497 4.5005
R4930 VCC.n6496 VCC.n6181 4.5005
R4931 VCC.n6533 VCC.n6532 4.5005
R4932 VCC.n6450 VCC.n6449 4.5005
R4933 VCC.n6463 VCC.n6462 4.5005
R4934 VCC.n6462 VCC.n6461 4.5005
R4935 VCC.n6212 VCC.n6208 4.5005
R4936 VCC.n6435 VCC.n6212 4.5005
R4937 VCC.n6426 VCC.n6425 4.5005
R4938 VCC.n6426 VCC.n6219 4.5005
R4939 VCC.n6478 VCC.n6477 4.5005
R4940 VCC.n6479 VCC.n6478 4.5005
R4941 VCC.n6470 VCC.n6191 4.5005
R4942 VCC.n6481 VCC.n6191 4.5005
R4943 VCC.n6485 VCC.n6183 4.5005
R4944 VCC.n6486 VCC.n6485 4.5005
R4945 VCC.n6506 VCC.n6505 4.5005
R4946 VCC.n6507 VCC.n6506 4.5005
R4947 VCC.n6172 VCC.n6170 4.5005
R4948 VCC.n6526 VCC.n6172 4.5005
R4949 VCC.n6112 VCC.n6107 4.5005
R4950 VCC.n6639 VCC.n6638 4.5005
R4951 VCC.n6549 VCC.n6548 4.5005
R4952 VCC.n6155 VCC.n6153 4.5005
R4953 VCC.n6574 VCC.n6573 4.5005
R4954 VCC.n6141 VCC.n6139 4.5005
R4955 VCC.n6139 VCC.n6138 4.5005
R4956 VCC.n6143 VCC.n6142 4.5005
R4957 VCC.n6557 VCC.n6145 4.5005
R4958 VCC.n6562 VCC.n6561 4.5005
R4959 VCC.n6546 VCC.n6545 4.5005
R4960 VCC.n6551 VCC.n6550 4.5005
R4961 VCC.n6114 VCC.n6113 4.5005
R4962 VCC.n6625 VCC.n6114 4.5005
R4963 VCC.n6613 VCC.n6612 4.5005
R4964 VCC.n6124 VCC.n6111 4.5005
R4965 VCC.n6603 VCC.n6602 4.5005
R4966 VCC.n6133 VCC.n6131 4.5005
R4967 VCC.n6604 VCC.n6126 4.5005
R4968 VCC.n6614 VCC.n6122 4.5005
R4969 VCC.n6616 VCC.n6615 4.5005
R4970 VCC.n6616 VCC.n6120 4.5005
R4971 VCC.n6637 VCC.n6106 4.5005
R4972 VCC.n6648 VCC.n6647 4.5005
R4973 VCC.n6148 VCC.n6146 4.5005
R4974 VCC.n7106 VCC.n6708 4.5005
R4975 VCC.n7109 VCC.n7108 4.5005
R4976 VCC.n7183 VCC.n6663 4.5005
R4977 VCC.n7185 VCC.n7184 4.5005
R4978 VCC.n6680 VCC.n6679 4.5005
R4979 VCC.n6700 VCC.n6698 4.5005
R4980 VCC.n6710 VCC.n6697 4.5005
R4981 VCC.n7139 VCC.n7138 4.5005
R4982 VCC.n7148 VCC.n7147 4.5005
R4983 VCC.n6691 VCC.n6690 4.5005
R4984 VCC.n6671 VCC.n6670 4.5005
R4985 VCC.n7174 VCC.n7173 4.5005
R4986 VCC.n7186 VCC.n6661 4.5005
R4987 VCC.n6675 VCC.n6673 4.5005
R4988 VCC.n7146 VCC.n7145 4.5005
R4989 VCC.n7107 VCC.n7105 4.5005
R4990 VCC.n7103 VCC.n7102 4.5005
R4991 VCC.n7118 VCC.n6709 4.5005
R4992 VCC.n7188 VCC.n7187 4.5005
R4993 VCC.n7188 VCC.n6659 4.5005
R4994 VCC.n6678 VCC.n6676 4.5005
R4995 VCC.n6683 VCC.n6676 4.5005
R4996 VCC.n7134 VCC.n7133 4.5005
R4997 VCC.n7135 VCC.n7134 4.5005
R4998 VCC.n7201 VCC.n7200 4.5005
R4999 VCC.n7088 VCC.n6725 4.5005
R5000 VCC.n7087 VCC.n7086 4.5005
R5001 VCC.n7052 VCC.n6737 4.5005
R5002 VCC.n7006 VCC.n7005 4.5005
R5003 VCC.n6980 VCC.n6979 4.5005
R5004 VCC.n6975 VCC.n6971 4.5005
R5005 VCC.n6981 VCC.n6777 4.5005
R5006 VCC.n6777 VCC.n6775 4.5005
R5007 VCC.n7099 VCC.n7098 4.5005
R5008 VCC.n7054 VCC.n7053 4.5005
R5009 VCC.n6974 VCC.n6973 4.5005
R5010 VCC.n6768 VCC.n6764 4.5005
R5011 VCC.n6991 VCC.n6768 4.5005
R5012 VCC.n7004 VCC.n7003 4.5005
R5013 VCC.n7019 VCC.n7018 4.5005
R5014 VCC.n7018 VCC.n7017 4.5005
R5015 VCC.n7034 VCC.n7033 4.5005
R5016 VCC.n7035 VCC.n7034 4.5005
R5017 VCC.n7026 VCC.n6747 4.5005
R5018 VCC.n7037 VCC.n6747 4.5005
R5019 VCC.n7041 VCC.n6739 4.5005
R5020 VCC.n7042 VCC.n7041 4.5005
R5021 VCC.n7062 VCC.n7061 4.5005
R5022 VCC.n7063 VCC.n7062 4.5005
R5023 VCC.n7090 VCC.n7089 4.5005
R5024 VCC.n6728 VCC.n6726 4.5005
R5025 VCC.n7083 VCC.n6728 4.5005
R5026 VCC.n6953 VCC.n6787 4.5005
R5027 VCC.n6952 VCC.n6951 4.5005
R5028 VCC.n6926 VCC.n6798 4.5005
R5029 VCC.n6891 VCC.n6890 4.5005
R5030 VCC.n6856 VCC.n6855 4.5005
R5031 VCC.n6852 VCC.n6849 4.5005
R5032 VCC.n6858 VCC.n6857 4.5005
R5033 VCC.n6859 VCC.n6858 4.5005
R5034 VCC.n6964 VCC.n6963 4.5005
R5035 VCC.n6928 VCC.n6927 4.5005
R5036 VCC.n6851 VCC.n6850 4.5005
R5037 VCC.n6873 VCC.n6826 4.5005
R5038 VCC.n6873 VCC.n6836 4.5005
R5039 VCC.n6888 VCC.n6827 4.5005
R5040 VCC.n6898 VCC.n6897 4.5005
R5041 VCC.n6899 VCC.n6898 4.5005
R5042 VCC.n6903 VCC.n6818 4.5005
R5043 VCC.n6903 VCC.n6807 4.5005
R5044 VCC.n6906 VCC.n6819 4.5005
R5045 VCC.n6914 VCC.n6913 4.5005
R5046 VCC.n6915 VCC.n6914 4.5005
R5047 VCC.n6810 VCC.n6800 4.5005
R5048 VCC.n6811 VCC.n6810 4.5005
R5049 VCC.n6936 VCC.n6935 4.5005
R5050 VCC.n6937 VCC.n6936 4.5005
R5051 VCC.n6955 VCC.n6954 4.5005
R5052 VCC.n6790 VCC.n6788 4.5005
R5053 VCC.n6948 VCC.n6790 4.5005
R5054 VCC.n7503 VCC.n7337 4.5005
R5055 VCC.n7502 VCC.n7501 4.5005
R5056 VCC.n7406 VCC.n7405 4.5005
R5057 VCC.n7402 VCC.n7399 4.5005
R5058 VCC.n7438 VCC.n7377 4.5005
R5059 VCC.n7448 VCC.n7447 4.5005
R5060 VCC.n7449 VCC.n7448 4.5005
R5061 VCC.n7401 VCC.n7400 4.5005
R5062 VCC.n7423 VCC.n7376 4.5005
R5063 VCC.n7423 VCC.n7386 4.5005
R5064 VCC.n7408 VCC.n7407 4.5005
R5065 VCC.n7409 VCC.n7408 4.5005
R5066 VCC.n7453 VCC.n7368 4.5005
R5067 VCC.n7453 VCC.n7357 4.5005
R5068 VCC.n7514 VCC.n7513 4.5005
R5069 VCC.n7478 VCC.n7477 4.5005
R5070 VCC.n7476 VCC.n7348 4.5005
R5071 VCC.n7456 VCC.n7369 4.5005
R5072 VCC.n7464 VCC.n7463 4.5005
R5073 VCC.n7465 VCC.n7464 4.5005
R5074 VCC.n7360 VCC.n7350 4.5005
R5075 VCC.n7361 VCC.n7360 4.5005
R5076 VCC.n7486 VCC.n7485 4.5005
R5077 VCC.n7487 VCC.n7486 4.5005
R5078 VCC.n7505 VCC.n7504 4.5005
R5079 VCC.n7340 VCC.n7338 4.5005
R5080 VCC.n7498 VCC.n7340 4.5005
R5081 VCC.n7441 VCC.n7440 4.5005
R5082 VCC.n7638 VCC.n7276 4.5005
R5083 VCC.n7637 VCC.n7636 4.5005
R5084 VCC.n7531 VCC.n7530 4.5005
R5085 VCC.n7526 VCC.n7523 4.5005
R5086 VCC.n7555 VCC.n7554 4.5005
R5087 VCC.n7525 VCC.n7524 4.5005
R5088 VCC.n7649 VCC.n7648 4.5005
R5089 VCC.n7605 VCC.n7604 4.5005
R5090 VCC.n7603 VCC.n7288 4.5005
R5091 VCC.n7640 VCC.n7639 4.5005
R5092 VCC.n7557 VCC.n7556 4.5005
R5093 VCC.n7570 VCC.n7569 4.5005
R5094 VCC.n7569 VCC.n7568 4.5005
R5095 VCC.n7319 VCC.n7315 4.5005
R5096 VCC.n7542 VCC.n7319 4.5005
R5097 VCC.n7533 VCC.n7532 4.5005
R5098 VCC.n7533 VCC.n7326 4.5005
R5099 VCC.n7585 VCC.n7584 4.5005
R5100 VCC.n7586 VCC.n7585 4.5005
R5101 VCC.n7577 VCC.n7298 4.5005
R5102 VCC.n7588 VCC.n7298 4.5005
R5103 VCC.n7592 VCC.n7290 4.5005
R5104 VCC.n7593 VCC.n7592 4.5005
R5105 VCC.n7613 VCC.n7612 4.5005
R5106 VCC.n7614 VCC.n7613 4.5005
R5107 VCC.n7279 VCC.n7277 4.5005
R5108 VCC.n7633 VCC.n7279 4.5005
R5109 VCC.n7219 VCC.n7214 4.5005
R5110 VCC.n7746 VCC.n7745 4.5005
R5111 VCC.n7656 VCC.n7655 4.5005
R5112 VCC.n7262 VCC.n7260 4.5005
R5113 VCC.n7681 VCC.n7680 4.5005
R5114 VCC.n7248 VCC.n7246 4.5005
R5115 VCC.n7246 VCC.n7245 4.5005
R5116 VCC.n7250 VCC.n7249 4.5005
R5117 VCC.n7664 VCC.n7252 4.5005
R5118 VCC.n7669 VCC.n7668 4.5005
R5119 VCC.n7653 VCC.n7652 4.5005
R5120 VCC.n7658 VCC.n7657 4.5005
R5121 VCC.n7221 VCC.n7220 4.5005
R5122 VCC.n7732 VCC.n7221 4.5005
R5123 VCC.n7720 VCC.n7719 4.5005
R5124 VCC.n7231 VCC.n7218 4.5005
R5125 VCC.n7710 VCC.n7709 4.5005
R5126 VCC.n7240 VCC.n7238 4.5005
R5127 VCC.n7711 VCC.n7233 4.5005
R5128 VCC.n7721 VCC.n7229 4.5005
R5129 VCC.n7723 VCC.n7722 4.5005
R5130 VCC.n7723 VCC.n7227 4.5005
R5131 VCC.n7744 VCC.n7213 4.5005
R5132 VCC.n7755 VCC.n7754 4.5005
R5133 VCC.n7255 VCC.n7253 4.5005
R5134 VCC.n8213 VCC.n7815 4.5005
R5135 VCC.n8216 VCC.n8215 4.5005
R5136 VCC.n8290 VCC.n7770 4.5005
R5137 VCC.n8292 VCC.n8291 4.5005
R5138 VCC.n7787 VCC.n7786 4.5005
R5139 VCC.n7807 VCC.n7805 4.5005
R5140 VCC.n7817 VCC.n7804 4.5005
R5141 VCC.n8246 VCC.n8245 4.5005
R5142 VCC.n8255 VCC.n8254 4.5005
R5143 VCC.n7798 VCC.n7797 4.5005
R5144 VCC.n7778 VCC.n7777 4.5005
R5145 VCC.n8281 VCC.n8280 4.5005
R5146 VCC.n8293 VCC.n7768 4.5005
R5147 VCC.n7782 VCC.n7780 4.5005
R5148 VCC.n8253 VCC.n8252 4.5005
R5149 VCC.n8214 VCC.n8212 4.5005
R5150 VCC.n8210 VCC.n8209 4.5005
R5151 VCC.n8225 VCC.n7816 4.5005
R5152 VCC.n8295 VCC.n8294 4.5005
R5153 VCC.n8295 VCC.n7766 4.5005
R5154 VCC.n7785 VCC.n7783 4.5005
R5155 VCC.n7790 VCC.n7783 4.5005
R5156 VCC.n8241 VCC.n8240 4.5005
R5157 VCC.n8242 VCC.n8241 4.5005
R5158 VCC.n8308 VCC.n8307 4.5005
R5159 VCC.n8195 VCC.n7832 4.5005
R5160 VCC.n8194 VCC.n8193 4.5005
R5161 VCC.n8159 VCC.n7844 4.5005
R5162 VCC.n8113 VCC.n8112 4.5005
R5163 VCC.n8087 VCC.n8086 4.5005
R5164 VCC.n8082 VCC.n8078 4.5005
R5165 VCC.n8088 VCC.n7884 4.5005
R5166 VCC.n7884 VCC.n7882 4.5005
R5167 VCC.n8206 VCC.n8205 4.5005
R5168 VCC.n8161 VCC.n8160 4.5005
R5169 VCC.n8081 VCC.n8080 4.5005
R5170 VCC.n7875 VCC.n7871 4.5005
R5171 VCC.n8098 VCC.n7875 4.5005
R5172 VCC.n8111 VCC.n8110 4.5005
R5173 VCC.n8126 VCC.n8125 4.5005
R5174 VCC.n8125 VCC.n8124 4.5005
R5175 VCC.n8141 VCC.n8140 4.5005
R5176 VCC.n8142 VCC.n8141 4.5005
R5177 VCC.n8133 VCC.n7854 4.5005
R5178 VCC.n8144 VCC.n7854 4.5005
R5179 VCC.n8148 VCC.n7846 4.5005
R5180 VCC.n8149 VCC.n8148 4.5005
R5181 VCC.n8169 VCC.n8168 4.5005
R5182 VCC.n8170 VCC.n8169 4.5005
R5183 VCC.n8197 VCC.n8196 4.5005
R5184 VCC.n7835 VCC.n7833 4.5005
R5185 VCC.n8190 VCC.n7835 4.5005
R5186 VCC.n8060 VCC.n7894 4.5005
R5187 VCC.n8059 VCC.n8058 4.5005
R5188 VCC.n8033 VCC.n7905 4.5005
R5189 VCC.n7998 VCC.n7997 4.5005
R5190 VCC.n7963 VCC.n7962 4.5005
R5191 VCC.n7959 VCC.n7956 4.5005
R5192 VCC.n7965 VCC.n7964 4.5005
R5193 VCC.n7966 VCC.n7965 4.5005
R5194 VCC.n8071 VCC.n8070 4.5005
R5195 VCC.n8035 VCC.n8034 4.5005
R5196 VCC.n7958 VCC.n7957 4.5005
R5197 VCC.n7980 VCC.n7933 4.5005
R5198 VCC.n7980 VCC.n7943 4.5005
R5199 VCC.n7995 VCC.n7934 4.5005
R5200 VCC.n8005 VCC.n8004 4.5005
R5201 VCC.n8006 VCC.n8005 4.5005
R5202 VCC.n8010 VCC.n7925 4.5005
R5203 VCC.n8010 VCC.n7914 4.5005
R5204 VCC.n8013 VCC.n7926 4.5005
R5205 VCC.n8021 VCC.n8020 4.5005
R5206 VCC.n8022 VCC.n8021 4.5005
R5207 VCC.n7917 VCC.n7907 4.5005
R5208 VCC.n7918 VCC.n7917 4.5005
R5209 VCC.n8043 VCC.n8042 4.5005
R5210 VCC.n8044 VCC.n8043 4.5005
R5211 VCC.n8062 VCC.n8061 4.5005
R5212 VCC.n7897 VCC.n7895 4.5005
R5213 VCC.n8055 VCC.n7897 4.5005
R5214 VCC.n8558 VCC.n8383 4.5005
R5215 VCC.n8557 VCC.n8556 4.5005
R5216 VCC.n8451 VCC.n8450 4.5005
R5217 VCC.n8446 VCC.n8443 4.5005
R5218 VCC.n8475 VCC.n8474 4.5005
R5219 VCC.n8445 VCC.n8444 4.5005
R5220 VCC.n8569 VCC.n8568 4.5005
R5221 VCC.n8525 VCC.n8524 4.5005
R5222 VCC.n8523 VCC.n8395 4.5005
R5223 VCC.n8560 VCC.n8559 4.5005
R5224 VCC.n8477 VCC.n8476 4.5005
R5225 VCC.n8490 VCC.n8489 4.5005
R5226 VCC.n8489 VCC.n8488 4.5005
R5227 VCC.n8426 VCC.n8422 4.5005
R5228 VCC.n8462 VCC.n8426 4.5005
R5229 VCC.n8453 VCC.n8452 4.5005
R5230 VCC.n8453 VCC.n8433 4.5005
R5231 VCC.n8505 VCC.n8504 4.5005
R5232 VCC.n8506 VCC.n8505 4.5005
R5233 VCC.n8497 VCC.n8405 4.5005
R5234 VCC.n8508 VCC.n8405 4.5005
R5235 VCC.n8512 VCC.n8397 4.5005
R5236 VCC.n8513 VCC.n8512 4.5005
R5237 VCC.n8533 VCC.n8532 4.5005
R5238 VCC.n8534 VCC.n8533 4.5005
R5239 VCC.n8386 VCC.n8384 4.5005
R5240 VCC.n8553 VCC.n8386 4.5005
R5241 VCC.n8326 VCC.n8321 4.5005
R5242 VCC.n8666 VCC.n8665 4.5005
R5243 VCC.n8576 VCC.n8575 4.5005
R5244 VCC.n8369 VCC.n8367 4.5005
R5245 VCC.n8601 VCC.n8600 4.5005
R5246 VCC.n8355 VCC.n8353 4.5005
R5247 VCC.n8353 VCC.n8352 4.5005
R5248 VCC.n8357 VCC.n8356 4.5005
R5249 VCC.n8584 VCC.n8359 4.5005
R5250 VCC.n8589 VCC.n8588 4.5005
R5251 VCC.n8573 VCC.n8572 4.5005
R5252 VCC.n8578 VCC.n8577 4.5005
R5253 VCC.n8328 VCC.n8327 4.5005
R5254 VCC.n8652 VCC.n8328 4.5005
R5255 VCC.n8640 VCC.n8639 4.5005
R5256 VCC.n8338 VCC.n8325 4.5005
R5257 VCC.n8630 VCC.n8629 4.5005
R5258 VCC.n8347 VCC.n8345 4.5005
R5259 VCC.n8631 VCC.n8340 4.5005
R5260 VCC.n8641 VCC.n8336 4.5005
R5261 VCC.n8643 VCC.n8642 4.5005
R5262 VCC.n8643 VCC.n8334 4.5005
R5263 VCC.n8664 VCC.n8320 4.5005
R5264 VCC.n8675 VCC.n8674 4.5005
R5265 VCC.n8362 VCC.n8360 4.5005
R5266 VCC.n548 VCC.n4 4.31039
R5267 VCC.n1102 VCC.n558 4.31039
R5268 VCC.n1655 VCC.n1111 4.31039
R5269 VCC.n2211 VCC.n1667 4.31039
R5270 VCC.n2764 VCC.n2220 4.31039
R5271 VCC.n3320 VCC.n2776 4.31039
R5272 VCC.n3873 VCC.n3329 4.31039
R5273 VCC.n4429 VCC.n3885 4.31039
R5274 VCC.n4982 VCC.n4438 4.31039
R5275 VCC.n5538 VCC.n4994 4.31039
R5276 VCC.n6090 VCC.n5546 4.31039
R5277 VCC.n6645 VCC.n6101 4.31039
R5278 VCC.n7197 VCC.n6653 4.31039
R5279 VCC.n7752 VCC.n7208 4.31039
R5280 VCC.n8304 VCC.n7760 4.31039
R5281 VCC.n8672 VCC.n8315 4.31039
R5282 VCC.n472 VCC.n41 3.51902
R5283 VCC.n525 VCC.n22 3.51902
R5284 VCC.n1024 VCC.n593 3.51902
R5285 VCC.n1077 VCC.n574 3.51902
R5286 VCC.n1585 VCC.n1584 3.51902
R5287 VCC.n1621 VCC.n1620 3.51902
R5288 VCC.n2133 VCC.n1702 3.51902
R5289 VCC.n2186 VCC.n1683 3.51902
R5290 VCC.n2694 VCC.n2693 3.51902
R5291 VCC.n2730 VCC.n2729 3.51902
R5292 VCC.n3242 VCC.n2811 3.51902
R5293 VCC.n3295 VCC.n2792 3.51902
R5294 VCC.n3803 VCC.n3802 3.51902
R5295 VCC.n3839 VCC.n3838 3.51902
R5296 VCC.n4351 VCC.n3920 3.51902
R5297 VCC.n4404 VCC.n3901 3.51902
R5298 VCC.n4912 VCC.n4911 3.51902
R5299 VCC.n4948 VCC.n4947 3.51902
R5300 VCC.n5460 VCC.n5029 3.51902
R5301 VCC.n5513 VCC.n5010 3.51902
R5302 VCC.n6020 VCC.n6019 3.51902
R5303 VCC.n6056 VCC.n6055 3.51902
R5304 VCC.n6567 VCC.n6136 3.51902
R5305 VCC.n6620 VCC.n6117 3.51902
R5306 VCC.n7127 VCC.n7126 3.51902
R5307 VCC.n7163 VCC.n7162 3.51902
R5308 VCC.n7674 VCC.n7243 3.51902
R5309 VCC.n7727 VCC.n7224 3.51902
R5310 VCC.n8234 VCC.n8233 3.51902
R5311 VCC.n8270 VCC.n8269 3.51902
R5312 VCC.n8594 VCC.n8350 3.51902
R5313 VCC.n8647 VCC.n8331 3.51902
R5314 VCC.n313 VCC.n312 3.42479
R5315 VCC.n315 VCC.n314 3.42479
R5316 VCC.n865 VCC.n864 3.42479
R5317 VCC.n867 VCC.n866 3.42479
R5318 VCC.n1425 VCC.n1424 3.42479
R5319 VCC.n1423 VCC.n1422 3.42479
R5320 VCC.n1974 VCC.n1973 3.42479
R5321 VCC.n1976 VCC.n1975 3.42479
R5322 VCC.n2534 VCC.n2533 3.42479
R5323 VCC.n2532 VCC.n2531 3.42479
R5324 VCC.n3083 VCC.n3082 3.42479
R5325 VCC.n3085 VCC.n3084 3.42479
R5326 VCC.n3643 VCC.n3642 3.42479
R5327 VCC.n3641 VCC.n3640 3.42479
R5328 VCC.n4192 VCC.n4191 3.42479
R5329 VCC.n4194 VCC.n4193 3.42479
R5330 VCC.n4752 VCC.n4751 3.42479
R5331 VCC.n4750 VCC.n4749 3.42479
R5332 VCC.n5301 VCC.n5300 3.42479
R5333 VCC.n5303 VCC.n5302 3.42479
R5334 VCC.n5860 VCC.n5859 3.42479
R5335 VCC.n5858 VCC.n5857 3.42479
R5336 VCC.n6408 VCC.n6407 3.42479
R5337 VCC.n6410 VCC.n6409 3.42479
R5338 VCC.n6967 VCC.n6966 3.42479
R5339 VCC.n6965 VCC.n6964 3.42479
R5340 VCC.n7515 VCC.n7514 3.42479
R5341 VCC.n7517 VCC.n7516 3.42479
R5342 VCC.n8074 VCC.n8073 3.42479
R5343 VCC.n8072 VCC.n8071 3.42479
R5344 VCC.n8437 VCC.n8436 3.42479
R5345 VCC.n192 VCC.n191 3.42389
R5346 VCC.n448 VCC.n447 3.42389
R5347 VCC.n450 VCC.n449 3.42389
R5348 VCC.n744 VCC.n743 3.42389
R5349 VCC.n1000 VCC.n999 3.42389
R5350 VCC.n1002 VCC.n1001 3.42389
R5351 VCC.n1560 VCC.n1559 3.42389
R5352 VCC.n1558 VCC.n1557 3.42389
R5353 VCC.n1302 VCC.n1301 3.42389
R5354 VCC.n1853 VCC.n1852 3.42389
R5355 VCC.n2109 VCC.n2108 3.42389
R5356 VCC.n2111 VCC.n2110 3.42389
R5357 VCC.n2669 VCC.n2668 3.42389
R5358 VCC.n2667 VCC.n2666 3.42389
R5359 VCC.n2411 VCC.n2410 3.42389
R5360 VCC.n2962 VCC.n2961 3.42389
R5361 VCC.n3218 VCC.n3217 3.42389
R5362 VCC.n3220 VCC.n3219 3.42389
R5363 VCC.n3778 VCC.n3777 3.42389
R5364 VCC.n3776 VCC.n3775 3.42389
R5365 VCC.n3520 VCC.n3519 3.42389
R5366 VCC.n4071 VCC.n4070 3.42389
R5367 VCC.n4327 VCC.n4326 3.42389
R5368 VCC.n4329 VCC.n4328 3.42389
R5369 VCC.n4887 VCC.n4886 3.42389
R5370 VCC.n4885 VCC.n4884 3.42389
R5371 VCC.n4629 VCC.n4628 3.42389
R5372 VCC.n5180 VCC.n5179 3.42389
R5373 VCC.n5436 VCC.n5435 3.42389
R5374 VCC.n5438 VCC.n5437 3.42389
R5375 VCC.n5995 VCC.n5994 3.42389
R5376 VCC.n5993 VCC.n5992 3.42389
R5377 VCC.n5737 VCC.n5736 3.42389
R5378 VCC.n6287 VCC.n6286 3.42389
R5379 VCC.n6543 VCC.n6542 3.42389
R5380 VCC.n6545 VCC.n6544 3.42389
R5381 VCC.n7102 VCC.n7101 3.42389
R5382 VCC.n7100 VCC.n7099 3.42389
R5383 VCC.n6844 VCC.n6843 3.42389
R5384 VCC.n7394 VCC.n7393 3.42389
R5385 VCC.n7650 VCC.n7649 3.42389
R5386 VCC.n7652 VCC.n7651 3.42389
R5387 VCC.n8209 VCC.n8208 3.42389
R5388 VCC.n8207 VCC.n8206 3.42389
R5389 VCC.n7951 VCC.n7950 3.42389
R5390 VCC.n8570 VCC.n8569 3.42389
R5391 VCC.n8572 VCC.n8571 3.42389
R5392 VCC.n552 VCC.n551 3.423
R5393 VCC.n1106 VCC.n1105 3.423
R5394 VCC.n1660 VCC.n1659 3.423
R5395 VCC.n2215 VCC.n2214 3.423
R5396 VCC.n2769 VCC.n2768 3.423
R5397 VCC.n3324 VCC.n3323 3.423
R5398 VCC.n3878 VCC.n3877 3.423
R5399 VCC.n4433 VCC.n4432 3.423
R5400 VCC.n4987 VCC.n4986 3.423
R5401 VCC.n5542 VCC.n5541 3.423
R5402 VCC.n6095 VCC.n6094 3.423
R5403 VCC.n6649 VCC.n6648 3.423
R5404 VCC.n7202 VCC.n7201 3.423
R5405 VCC.n7756 VCC.n7755 3.423
R5406 VCC.n8309 VCC.n8308 3.423
R5407 VCC.n8676 VCC.n8675 3.423
R5408 VCC.n514 VCC.n513 3.4105
R5409 VCC.n536 VCC.n535 3.4105
R5410 VCC.n535 VCC.n534 3.4105
R5411 VCC.n504 VCC.n33 3.4105
R5412 VCC.n33 VCC.n32 3.4105
R5413 VCC.n506 VCC.n505 3.4105
R5414 VCC.n512 VCC.n511 3.4105
R5415 VCC.n511 VCC.n510 3.4105
R5416 VCC.n486 VCC.n485 3.4105
R5417 VCC.n486 VCC.n45 3.4105
R5418 VCC.n482 VCC.n35 3.4105
R5419 VCC.n503 VCC.n502 3.4105
R5420 VCC.n502 VCC.n501 3.4105
R5421 VCC.n464 VCC.n461 3.4105
R5422 VCC.n464 VCC.n463 3.4105
R5423 VCC.n481 VCC.n480 3.4105
R5424 VCC.n444 VCC.n443 3.4105
R5425 VCC.n445 VCC.n444 3.4105
R5426 VCC.n409 VCC.n408 3.4105
R5427 VCC.n442 VCC.n441 3.4105
R5428 VCC.n441 VCC.n440 3.4105
R5429 VCC.n379 VCC.n378 3.4105
R5430 VCC.n378 VCC.n377 3.4105
R5431 VCC.n374 VCC.n372 3.4105
R5432 VCC.n407 VCC.n406 3.4105
R5433 VCC.n406 VCC.n405 3.4105
R5434 VCC.n103 VCC.n102 3.4105
R5435 VCC.n350 VCC.n103 3.4105
R5436 VCC.n371 VCC.n100 3.4105
R5437 VCC.n381 VCC.n380 3.4105
R5438 VCC.n381 VCC.n99 3.4105
R5439 VCC.n344 VCC.n114 3.4105
R5440 VCC.n344 VCC.n343 3.4105
R5441 VCC.n348 VCC.n347 3.4105
R5442 VCC.n318 VCC.n317 3.4105
R5443 VCC.n318 VCC.n125 3.4105
R5444 VCC.n309 VCC.n308 3.4105
R5445 VCC.n310 VCC.n309 3.4105
R5446 VCC.n282 VCC.n281 3.4105
R5447 VCC.n307 VCC.n306 3.4105
R5448 VCC.n306 VCC.n305 3.4105
R5449 VCC.n258 VCC.n163 3.4105
R5450 VCC.n163 VCC.n157 3.4105
R5451 VCC.n260 VCC.n259 3.4105
R5452 VCC.n280 VCC.n279 3.4105
R5453 VCC.n279 VCC.n278 3.4105
R5454 VCC.n242 VCC.n171 3.4105
R5455 VCC.n171 VCC.n170 3.4105
R5456 VCC.n172 VCC.n165 3.4105
R5457 VCC.n257 VCC.n256 3.4105
R5458 VCC.n256 VCC.n255 3.4105
R5459 VCC.n219 VCC.n218 3.4105
R5460 VCC.n220 VCC.n219 3.4105
R5461 VCC.n241 VCC.n240 3.4105
R5462 VCC.n217 VCC.n216 3.4105
R5463 VCC.n216 VCC.n215 3.4105
R5464 VCC.n460 VCC.n459 3.4105
R5465 VCC.n459 VCC.n458 3.4105
R5466 VCC.n538 VCC.n537 3.4105
R5467 VCC.n538 VCC.n2 3.4105
R5468 VCC.n1090 VCC.n1089 3.4105
R5469 VCC.n1090 VCC.n556 3.4105
R5470 VCC.n1066 VCC.n1065 3.4105
R5471 VCC.n1088 VCC.n1087 3.4105
R5472 VCC.n1087 VCC.n1086 3.4105
R5473 VCC.n1056 VCC.n585 3.4105
R5474 VCC.n585 VCC.n584 3.4105
R5475 VCC.n1058 VCC.n1057 3.4105
R5476 VCC.n1064 VCC.n1063 3.4105
R5477 VCC.n1063 VCC.n1062 3.4105
R5478 VCC.n1038 VCC.n1037 3.4105
R5479 VCC.n1038 VCC.n597 3.4105
R5480 VCC.n1034 VCC.n587 3.4105
R5481 VCC.n1055 VCC.n1054 3.4105
R5482 VCC.n1054 VCC.n1053 3.4105
R5483 VCC.n1016 VCC.n1013 3.4105
R5484 VCC.n1016 VCC.n1015 3.4105
R5485 VCC.n1033 VCC.n1032 3.4105
R5486 VCC.n1012 VCC.n1011 3.4105
R5487 VCC.n1011 VCC.n1010 3.4105
R5488 VCC.n996 VCC.n995 3.4105
R5489 VCC.n997 VCC.n996 3.4105
R5490 VCC.n961 VCC.n960 3.4105
R5491 VCC.n994 VCC.n993 3.4105
R5492 VCC.n993 VCC.n992 3.4105
R5493 VCC.n931 VCC.n930 3.4105
R5494 VCC.n930 VCC.n929 3.4105
R5495 VCC.n926 VCC.n924 3.4105
R5496 VCC.n959 VCC.n958 3.4105
R5497 VCC.n958 VCC.n957 3.4105
R5498 VCC.n655 VCC.n654 3.4105
R5499 VCC.n902 VCC.n655 3.4105
R5500 VCC.n923 VCC.n652 3.4105
R5501 VCC.n933 VCC.n932 3.4105
R5502 VCC.n933 VCC.n651 3.4105
R5503 VCC.n896 VCC.n666 3.4105
R5504 VCC.n896 VCC.n895 3.4105
R5505 VCC.n900 VCC.n899 3.4105
R5506 VCC.n870 VCC.n869 3.4105
R5507 VCC.n870 VCC.n677 3.4105
R5508 VCC.n861 VCC.n860 3.4105
R5509 VCC.n862 VCC.n861 3.4105
R5510 VCC.n834 VCC.n833 3.4105
R5511 VCC.n859 VCC.n858 3.4105
R5512 VCC.n858 VCC.n857 3.4105
R5513 VCC.n810 VCC.n715 3.4105
R5514 VCC.n715 VCC.n709 3.4105
R5515 VCC.n812 VCC.n811 3.4105
R5516 VCC.n832 VCC.n831 3.4105
R5517 VCC.n831 VCC.n830 3.4105
R5518 VCC.n794 VCC.n723 3.4105
R5519 VCC.n723 VCC.n722 3.4105
R5520 VCC.n724 VCC.n717 3.4105
R5521 VCC.n809 VCC.n808 3.4105
R5522 VCC.n808 VCC.n807 3.4105
R5523 VCC.n771 VCC.n770 3.4105
R5524 VCC.n772 VCC.n771 3.4105
R5525 VCC.n793 VCC.n792 3.4105
R5526 VCC.n769 VCC.n768 3.4105
R5527 VCC.n768 VCC.n767 3.4105
R5528 VCC.n1419 VCC.n1418 3.4105
R5529 VCC.n1420 VCC.n1419 3.4105
R5530 VCC.n1392 VCC.n1391 3.4105
R5531 VCC.n1417 VCC.n1416 3.4105
R5532 VCC.n1416 VCC.n1415 3.4105
R5533 VCC.n1368 VCC.n1273 3.4105
R5534 VCC.n1273 VCC.n1267 3.4105
R5535 VCC.n1370 VCC.n1369 3.4105
R5536 VCC.n1390 VCC.n1389 3.4105
R5537 VCC.n1389 VCC.n1388 3.4105
R5538 VCC.n1352 VCC.n1281 3.4105
R5539 VCC.n1281 VCC.n1280 3.4105
R5540 VCC.n1282 VCC.n1275 3.4105
R5541 VCC.n1367 VCC.n1366 3.4105
R5542 VCC.n1366 VCC.n1365 3.4105
R5543 VCC.n1329 VCC.n1328 3.4105
R5544 VCC.n1330 VCC.n1329 3.4105
R5545 VCC.n1351 VCC.n1350 3.4105
R5546 VCC.n1327 VCC.n1326 3.4105
R5547 VCC.n1326 VCC.n1325 3.4105
R5548 VCC.n1571 VCC.n1570 3.4105
R5549 VCC.n1570 VCC.n1569 3.4105
R5550 VCC.n1630 VCC.n1629 3.4105
R5551 VCC.n1635 VCC.n1634 3.4105
R5552 VCC.n1634 VCC.n1633 3.4105
R5553 VCC.n1613 VCC.n1612 3.4105
R5554 VCC.n1614 VCC.n1613 3.4105
R5555 VCC.n1611 VCC.n1610 3.4105
R5556 VCC.n1628 VCC.n1627 3.4105
R5557 VCC.n1627 VCC.n1626 3.4105
R5558 VCC.n1600 VCC.n1153 3.4105
R5559 VCC.n1153 VCC.n1152 3.4105
R5560 VCC.n1151 VCC.n1150 3.4105
R5561 VCC.n1608 VCC.n1607 3.4105
R5562 VCC.n1607 VCC.n1146 3.4105
R5563 VCC.n1573 VCC.n1572 3.4105
R5564 VCC.n1573 VCC.n1169 3.4105
R5565 VCC.n1599 VCC.n1598 3.4105
R5566 VCC.n1637 VCC.n1636 3.4105
R5567 VCC.n1637 VCC.n1110 3.4105
R5568 VCC.n1554 VCC.n1553 3.4105
R5569 VCC.n1555 VCC.n1554 3.4105
R5570 VCC.n1518 VCC.n1517 3.4105
R5571 VCC.n1552 VCC.n1551 3.4105
R5572 VCC.n1551 VCC.n1550 3.4105
R5573 VCC.n1488 VCC.n1487 3.4105
R5574 VCC.n1487 VCC.n1486 3.4105
R5575 VCC.n1483 VCC.n1481 3.4105
R5576 VCC.n1516 VCC.n1515 3.4105
R5577 VCC.n1515 VCC.n1514 3.4105
R5578 VCC.n1212 VCC.n1211 3.4105
R5579 VCC.n1459 VCC.n1212 3.4105
R5580 VCC.n1480 VCC.n1209 3.4105
R5581 VCC.n1490 VCC.n1489 3.4105
R5582 VCC.n1490 VCC.n1208 3.4105
R5583 VCC.n1453 VCC.n1223 3.4105
R5584 VCC.n1453 VCC.n1452 3.4105
R5585 VCC.n1457 VCC.n1456 3.4105
R5586 VCC.n1428 VCC.n1427 3.4105
R5587 VCC.n1428 VCC.n1234 3.4105
R5588 VCC.n2199 VCC.n2198 3.4105
R5589 VCC.n2199 VCC.n1665 3.4105
R5590 VCC.n2175 VCC.n2174 3.4105
R5591 VCC.n2197 VCC.n2196 3.4105
R5592 VCC.n2196 VCC.n2195 3.4105
R5593 VCC.n2165 VCC.n1694 3.4105
R5594 VCC.n1694 VCC.n1693 3.4105
R5595 VCC.n2167 VCC.n2166 3.4105
R5596 VCC.n2173 VCC.n2172 3.4105
R5597 VCC.n2172 VCC.n2171 3.4105
R5598 VCC.n2147 VCC.n2146 3.4105
R5599 VCC.n2147 VCC.n1706 3.4105
R5600 VCC.n2143 VCC.n1696 3.4105
R5601 VCC.n2164 VCC.n2163 3.4105
R5602 VCC.n2163 VCC.n2162 3.4105
R5603 VCC.n2125 VCC.n2122 3.4105
R5604 VCC.n2125 VCC.n2124 3.4105
R5605 VCC.n2142 VCC.n2141 3.4105
R5606 VCC.n2121 VCC.n2120 3.4105
R5607 VCC.n2120 VCC.n2119 3.4105
R5608 VCC.n2105 VCC.n2104 3.4105
R5609 VCC.n2106 VCC.n2105 3.4105
R5610 VCC.n2070 VCC.n2069 3.4105
R5611 VCC.n2103 VCC.n2102 3.4105
R5612 VCC.n2102 VCC.n2101 3.4105
R5613 VCC.n2040 VCC.n2039 3.4105
R5614 VCC.n2039 VCC.n2038 3.4105
R5615 VCC.n2035 VCC.n2033 3.4105
R5616 VCC.n2068 VCC.n2067 3.4105
R5617 VCC.n2067 VCC.n2066 3.4105
R5618 VCC.n1764 VCC.n1763 3.4105
R5619 VCC.n2011 VCC.n1764 3.4105
R5620 VCC.n2032 VCC.n1761 3.4105
R5621 VCC.n2042 VCC.n2041 3.4105
R5622 VCC.n2042 VCC.n1760 3.4105
R5623 VCC.n2005 VCC.n1775 3.4105
R5624 VCC.n2005 VCC.n2004 3.4105
R5625 VCC.n2009 VCC.n2008 3.4105
R5626 VCC.n1979 VCC.n1978 3.4105
R5627 VCC.n1979 VCC.n1786 3.4105
R5628 VCC.n1970 VCC.n1969 3.4105
R5629 VCC.n1971 VCC.n1970 3.4105
R5630 VCC.n1943 VCC.n1942 3.4105
R5631 VCC.n1968 VCC.n1967 3.4105
R5632 VCC.n1967 VCC.n1966 3.4105
R5633 VCC.n1919 VCC.n1824 3.4105
R5634 VCC.n1824 VCC.n1818 3.4105
R5635 VCC.n1921 VCC.n1920 3.4105
R5636 VCC.n1941 VCC.n1940 3.4105
R5637 VCC.n1940 VCC.n1939 3.4105
R5638 VCC.n1903 VCC.n1832 3.4105
R5639 VCC.n1832 VCC.n1831 3.4105
R5640 VCC.n1833 VCC.n1826 3.4105
R5641 VCC.n1918 VCC.n1917 3.4105
R5642 VCC.n1917 VCC.n1916 3.4105
R5643 VCC.n1880 VCC.n1879 3.4105
R5644 VCC.n1881 VCC.n1880 3.4105
R5645 VCC.n1902 VCC.n1901 3.4105
R5646 VCC.n1878 VCC.n1877 3.4105
R5647 VCC.n1877 VCC.n1876 3.4105
R5648 VCC.n2528 VCC.n2527 3.4105
R5649 VCC.n2529 VCC.n2528 3.4105
R5650 VCC.n2501 VCC.n2500 3.4105
R5651 VCC.n2526 VCC.n2525 3.4105
R5652 VCC.n2525 VCC.n2524 3.4105
R5653 VCC.n2477 VCC.n2382 3.4105
R5654 VCC.n2382 VCC.n2376 3.4105
R5655 VCC.n2479 VCC.n2478 3.4105
R5656 VCC.n2499 VCC.n2498 3.4105
R5657 VCC.n2498 VCC.n2497 3.4105
R5658 VCC.n2461 VCC.n2390 3.4105
R5659 VCC.n2390 VCC.n2389 3.4105
R5660 VCC.n2391 VCC.n2384 3.4105
R5661 VCC.n2476 VCC.n2475 3.4105
R5662 VCC.n2475 VCC.n2474 3.4105
R5663 VCC.n2438 VCC.n2437 3.4105
R5664 VCC.n2439 VCC.n2438 3.4105
R5665 VCC.n2460 VCC.n2459 3.4105
R5666 VCC.n2436 VCC.n2435 3.4105
R5667 VCC.n2435 VCC.n2434 3.4105
R5668 VCC.n2680 VCC.n2679 3.4105
R5669 VCC.n2679 VCC.n2678 3.4105
R5670 VCC.n2739 VCC.n2738 3.4105
R5671 VCC.n2744 VCC.n2743 3.4105
R5672 VCC.n2743 VCC.n2742 3.4105
R5673 VCC.n2722 VCC.n2721 3.4105
R5674 VCC.n2723 VCC.n2722 3.4105
R5675 VCC.n2720 VCC.n2719 3.4105
R5676 VCC.n2737 VCC.n2736 3.4105
R5677 VCC.n2736 VCC.n2735 3.4105
R5678 VCC.n2709 VCC.n2262 3.4105
R5679 VCC.n2262 VCC.n2261 3.4105
R5680 VCC.n2260 VCC.n2259 3.4105
R5681 VCC.n2717 VCC.n2716 3.4105
R5682 VCC.n2716 VCC.n2255 3.4105
R5683 VCC.n2682 VCC.n2681 3.4105
R5684 VCC.n2682 VCC.n2278 3.4105
R5685 VCC.n2708 VCC.n2707 3.4105
R5686 VCC.n2746 VCC.n2745 3.4105
R5687 VCC.n2746 VCC.n2219 3.4105
R5688 VCC.n2663 VCC.n2662 3.4105
R5689 VCC.n2664 VCC.n2663 3.4105
R5690 VCC.n2627 VCC.n2626 3.4105
R5691 VCC.n2661 VCC.n2660 3.4105
R5692 VCC.n2660 VCC.n2659 3.4105
R5693 VCC.n2597 VCC.n2596 3.4105
R5694 VCC.n2596 VCC.n2595 3.4105
R5695 VCC.n2592 VCC.n2590 3.4105
R5696 VCC.n2625 VCC.n2624 3.4105
R5697 VCC.n2624 VCC.n2623 3.4105
R5698 VCC.n2321 VCC.n2320 3.4105
R5699 VCC.n2568 VCC.n2321 3.4105
R5700 VCC.n2589 VCC.n2318 3.4105
R5701 VCC.n2599 VCC.n2598 3.4105
R5702 VCC.n2599 VCC.n2317 3.4105
R5703 VCC.n2562 VCC.n2332 3.4105
R5704 VCC.n2562 VCC.n2561 3.4105
R5705 VCC.n2566 VCC.n2565 3.4105
R5706 VCC.n2537 VCC.n2536 3.4105
R5707 VCC.n2537 VCC.n2343 3.4105
R5708 VCC.n3308 VCC.n3307 3.4105
R5709 VCC.n3308 VCC.n2774 3.4105
R5710 VCC.n3284 VCC.n3283 3.4105
R5711 VCC.n3306 VCC.n3305 3.4105
R5712 VCC.n3305 VCC.n3304 3.4105
R5713 VCC.n3274 VCC.n2803 3.4105
R5714 VCC.n2803 VCC.n2802 3.4105
R5715 VCC.n3276 VCC.n3275 3.4105
R5716 VCC.n3282 VCC.n3281 3.4105
R5717 VCC.n3281 VCC.n3280 3.4105
R5718 VCC.n3256 VCC.n3255 3.4105
R5719 VCC.n3256 VCC.n2815 3.4105
R5720 VCC.n3252 VCC.n2805 3.4105
R5721 VCC.n3273 VCC.n3272 3.4105
R5722 VCC.n3272 VCC.n3271 3.4105
R5723 VCC.n3234 VCC.n3231 3.4105
R5724 VCC.n3234 VCC.n3233 3.4105
R5725 VCC.n3251 VCC.n3250 3.4105
R5726 VCC.n3230 VCC.n3229 3.4105
R5727 VCC.n3229 VCC.n3228 3.4105
R5728 VCC.n3214 VCC.n3213 3.4105
R5729 VCC.n3215 VCC.n3214 3.4105
R5730 VCC.n3179 VCC.n3178 3.4105
R5731 VCC.n3212 VCC.n3211 3.4105
R5732 VCC.n3211 VCC.n3210 3.4105
R5733 VCC.n3149 VCC.n3148 3.4105
R5734 VCC.n3148 VCC.n3147 3.4105
R5735 VCC.n3144 VCC.n3142 3.4105
R5736 VCC.n3177 VCC.n3176 3.4105
R5737 VCC.n3176 VCC.n3175 3.4105
R5738 VCC.n2873 VCC.n2872 3.4105
R5739 VCC.n3120 VCC.n2873 3.4105
R5740 VCC.n3141 VCC.n2870 3.4105
R5741 VCC.n3151 VCC.n3150 3.4105
R5742 VCC.n3151 VCC.n2869 3.4105
R5743 VCC.n3114 VCC.n2884 3.4105
R5744 VCC.n3114 VCC.n3113 3.4105
R5745 VCC.n3118 VCC.n3117 3.4105
R5746 VCC.n3088 VCC.n3087 3.4105
R5747 VCC.n3088 VCC.n2895 3.4105
R5748 VCC.n3079 VCC.n3078 3.4105
R5749 VCC.n3080 VCC.n3079 3.4105
R5750 VCC.n3052 VCC.n3051 3.4105
R5751 VCC.n3077 VCC.n3076 3.4105
R5752 VCC.n3076 VCC.n3075 3.4105
R5753 VCC.n3028 VCC.n2933 3.4105
R5754 VCC.n2933 VCC.n2927 3.4105
R5755 VCC.n3030 VCC.n3029 3.4105
R5756 VCC.n3050 VCC.n3049 3.4105
R5757 VCC.n3049 VCC.n3048 3.4105
R5758 VCC.n3012 VCC.n2941 3.4105
R5759 VCC.n2941 VCC.n2940 3.4105
R5760 VCC.n2942 VCC.n2935 3.4105
R5761 VCC.n3027 VCC.n3026 3.4105
R5762 VCC.n3026 VCC.n3025 3.4105
R5763 VCC.n2989 VCC.n2988 3.4105
R5764 VCC.n2990 VCC.n2989 3.4105
R5765 VCC.n3011 VCC.n3010 3.4105
R5766 VCC.n2987 VCC.n2986 3.4105
R5767 VCC.n2986 VCC.n2985 3.4105
R5768 VCC.n3637 VCC.n3636 3.4105
R5769 VCC.n3638 VCC.n3637 3.4105
R5770 VCC.n3610 VCC.n3609 3.4105
R5771 VCC.n3635 VCC.n3634 3.4105
R5772 VCC.n3634 VCC.n3633 3.4105
R5773 VCC.n3586 VCC.n3491 3.4105
R5774 VCC.n3491 VCC.n3485 3.4105
R5775 VCC.n3588 VCC.n3587 3.4105
R5776 VCC.n3608 VCC.n3607 3.4105
R5777 VCC.n3607 VCC.n3606 3.4105
R5778 VCC.n3570 VCC.n3499 3.4105
R5779 VCC.n3499 VCC.n3498 3.4105
R5780 VCC.n3500 VCC.n3493 3.4105
R5781 VCC.n3585 VCC.n3584 3.4105
R5782 VCC.n3584 VCC.n3583 3.4105
R5783 VCC.n3547 VCC.n3546 3.4105
R5784 VCC.n3548 VCC.n3547 3.4105
R5785 VCC.n3569 VCC.n3568 3.4105
R5786 VCC.n3545 VCC.n3544 3.4105
R5787 VCC.n3544 VCC.n3543 3.4105
R5788 VCC.n3789 VCC.n3788 3.4105
R5789 VCC.n3788 VCC.n3787 3.4105
R5790 VCC.n3848 VCC.n3847 3.4105
R5791 VCC.n3853 VCC.n3852 3.4105
R5792 VCC.n3852 VCC.n3851 3.4105
R5793 VCC.n3831 VCC.n3830 3.4105
R5794 VCC.n3832 VCC.n3831 3.4105
R5795 VCC.n3829 VCC.n3828 3.4105
R5796 VCC.n3846 VCC.n3845 3.4105
R5797 VCC.n3845 VCC.n3844 3.4105
R5798 VCC.n3818 VCC.n3371 3.4105
R5799 VCC.n3371 VCC.n3370 3.4105
R5800 VCC.n3369 VCC.n3368 3.4105
R5801 VCC.n3826 VCC.n3825 3.4105
R5802 VCC.n3825 VCC.n3364 3.4105
R5803 VCC.n3791 VCC.n3790 3.4105
R5804 VCC.n3791 VCC.n3387 3.4105
R5805 VCC.n3817 VCC.n3816 3.4105
R5806 VCC.n3855 VCC.n3854 3.4105
R5807 VCC.n3855 VCC.n3328 3.4105
R5808 VCC.n3772 VCC.n3771 3.4105
R5809 VCC.n3773 VCC.n3772 3.4105
R5810 VCC.n3736 VCC.n3735 3.4105
R5811 VCC.n3770 VCC.n3769 3.4105
R5812 VCC.n3769 VCC.n3768 3.4105
R5813 VCC.n3706 VCC.n3705 3.4105
R5814 VCC.n3705 VCC.n3704 3.4105
R5815 VCC.n3701 VCC.n3699 3.4105
R5816 VCC.n3734 VCC.n3733 3.4105
R5817 VCC.n3733 VCC.n3732 3.4105
R5818 VCC.n3430 VCC.n3429 3.4105
R5819 VCC.n3677 VCC.n3430 3.4105
R5820 VCC.n3698 VCC.n3427 3.4105
R5821 VCC.n3708 VCC.n3707 3.4105
R5822 VCC.n3708 VCC.n3426 3.4105
R5823 VCC.n3671 VCC.n3441 3.4105
R5824 VCC.n3671 VCC.n3670 3.4105
R5825 VCC.n3675 VCC.n3674 3.4105
R5826 VCC.n3646 VCC.n3645 3.4105
R5827 VCC.n3646 VCC.n3452 3.4105
R5828 VCC.n4417 VCC.n4416 3.4105
R5829 VCC.n4417 VCC.n3883 3.4105
R5830 VCC.n4393 VCC.n4392 3.4105
R5831 VCC.n4415 VCC.n4414 3.4105
R5832 VCC.n4414 VCC.n4413 3.4105
R5833 VCC.n4383 VCC.n3912 3.4105
R5834 VCC.n3912 VCC.n3911 3.4105
R5835 VCC.n4385 VCC.n4384 3.4105
R5836 VCC.n4391 VCC.n4390 3.4105
R5837 VCC.n4390 VCC.n4389 3.4105
R5838 VCC.n4365 VCC.n4364 3.4105
R5839 VCC.n4365 VCC.n3924 3.4105
R5840 VCC.n4361 VCC.n3914 3.4105
R5841 VCC.n4382 VCC.n4381 3.4105
R5842 VCC.n4381 VCC.n4380 3.4105
R5843 VCC.n4343 VCC.n4340 3.4105
R5844 VCC.n4343 VCC.n4342 3.4105
R5845 VCC.n4360 VCC.n4359 3.4105
R5846 VCC.n4339 VCC.n4338 3.4105
R5847 VCC.n4338 VCC.n4337 3.4105
R5848 VCC.n4323 VCC.n4322 3.4105
R5849 VCC.n4324 VCC.n4323 3.4105
R5850 VCC.n4288 VCC.n4287 3.4105
R5851 VCC.n4321 VCC.n4320 3.4105
R5852 VCC.n4320 VCC.n4319 3.4105
R5853 VCC.n4258 VCC.n4257 3.4105
R5854 VCC.n4257 VCC.n4256 3.4105
R5855 VCC.n4253 VCC.n4251 3.4105
R5856 VCC.n4286 VCC.n4285 3.4105
R5857 VCC.n4285 VCC.n4284 3.4105
R5858 VCC.n3982 VCC.n3981 3.4105
R5859 VCC.n4229 VCC.n3982 3.4105
R5860 VCC.n4250 VCC.n3979 3.4105
R5861 VCC.n4260 VCC.n4259 3.4105
R5862 VCC.n4260 VCC.n3978 3.4105
R5863 VCC.n4223 VCC.n3993 3.4105
R5864 VCC.n4223 VCC.n4222 3.4105
R5865 VCC.n4227 VCC.n4226 3.4105
R5866 VCC.n4197 VCC.n4196 3.4105
R5867 VCC.n4197 VCC.n4004 3.4105
R5868 VCC.n4188 VCC.n4187 3.4105
R5869 VCC.n4189 VCC.n4188 3.4105
R5870 VCC.n4161 VCC.n4160 3.4105
R5871 VCC.n4186 VCC.n4185 3.4105
R5872 VCC.n4185 VCC.n4184 3.4105
R5873 VCC.n4137 VCC.n4042 3.4105
R5874 VCC.n4042 VCC.n4036 3.4105
R5875 VCC.n4139 VCC.n4138 3.4105
R5876 VCC.n4159 VCC.n4158 3.4105
R5877 VCC.n4158 VCC.n4157 3.4105
R5878 VCC.n4121 VCC.n4050 3.4105
R5879 VCC.n4050 VCC.n4049 3.4105
R5880 VCC.n4051 VCC.n4044 3.4105
R5881 VCC.n4136 VCC.n4135 3.4105
R5882 VCC.n4135 VCC.n4134 3.4105
R5883 VCC.n4098 VCC.n4097 3.4105
R5884 VCC.n4099 VCC.n4098 3.4105
R5885 VCC.n4120 VCC.n4119 3.4105
R5886 VCC.n4096 VCC.n4095 3.4105
R5887 VCC.n4095 VCC.n4094 3.4105
R5888 VCC.n4746 VCC.n4745 3.4105
R5889 VCC.n4747 VCC.n4746 3.4105
R5890 VCC.n4719 VCC.n4718 3.4105
R5891 VCC.n4744 VCC.n4743 3.4105
R5892 VCC.n4743 VCC.n4742 3.4105
R5893 VCC.n4695 VCC.n4600 3.4105
R5894 VCC.n4600 VCC.n4594 3.4105
R5895 VCC.n4697 VCC.n4696 3.4105
R5896 VCC.n4717 VCC.n4716 3.4105
R5897 VCC.n4716 VCC.n4715 3.4105
R5898 VCC.n4679 VCC.n4608 3.4105
R5899 VCC.n4608 VCC.n4607 3.4105
R5900 VCC.n4609 VCC.n4602 3.4105
R5901 VCC.n4694 VCC.n4693 3.4105
R5902 VCC.n4693 VCC.n4692 3.4105
R5903 VCC.n4656 VCC.n4655 3.4105
R5904 VCC.n4657 VCC.n4656 3.4105
R5905 VCC.n4678 VCC.n4677 3.4105
R5906 VCC.n4654 VCC.n4653 3.4105
R5907 VCC.n4653 VCC.n4652 3.4105
R5908 VCC.n4898 VCC.n4897 3.4105
R5909 VCC.n4897 VCC.n4896 3.4105
R5910 VCC.n4957 VCC.n4956 3.4105
R5911 VCC.n4962 VCC.n4961 3.4105
R5912 VCC.n4961 VCC.n4960 3.4105
R5913 VCC.n4940 VCC.n4939 3.4105
R5914 VCC.n4941 VCC.n4940 3.4105
R5915 VCC.n4938 VCC.n4937 3.4105
R5916 VCC.n4955 VCC.n4954 3.4105
R5917 VCC.n4954 VCC.n4953 3.4105
R5918 VCC.n4927 VCC.n4480 3.4105
R5919 VCC.n4480 VCC.n4479 3.4105
R5920 VCC.n4478 VCC.n4477 3.4105
R5921 VCC.n4935 VCC.n4934 3.4105
R5922 VCC.n4934 VCC.n4473 3.4105
R5923 VCC.n4900 VCC.n4899 3.4105
R5924 VCC.n4900 VCC.n4496 3.4105
R5925 VCC.n4926 VCC.n4925 3.4105
R5926 VCC.n4964 VCC.n4963 3.4105
R5927 VCC.n4964 VCC.n4437 3.4105
R5928 VCC.n4881 VCC.n4880 3.4105
R5929 VCC.n4882 VCC.n4881 3.4105
R5930 VCC.n4845 VCC.n4844 3.4105
R5931 VCC.n4879 VCC.n4878 3.4105
R5932 VCC.n4878 VCC.n4877 3.4105
R5933 VCC.n4815 VCC.n4814 3.4105
R5934 VCC.n4814 VCC.n4813 3.4105
R5935 VCC.n4810 VCC.n4808 3.4105
R5936 VCC.n4843 VCC.n4842 3.4105
R5937 VCC.n4842 VCC.n4841 3.4105
R5938 VCC.n4539 VCC.n4538 3.4105
R5939 VCC.n4786 VCC.n4539 3.4105
R5940 VCC.n4807 VCC.n4536 3.4105
R5941 VCC.n4817 VCC.n4816 3.4105
R5942 VCC.n4817 VCC.n4535 3.4105
R5943 VCC.n4780 VCC.n4550 3.4105
R5944 VCC.n4780 VCC.n4779 3.4105
R5945 VCC.n4784 VCC.n4783 3.4105
R5946 VCC.n4755 VCC.n4754 3.4105
R5947 VCC.n4755 VCC.n4561 3.4105
R5948 VCC.n5526 VCC.n5525 3.4105
R5949 VCC.n5526 VCC.n4992 3.4105
R5950 VCC.n5502 VCC.n5501 3.4105
R5951 VCC.n5524 VCC.n5523 3.4105
R5952 VCC.n5523 VCC.n5522 3.4105
R5953 VCC.n5492 VCC.n5021 3.4105
R5954 VCC.n5021 VCC.n5020 3.4105
R5955 VCC.n5494 VCC.n5493 3.4105
R5956 VCC.n5500 VCC.n5499 3.4105
R5957 VCC.n5499 VCC.n5498 3.4105
R5958 VCC.n5474 VCC.n5473 3.4105
R5959 VCC.n5474 VCC.n5033 3.4105
R5960 VCC.n5470 VCC.n5023 3.4105
R5961 VCC.n5491 VCC.n5490 3.4105
R5962 VCC.n5490 VCC.n5489 3.4105
R5963 VCC.n5452 VCC.n5449 3.4105
R5964 VCC.n5452 VCC.n5451 3.4105
R5965 VCC.n5469 VCC.n5468 3.4105
R5966 VCC.n5448 VCC.n5447 3.4105
R5967 VCC.n5447 VCC.n5446 3.4105
R5968 VCC.n5432 VCC.n5431 3.4105
R5969 VCC.n5433 VCC.n5432 3.4105
R5970 VCC.n5397 VCC.n5396 3.4105
R5971 VCC.n5430 VCC.n5429 3.4105
R5972 VCC.n5429 VCC.n5428 3.4105
R5973 VCC.n5367 VCC.n5366 3.4105
R5974 VCC.n5366 VCC.n5365 3.4105
R5975 VCC.n5362 VCC.n5360 3.4105
R5976 VCC.n5395 VCC.n5394 3.4105
R5977 VCC.n5394 VCC.n5393 3.4105
R5978 VCC.n5091 VCC.n5090 3.4105
R5979 VCC.n5338 VCC.n5091 3.4105
R5980 VCC.n5359 VCC.n5088 3.4105
R5981 VCC.n5369 VCC.n5368 3.4105
R5982 VCC.n5369 VCC.n5087 3.4105
R5983 VCC.n5332 VCC.n5102 3.4105
R5984 VCC.n5332 VCC.n5331 3.4105
R5985 VCC.n5336 VCC.n5335 3.4105
R5986 VCC.n5306 VCC.n5305 3.4105
R5987 VCC.n5306 VCC.n5113 3.4105
R5988 VCC.n5297 VCC.n5296 3.4105
R5989 VCC.n5298 VCC.n5297 3.4105
R5990 VCC.n5270 VCC.n5269 3.4105
R5991 VCC.n5295 VCC.n5294 3.4105
R5992 VCC.n5294 VCC.n5293 3.4105
R5993 VCC.n5246 VCC.n5151 3.4105
R5994 VCC.n5151 VCC.n5145 3.4105
R5995 VCC.n5248 VCC.n5247 3.4105
R5996 VCC.n5268 VCC.n5267 3.4105
R5997 VCC.n5267 VCC.n5266 3.4105
R5998 VCC.n5230 VCC.n5159 3.4105
R5999 VCC.n5159 VCC.n5158 3.4105
R6000 VCC.n5160 VCC.n5153 3.4105
R6001 VCC.n5245 VCC.n5244 3.4105
R6002 VCC.n5244 VCC.n5243 3.4105
R6003 VCC.n5207 VCC.n5206 3.4105
R6004 VCC.n5208 VCC.n5207 3.4105
R6005 VCC.n5229 VCC.n5228 3.4105
R6006 VCC.n5205 VCC.n5204 3.4105
R6007 VCC.n5204 VCC.n5203 3.4105
R6008 VCC.n5854 VCC.n5853 3.4105
R6009 VCC.n5855 VCC.n5854 3.4105
R6010 VCC.n5827 VCC.n5826 3.4105
R6011 VCC.n5852 VCC.n5851 3.4105
R6012 VCC.n5851 VCC.n5850 3.4105
R6013 VCC.n5803 VCC.n5708 3.4105
R6014 VCC.n5708 VCC.n5702 3.4105
R6015 VCC.n5805 VCC.n5804 3.4105
R6016 VCC.n5825 VCC.n5824 3.4105
R6017 VCC.n5824 VCC.n5823 3.4105
R6018 VCC.n5787 VCC.n5716 3.4105
R6019 VCC.n5716 VCC.n5715 3.4105
R6020 VCC.n5717 VCC.n5710 3.4105
R6021 VCC.n5802 VCC.n5801 3.4105
R6022 VCC.n5801 VCC.n5800 3.4105
R6023 VCC.n5764 VCC.n5763 3.4105
R6024 VCC.n5765 VCC.n5764 3.4105
R6025 VCC.n5786 VCC.n5785 3.4105
R6026 VCC.n5762 VCC.n5761 3.4105
R6027 VCC.n5761 VCC.n5760 3.4105
R6028 VCC.n6006 VCC.n6005 3.4105
R6029 VCC.n6005 VCC.n6004 3.4105
R6030 VCC.n6065 VCC.n6064 3.4105
R6031 VCC.n6070 VCC.n6069 3.4105
R6032 VCC.n6069 VCC.n6068 3.4105
R6033 VCC.n6048 VCC.n6047 3.4105
R6034 VCC.n6049 VCC.n6048 3.4105
R6035 VCC.n6046 VCC.n6045 3.4105
R6036 VCC.n6063 VCC.n6062 3.4105
R6037 VCC.n6062 VCC.n6061 3.4105
R6038 VCC.n6035 VCC.n5588 3.4105
R6039 VCC.n5588 VCC.n5587 3.4105
R6040 VCC.n5586 VCC.n5585 3.4105
R6041 VCC.n6043 VCC.n6042 3.4105
R6042 VCC.n6042 VCC.n5581 3.4105
R6043 VCC.n6008 VCC.n6007 3.4105
R6044 VCC.n6008 VCC.n5604 3.4105
R6045 VCC.n6034 VCC.n6033 3.4105
R6046 VCC.n6072 VCC.n6071 3.4105
R6047 VCC.n6072 VCC.n5545 3.4105
R6048 VCC.n5989 VCC.n5988 3.4105
R6049 VCC.n5990 VCC.n5989 3.4105
R6050 VCC.n5953 VCC.n5952 3.4105
R6051 VCC.n5987 VCC.n5986 3.4105
R6052 VCC.n5986 VCC.n5985 3.4105
R6053 VCC.n5923 VCC.n5922 3.4105
R6054 VCC.n5922 VCC.n5921 3.4105
R6055 VCC.n5918 VCC.n5916 3.4105
R6056 VCC.n5951 VCC.n5950 3.4105
R6057 VCC.n5950 VCC.n5949 3.4105
R6058 VCC.n5647 VCC.n5646 3.4105
R6059 VCC.n5894 VCC.n5647 3.4105
R6060 VCC.n5915 VCC.n5644 3.4105
R6061 VCC.n5925 VCC.n5924 3.4105
R6062 VCC.n5925 VCC.n5643 3.4105
R6063 VCC.n5888 VCC.n5658 3.4105
R6064 VCC.n5888 VCC.n5887 3.4105
R6065 VCC.n5892 VCC.n5891 3.4105
R6066 VCC.n5863 VCC.n5862 3.4105
R6067 VCC.n5863 VCC.n5669 3.4105
R6068 VCC.n6633 VCC.n6632 3.4105
R6069 VCC.n6633 VCC.n6099 3.4105
R6070 VCC.n6609 VCC.n6608 3.4105
R6071 VCC.n6631 VCC.n6630 3.4105
R6072 VCC.n6630 VCC.n6629 3.4105
R6073 VCC.n6599 VCC.n6128 3.4105
R6074 VCC.n6128 VCC.n6127 3.4105
R6075 VCC.n6601 VCC.n6600 3.4105
R6076 VCC.n6607 VCC.n6606 3.4105
R6077 VCC.n6606 VCC.n6605 3.4105
R6078 VCC.n6581 VCC.n6580 3.4105
R6079 VCC.n6581 VCC.n6140 3.4105
R6080 VCC.n6577 VCC.n6130 3.4105
R6081 VCC.n6598 VCC.n6597 3.4105
R6082 VCC.n6597 VCC.n6596 3.4105
R6083 VCC.n6559 VCC.n6556 3.4105
R6084 VCC.n6559 VCC.n6558 3.4105
R6085 VCC.n6576 VCC.n6575 3.4105
R6086 VCC.n6555 VCC.n6554 3.4105
R6087 VCC.n6554 VCC.n6553 3.4105
R6088 VCC.n6539 VCC.n6538 3.4105
R6089 VCC.n6540 VCC.n6539 3.4105
R6090 VCC.n6504 VCC.n6503 3.4105
R6091 VCC.n6537 VCC.n6536 3.4105
R6092 VCC.n6536 VCC.n6535 3.4105
R6093 VCC.n6474 VCC.n6473 3.4105
R6094 VCC.n6473 VCC.n6472 3.4105
R6095 VCC.n6469 VCC.n6467 3.4105
R6096 VCC.n6502 VCC.n6501 3.4105
R6097 VCC.n6501 VCC.n6500 3.4105
R6098 VCC.n6198 VCC.n6197 3.4105
R6099 VCC.n6445 VCC.n6198 3.4105
R6100 VCC.n6466 VCC.n6195 3.4105
R6101 VCC.n6476 VCC.n6475 3.4105
R6102 VCC.n6476 VCC.n6194 3.4105
R6103 VCC.n6439 VCC.n6209 3.4105
R6104 VCC.n6439 VCC.n6438 3.4105
R6105 VCC.n6443 VCC.n6442 3.4105
R6106 VCC.n6413 VCC.n6412 3.4105
R6107 VCC.n6413 VCC.n6220 3.4105
R6108 VCC.n6404 VCC.n6403 3.4105
R6109 VCC.n6405 VCC.n6404 3.4105
R6110 VCC.n6377 VCC.n6376 3.4105
R6111 VCC.n6402 VCC.n6401 3.4105
R6112 VCC.n6401 VCC.n6400 3.4105
R6113 VCC.n6353 VCC.n6258 3.4105
R6114 VCC.n6258 VCC.n6252 3.4105
R6115 VCC.n6355 VCC.n6354 3.4105
R6116 VCC.n6375 VCC.n6374 3.4105
R6117 VCC.n6374 VCC.n6373 3.4105
R6118 VCC.n6337 VCC.n6266 3.4105
R6119 VCC.n6266 VCC.n6265 3.4105
R6120 VCC.n6267 VCC.n6260 3.4105
R6121 VCC.n6352 VCC.n6351 3.4105
R6122 VCC.n6351 VCC.n6350 3.4105
R6123 VCC.n6314 VCC.n6313 3.4105
R6124 VCC.n6315 VCC.n6314 3.4105
R6125 VCC.n6336 VCC.n6335 3.4105
R6126 VCC.n6312 VCC.n6311 3.4105
R6127 VCC.n6311 VCC.n6310 3.4105
R6128 VCC.n6961 VCC.n6960 3.4105
R6129 VCC.n6962 VCC.n6961 3.4105
R6130 VCC.n6934 VCC.n6933 3.4105
R6131 VCC.n6959 VCC.n6958 3.4105
R6132 VCC.n6958 VCC.n6957 3.4105
R6133 VCC.n6910 VCC.n6815 3.4105
R6134 VCC.n6815 VCC.n6809 3.4105
R6135 VCC.n6912 VCC.n6911 3.4105
R6136 VCC.n6932 VCC.n6931 3.4105
R6137 VCC.n6931 VCC.n6930 3.4105
R6138 VCC.n6894 VCC.n6823 3.4105
R6139 VCC.n6823 VCC.n6822 3.4105
R6140 VCC.n6824 VCC.n6817 3.4105
R6141 VCC.n6909 VCC.n6908 3.4105
R6142 VCC.n6908 VCC.n6907 3.4105
R6143 VCC.n6871 VCC.n6870 3.4105
R6144 VCC.n6872 VCC.n6871 3.4105
R6145 VCC.n6893 VCC.n6892 3.4105
R6146 VCC.n6869 VCC.n6868 3.4105
R6147 VCC.n6868 VCC.n6867 3.4105
R6148 VCC.n7113 VCC.n7112 3.4105
R6149 VCC.n7112 VCC.n7111 3.4105
R6150 VCC.n7172 VCC.n7171 3.4105
R6151 VCC.n7177 VCC.n7176 3.4105
R6152 VCC.n7176 VCC.n7175 3.4105
R6153 VCC.n7155 VCC.n7154 3.4105
R6154 VCC.n7156 VCC.n7155 3.4105
R6155 VCC.n7153 VCC.n7152 3.4105
R6156 VCC.n7170 VCC.n7169 3.4105
R6157 VCC.n7169 VCC.n7168 3.4105
R6158 VCC.n7142 VCC.n6695 3.4105
R6159 VCC.n6695 VCC.n6694 3.4105
R6160 VCC.n6693 VCC.n6692 3.4105
R6161 VCC.n7150 VCC.n7149 3.4105
R6162 VCC.n7149 VCC.n6688 3.4105
R6163 VCC.n7115 VCC.n7114 3.4105
R6164 VCC.n7115 VCC.n6711 3.4105
R6165 VCC.n7141 VCC.n7140 3.4105
R6166 VCC.n7179 VCC.n7178 3.4105
R6167 VCC.n7179 VCC.n6652 3.4105
R6168 VCC.n7096 VCC.n7095 3.4105
R6169 VCC.n7097 VCC.n7096 3.4105
R6170 VCC.n7060 VCC.n7059 3.4105
R6171 VCC.n7094 VCC.n7093 3.4105
R6172 VCC.n7093 VCC.n7092 3.4105
R6173 VCC.n7030 VCC.n7029 3.4105
R6174 VCC.n7029 VCC.n7028 3.4105
R6175 VCC.n7025 VCC.n7023 3.4105
R6176 VCC.n7058 VCC.n7057 3.4105
R6177 VCC.n7057 VCC.n7056 3.4105
R6178 VCC.n6754 VCC.n6753 3.4105
R6179 VCC.n7001 VCC.n6754 3.4105
R6180 VCC.n7022 VCC.n6751 3.4105
R6181 VCC.n7032 VCC.n7031 3.4105
R6182 VCC.n7032 VCC.n6750 3.4105
R6183 VCC.n6995 VCC.n6765 3.4105
R6184 VCC.n6995 VCC.n6994 3.4105
R6185 VCC.n6999 VCC.n6998 3.4105
R6186 VCC.n6970 VCC.n6969 3.4105
R6187 VCC.n6970 VCC.n6776 3.4105
R6188 VCC.n7740 VCC.n7739 3.4105
R6189 VCC.n7740 VCC.n7206 3.4105
R6190 VCC.n7716 VCC.n7715 3.4105
R6191 VCC.n7738 VCC.n7737 3.4105
R6192 VCC.n7737 VCC.n7736 3.4105
R6193 VCC.n7706 VCC.n7235 3.4105
R6194 VCC.n7235 VCC.n7234 3.4105
R6195 VCC.n7708 VCC.n7707 3.4105
R6196 VCC.n7714 VCC.n7713 3.4105
R6197 VCC.n7713 VCC.n7712 3.4105
R6198 VCC.n7688 VCC.n7687 3.4105
R6199 VCC.n7688 VCC.n7247 3.4105
R6200 VCC.n7684 VCC.n7237 3.4105
R6201 VCC.n7705 VCC.n7704 3.4105
R6202 VCC.n7704 VCC.n7703 3.4105
R6203 VCC.n7666 VCC.n7663 3.4105
R6204 VCC.n7666 VCC.n7665 3.4105
R6205 VCC.n7683 VCC.n7682 3.4105
R6206 VCC.n7662 VCC.n7661 3.4105
R6207 VCC.n7661 VCC.n7660 3.4105
R6208 VCC.n7646 VCC.n7645 3.4105
R6209 VCC.n7647 VCC.n7646 3.4105
R6210 VCC.n7611 VCC.n7610 3.4105
R6211 VCC.n7644 VCC.n7643 3.4105
R6212 VCC.n7643 VCC.n7642 3.4105
R6213 VCC.n7581 VCC.n7580 3.4105
R6214 VCC.n7580 VCC.n7579 3.4105
R6215 VCC.n7576 VCC.n7574 3.4105
R6216 VCC.n7609 VCC.n7608 3.4105
R6217 VCC.n7608 VCC.n7607 3.4105
R6218 VCC.n7305 VCC.n7304 3.4105
R6219 VCC.n7552 VCC.n7305 3.4105
R6220 VCC.n7573 VCC.n7302 3.4105
R6221 VCC.n7583 VCC.n7582 3.4105
R6222 VCC.n7583 VCC.n7301 3.4105
R6223 VCC.n7546 VCC.n7316 3.4105
R6224 VCC.n7546 VCC.n7545 3.4105
R6225 VCC.n7550 VCC.n7549 3.4105
R6226 VCC.n7520 VCC.n7519 3.4105
R6227 VCC.n7520 VCC.n7327 3.4105
R6228 VCC.n7511 VCC.n7510 3.4105
R6229 VCC.n7512 VCC.n7511 3.4105
R6230 VCC.n7484 VCC.n7483 3.4105
R6231 VCC.n7509 VCC.n7508 3.4105
R6232 VCC.n7508 VCC.n7507 3.4105
R6233 VCC.n7460 VCC.n7365 3.4105
R6234 VCC.n7365 VCC.n7359 3.4105
R6235 VCC.n7462 VCC.n7461 3.4105
R6236 VCC.n7482 VCC.n7481 3.4105
R6237 VCC.n7481 VCC.n7480 3.4105
R6238 VCC.n7444 VCC.n7373 3.4105
R6239 VCC.n7373 VCC.n7372 3.4105
R6240 VCC.n7374 VCC.n7367 3.4105
R6241 VCC.n7459 VCC.n7458 3.4105
R6242 VCC.n7458 VCC.n7457 3.4105
R6243 VCC.n7421 VCC.n7420 3.4105
R6244 VCC.n7422 VCC.n7421 3.4105
R6245 VCC.n7443 VCC.n7442 3.4105
R6246 VCC.n7419 VCC.n7418 3.4105
R6247 VCC.n7418 VCC.n7417 3.4105
R6248 VCC.n8068 VCC.n8067 3.4105
R6249 VCC.n8069 VCC.n8068 3.4105
R6250 VCC.n8041 VCC.n8040 3.4105
R6251 VCC.n8066 VCC.n8065 3.4105
R6252 VCC.n8065 VCC.n8064 3.4105
R6253 VCC.n8017 VCC.n7922 3.4105
R6254 VCC.n7922 VCC.n7916 3.4105
R6255 VCC.n8019 VCC.n8018 3.4105
R6256 VCC.n8039 VCC.n8038 3.4105
R6257 VCC.n8038 VCC.n8037 3.4105
R6258 VCC.n8001 VCC.n7930 3.4105
R6259 VCC.n7930 VCC.n7929 3.4105
R6260 VCC.n7931 VCC.n7924 3.4105
R6261 VCC.n8016 VCC.n8015 3.4105
R6262 VCC.n8015 VCC.n8014 3.4105
R6263 VCC.n7978 VCC.n7977 3.4105
R6264 VCC.n7979 VCC.n7978 3.4105
R6265 VCC.n8000 VCC.n7999 3.4105
R6266 VCC.n7976 VCC.n7975 3.4105
R6267 VCC.n7975 VCC.n7974 3.4105
R6268 VCC.n8220 VCC.n8219 3.4105
R6269 VCC.n8219 VCC.n8218 3.4105
R6270 VCC.n8279 VCC.n8278 3.4105
R6271 VCC.n8284 VCC.n8283 3.4105
R6272 VCC.n8283 VCC.n8282 3.4105
R6273 VCC.n8262 VCC.n8261 3.4105
R6274 VCC.n8263 VCC.n8262 3.4105
R6275 VCC.n8260 VCC.n8259 3.4105
R6276 VCC.n8277 VCC.n8276 3.4105
R6277 VCC.n8276 VCC.n8275 3.4105
R6278 VCC.n8249 VCC.n7802 3.4105
R6279 VCC.n7802 VCC.n7801 3.4105
R6280 VCC.n7800 VCC.n7799 3.4105
R6281 VCC.n8257 VCC.n8256 3.4105
R6282 VCC.n8256 VCC.n7795 3.4105
R6283 VCC.n8222 VCC.n8221 3.4105
R6284 VCC.n8222 VCC.n7818 3.4105
R6285 VCC.n8248 VCC.n8247 3.4105
R6286 VCC.n8286 VCC.n8285 3.4105
R6287 VCC.n8286 VCC.n7759 3.4105
R6288 VCC.n8203 VCC.n8202 3.4105
R6289 VCC.n8204 VCC.n8203 3.4105
R6290 VCC.n8167 VCC.n8166 3.4105
R6291 VCC.n8201 VCC.n8200 3.4105
R6292 VCC.n8200 VCC.n8199 3.4105
R6293 VCC.n8137 VCC.n8136 3.4105
R6294 VCC.n8136 VCC.n8135 3.4105
R6295 VCC.n8132 VCC.n8130 3.4105
R6296 VCC.n8165 VCC.n8164 3.4105
R6297 VCC.n8164 VCC.n8163 3.4105
R6298 VCC.n7861 VCC.n7860 3.4105
R6299 VCC.n8108 VCC.n7861 3.4105
R6300 VCC.n8129 VCC.n7858 3.4105
R6301 VCC.n8139 VCC.n8138 3.4105
R6302 VCC.n8139 VCC.n7857 3.4105
R6303 VCC.n8102 VCC.n7872 3.4105
R6304 VCC.n8102 VCC.n8101 3.4105
R6305 VCC.n8106 VCC.n8105 3.4105
R6306 VCC.n8077 VCC.n8076 3.4105
R6307 VCC.n8077 VCC.n7883 3.4105
R6308 VCC.n8660 VCC.n8659 3.4105
R6309 VCC.n8660 VCC.n8313 3.4105
R6310 VCC.n8636 VCC.n8635 3.4105
R6311 VCC.n8658 VCC.n8657 3.4105
R6312 VCC.n8657 VCC.n8656 3.4105
R6313 VCC.n8626 VCC.n8342 3.4105
R6314 VCC.n8342 VCC.n8341 3.4105
R6315 VCC.n8628 VCC.n8627 3.4105
R6316 VCC.n8634 VCC.n8633 3.4105
R6317 VCC.n8633 VCC.n8632 3.4105
R6318 VCC.n8608 VCC.n8607 3.4105
R6319 VCC.n8608 VCC.n8354 3.4105
R6320 VCC.n8604 VCC.n8344 3.4105
R6321 VCC.n8625 VCC.n8624 3.4105
R6322 VCC.n8624 VCC.n8623 3.4105
R6323 VCC.n8586 VCC.n8583 3.4105
R6324 VCC.n8586 VCC.n8585 3.4105
R6325 VCC.n8603 VCC.n8602 3.4105
R6326 VCC.n8582 VCC.n8581 3.4105
R6327 VCC.n8581 VCC.n8580 3.4105
R6328 VCC.n8566 VCC.n8565 3.4105
R6329 VCC.n8567 VCC.n8566 3.4105
R6330 VCC.n8531 VCC.n8530 3.4105
R6331 VCC.n8564 VCC.n8563 3.4105
R6332 VCC.n8563 VCC.n8562 3.4105
R6333 VCC.n8501 VCC.n8500 3.4105
R6334 VCC.n8500 VCC.n8499 3.4105
R6335 VCC.n8496 VCC.n8494 3.4105
R6336 VCC.n8529 VCC.n8528 3.4105
R6337 VCC.n8528 VCC.n8527 3.4105
R6338 VCC.n8412 VCC.n8411 3.4105
R6339 VCC.n8472 VCC.n8412 3.4105
R6340 VCC.n8493 VCC.n8409 3.4105
R6341 VCC.n8503 VCC.n8502 3.4105
R6342 VCC.n8503 VCC.n8408 3.4105
R6343 VCC.n8466 VCC.n8423 3.4105
R6344 VCC.n8466 VCC.n8465 3.4105
R6345 VCC.n8470 VCC.n8469 3.4105
R6346 VCC.n8440 VCC.n8439 3.4105
R6347 VCC.n8440 VCC.n8434 3.4105
R6348 VCC.n421 VCC.n57 3.29193
R6349 VCC.n476 VCC.n475 3.29193
R6350 VCC.n515 VCC.n20 3.29193
R6351 VCC.n973 VCC.n609 3.29193
R6352 VCC.n1028 VCC.n1027 3.29193
R6353 VCC.n1067 VCC.n572 3.29193
R6354 VCC.n1531 VCC.n1165 3.29193
R6355 VCC.n1594 VCC.n1159 3.29193
R6356 VCC.n1140 VCC.n1116 3.29193
R6357 VCC.n2082 VCC.n1718 3.29193
R6358 VCC.n2137 VCC.n2136 3.29193
R6359 VCC.n2176 VCC.n1681 3.29193
R6360 VCC.n2640 VCC.n2274 3.29193
R6361 VCC.n2703 VCC.n2268 3.29193
R6362 VCC.n2249 VCC.n2225 3.29193
R6363 VCC.n3191 VCC.n2827 3.29193
R6364 VCC.n3246 VCC.n3245 3.29193
R6365 VCC.n3285 VCC.n2790 3.29193
R6366 VCC.n3749 VCC.n3383 3.29193
R6367 VCC.n3812 VCC.n3377 3.29193
R6368 VCC.n3358 VCC.n3334 3.29193
R6369 VCC.n4300 VCC.n3936 3.29193
R6370 VCC.n4355 VCC.n4354 3.29193
R6371 VCC.n4394 VCC.n3899 3.29193
R6372 VCC.n4858 VCC.n4492 3.29193
R6373 VCC.n4921 VCC.n4486 3.29193
R6374 VCC.n4467 VCC.n4443 3.29193
R6375 VCC.n5409 VCC.n5045 3.29193
R6376 VCC.n5464 VCC.n5463 3.29193
R6377 VCC.n5503 VCC.n5008 3.29193
R6378 VCC.n5966 VCC.n5600 3.29193
R6379 VCC.n6029 VCC.n5594 3.29193
R6380 VCC.n5575 VCC.n5551 3.29193
R6381 VCC.n6516 VCC.n6152 3.29193
R6382 VCC.n6571 VCC.n6570 3.29193
R6383 VCC.n6610 VCC.n6115 3.29193
R6384 VCC.n7073 VCC.n6707 3.29193
R6385 VCC.n7136 VCC.n6701 3.29193
R6386 VCC.n6682 VCC.n6658 3.29193
R6387 VCC.n7623 VCC.n7259 3.29193
R6388 VCC.n7678 VCC.n7677 3.29193
R6389 VCC.n7717 VCC.n7222 3.29193
R6390 VCC.n8180 VCC.n7814 3.29193
R6391 VCC.n8243 VCC.n7808 3.29193
R6392 VCC.n7789 VCC.n7765 3.29193
R6393 VCC.n8543 VCC.n8366 3.29193
R6394 VCC.n8598 VCC.n8597 3.29193
R6395 VCC.n8637 VCC.n8329 3.29193
R6396 VCC.n469 VCC.n55 3.25764
R6397 VCC.n528 VCC.n6 3.25764
R6398 VCC.n1021 VCC.n607 3.25764
R6399 VCC.n1080 VCC.n560 3.25764
R6400 VCC.n1579 VCC.n1164 3.25764
R6401 VCC.n1650 VCC.n1113 3.25764
R6402 VCC.n2130 VCC.n1716 3.25764
R6403 VCC.n2189 VCC.n1669 3.25764
R6404 VCC.n2688 VCC.n2273 3.25764
R6405 VCC.n2759 VCC.n2222 3.25764
R6406 VCC.n3239 VCC.n2825 3.25764
R6407 VCC.n3298 VCC.n2778 3.25764
R6408 VCC.n3797 VCC.n3382 3.25764
R6409 VCC.n3868 VCC.n3331 3.25764
R6410 VCC.n4348 VCC.n3934 3.25764
R6411 VCC.n4407 VCC.n3887 3.25764
R6412 VCC.n4906 VCC.n4491 3.25764
R6413 VCC.n4977 VCC.n4440 3.25764
R6414 VCC.n5457 VCC.n5043 3.25764
R6415 VCC.n5516 VCC.n4996 3.25764
R6416 VCC.n6014 VCC.n5599 3.25764
R6417 VCC.n6085 VCC.n5548 3.25764
R6418 VCC.n6564 VCC.n6150 3.25764
R6419 VCC.n6623 VCC.n6103 3.25764
R6420 VCC.n7121 VCC.n6706 3.25764
R6421 VCC.n7192 VCC.n6655 3.25764
R6422 VCC.n7671 VCC.n7257 3.25764
R6423 VCC.n7730 VCC.n7210 3.25764
R6424 VCC.n8228 VCC.n7813 3.25764
R6425 VCC.n8299 VCC.n7762 3.25764
R6426 VCC.n8591 VCC.n8364 3.25764
R6427 VCC.n8650 VCC.n8317 3.25764
R6428 VCC.n545 VCC.n544 3.2005
R6429 VCC.n1099 VCC.n1098 3.2005
R6430 VCC.n1124 VCC.n1112 3.2005
R6431 VCC.n2208 VCC.n2207 3.2005
R6432 VCC.n2233 VCC.n2221 3.2005
R6433 VCC.n3317 VCC.n3316 3.2005
R6434 VCC.n3342 VCC.n3330 3.2005
R6435 VCC.n4426 VCC.n4425 3.2005
R6436 VCC.n4451 VCC.n4439 3.2005
R6437 VCC.n5535 VCC.n5534 3.2005
R6438 VCC.n5559 VCC.n5547 3.2005
R6439 VCC.n6642 VCC.n6641 3.2005
R6440 VCC.n6666 VCC.n6654 3.2005
R6441 VCC.n7749 VCC.n7748 3.2005
R6442 VCC.n7773 VCC.n7761 3.2005
R6443 VCC.n8669 VCC.n8668 3.2005
R6444 VCC.n500 VCC.n499 3.03311
R6445 VCC.n468 VCC.n467 3.03311
R6446 VCC.n1020 VCC.n1019 3.03311
R6447 VCC.n1052 VCC.n1051 3.03311
R6448 VCC.n1616 VCC.n1615 3.03311
R6449 VCC.n1577 VCC.n1576 3.03311
R6450 VCC.n2129 VCC.n2128 3.03311
R6451 VCC.n2161 VCC.n2160 3.03311
R6452 VCC.n2725 VCC.n2724 3.03311
R6453 VCC.n2686 VCC.n2685 3.03311
R6454 VCC.n3238 VCC.n3237 3.03311
R6455 VCC.n3270 VCC.n3269 3.03311
R6456 VCC.n3834 VCC.n3833 3.03311
R6457 VCC.n3795 VCC.n3794 3.03311
R6458 VCC.n4347 VCC.n4346 3.03311
R6459 VCC.n4379 VCC.n4378 3.03311
R6460 VCC.n4943 VCC.n4942 3.03311
R6461 VCC.n4904 VCC.n4903 3.03311
R6462 VCC.n5456 VCC.n5455 3.03311
R6463 VCC.n5488 VCC.n5487 3.03311
R6464 VCC.n6051 VCC.n6050 3.03311
R6465 VCC.n6012 VCC.n6011 3.03311
R6466 VCC.n6563 VCC.n6562 3.03311
R6467 VCC.n6595 VCC.n6594 3.03311
R6468 VCC.n7158 VCC.n7157 3.03311
R6469 VCC.n7119 VCC.n7118 3.03311
R6470 VCC.n7670 VCC.n7669 3.03311
R6471 VCC.n7702 VCC.n7701 3.03311
R6472 VCC.n8265 VCC.n8264 3.03311
R6473 VCC.n8226 VCC.n8225 3.03311
R6474 VCC.n8590 VCC.n8589 3.03311
R6475 VCC.n8622 VCC.n8621 3.03311
R6476 VCC.n225 VCC.n182 2.8505
R6477 VCC.n292 VCC.n140 2.8505
R6478 VCC.n338 VCC.n119 2.8505
R6479 VCC.n416 VCC.n80 2.8505
R6480 VCC.n777 VCC.n734 2.8505
R6481 VCC.n844 VCC.n692 2.8505
R6482 VCC.n890 VCC.n671 2.8505
R6483 VCC.n968 VCC.n632 2.8505
R6484 VCC.n1447 VCC.n1228 2.8505
R6485 VCC.n1525 VCC.n1189 2.8505
R6486 VCC.n1335 VCC.n1292 2.8505
R6487 VCC.n1402 VCC.n1250 2.8505
R6488 VCC.n1886 VCC.n1843 2.8505
R6489 VCC.n1953 VCC.n1801 2.8505
R6490 VCC.n1999 VCC.n1780 2.8505
R6491 VCC.n2077 VCC.n1741 2.8505
R6492 VCC.n2556 VCC.n2337 2.8505
R6493 VCC.n2634 VCC.n2298 2.8505
R6494 VCC.n2444 VCC.n2401 2.8505
R6495 VCC.n2511 VCC.n2359 2.8505
R6496 VCC.n2995 VCC.n2952 2.8505
R6497 VCC.n3062 VCC.n2910 2.8505
R6498 VCC.n3108 VCC.n2889 2.8505
R6499 VCC.n3186 VCC.n2850 2.8505
R6500 VCC.n3665 VCC.n3446 2.8505
R6501 VCC.n3743 VCC.n3407 2.8505
R6502 VCC.n3553 VCC.n3510 2.8505
R6503 VCC.n3620 VCC.n3468 2.8505
R6504 VCC.n4104 VCC.n4061 2.8505
R6505 VCC.n4171 VCC.n4019 2.8505
R6506 VCC.n4217 VCC.n3998 2.8505
R6507 VCC.n4295 VCC.n3959 2.8505
R6508 VCC.n4774 VCC.n4555 2.8505
R6509 VCC.n4852 VCC.n4516 2.8505
R6510 VCC.n4662 VCC.n4619 2.8505
R6511 VCC.n4729 VCC.n4577 2.8505
R6512 VCC.n5213 VCC.n5170 2.8505
R6513 VCC.n5280 VCC.n5128 2.8505
R6514 VCC.n5326 VCC.n5107 2.8505
R6515 VCC.n5404 VCC.n5068 2.8505
R6516 VCC.n5882 VCC.n5663 2.8505
R6517 VCC.n5960 VCC.n5624 2.8505
R6518 VCC.n5770 VCC.n5727 2.8505
R6519 VCC.n5837 VCC.n5685 2.8505
R6520 VCC.n6320 VCC.n6277 2.8505
R6521 VCC.n6387 VCC.n6235 2.8505
R6522 VCC.n6433 VCC.n6214 2.8505
R6523 VCC.n6511 VCC.n6175 2.8505
R6524 VCC.n6989 VCC.n6770 2.8505
R6525 VCC.n7067 VCC.n6731 2.8505
R6526 VCC.n6877 VCC.n6834 2.8505
R6527 VCC.n6944 VCC.n6792 2.8505
R6528 VCC.n7427 VCC.n7384 2.8505
R6529 VCC.n7494 VCC.n7342 2.8505
R6530 VCC.n7540 VCC.n7321 2.8505
R6531 VCC.n7618 VCC.n7282 2.8505
R6532 VCC.n8096 VCC.n7877 2.8505
R6533 VCC.n8174 VCC.n7838 2.8505
R6534 VCC.n7984 VCC.n7941 2.8505
R6535 VCC.n8051 VCC.n7899 2.8505
R6536 VCC.n8460 VCC.n8428 2.8505
R6537 VCC.n8538 VCC.n8389 2.8505
R6538 VCC.n272 VCC.n271 2.5605
R6539 VCC.n399 VCC.n398 2.5605
R6540 VCC.n824 VCC.n823 2.5605
R6541 VCC.n951 VCC.n950 2.5605
R6542 VCC.n1508 VCC.n1507 2.5605
R6543 VCC.n1382 VCC.n1381 2.5605
R6544 VCC.n1933 VCC.n1932 2.5605
R6545 VCC.n2060 VCC.n2059 2.5605
R6546 VCC.n2617 VCC.n2616 2.5605
R6547 VCC.n2491 VCC.n2490 2.5605
R6548 VCC.n3042 VCC.n3041 2.5605
R6549 VCC.n3169 VCC.n3168 2.5605
R6550 VCC.n3726 VCC.n3725 2.5605
R6551 VCC.n3600 VCC.n3599 2.5605
R6552 VCC.n4151 VCC.n4150 2.5605
R6553 VCC.n4278 VCC.n4277 2.5605
R6554 VCC.n4835 VCC.n4834 2.5605
R6555 VCC.n4709 VCC.n4708 2.5605
R6556 VCC.n5260 VCC.n5259 2.5605
R6557 VCC.n5387 VCC.n5386 2.5605
R6558 VCC.n5943 VCC.n5942 2.5605
R6559 VCC.n5817 VCC.n5816 2.5605
R6560 VCC.n6367 VCC.n6366 2.5605
R6561 VCC.n6494 VCC.n6493 2.5605
R6562 VCC.n7050 VCC.n7049 2.5605
R6563 VCC.n6924 VCC.n6923 2.5605
R6564 VCC.n7474 VCC.n7473 2.5605
R6565 VCC.n7601 VCC.n7600 2.5605
R6566 VCC.n8157 VCC.n8156 2.5605
R6567 VCC.n8031 VCC.n8030 2.5605
R6568 VCC.n8521 VCC.n8520 2.5605
R6569 VCC.n232 VCC.n231 2.46907
R6570 VCC.n358 VCC.n357 2.46907
R6571 VCC.n784 VCC.n783 2.46907
R6572 VCC.n910 VCC.n909 2.46907
R6573 VCC.n1467 VCC.n1466 2.46907
R6574 VCC.n1342 VCC.n1341 2.46907
R6575 VCC.n1893 VCC.n1892 2.46907
R6576 VCC.n2019 VCC.n2018 2.46907
R6577 VCC.n2576 VCC.n2575 2.46907
R6578 VCC.n2451 VCC.n2450 2.46907
R6579 VCC.n3002 VCC.n3001 2.46907
R6580 VCC.n3128 VCC.n3127 2.46907
R6581 VCC.n3685 VCC.n3684 2.46907
R6582 VCC.n3560 VCC.n3559 2.46907
R6583 VCC.n4111 VCC.n4110 2.46907
R6584 VCC.n4237 VCC.n4236 2.46907
R6585 VCC.n4794 VCC.n4793 2.46907
R6586 VCC.n4669 VCC.n4668 2.46907
R6587 VCC.n5220 VCC.n5219 2.46907
R6588 VCC.n5346 VCC.n5345 2.46907
R6589 VCC.n5902 VCC.n5901 2.46907
R6590 VCC.n5777 VCC.n5776 2.46907
R6591 VCC.n6327 VCC.n6326 2.46907
R6592 VCC.n6453 VCC.n6452 2.46907
R6593 VCC.n7009 VCC.n7008 2.46907
R6594 VCC.n6884 VCC.n6883 2.46907
R6595 VCC.n7434 VCC.n7433 2.46907
R6596 VCC.n7560 VCC.n7559 2.46907
R6597 VCC.n8116 VCC.n8115 2.46907
R6598 VCC.n7991 VCC.n7990 2.46907
R6599 VCC.n8480 VCC.n8479 2.46907
R6600 VCC.n141 VCC.n139 2.37764
R6601 VCC.n414 VCC.n78 2.37764
R6602 VCC.n693 VCC.n691 2.37764
R6603 VCC.n966 VCC.n630 2.37764
R6604 VCC.n1523 VCC.n1187 2.37764
R6605 VCC.n1251 VCC.n1249 2.37764
R6606 VCC.n1802 VCC.n1800 2.37764
R6607 VCC.n2075 VCC.n1739 2.37764
R6608 VCC.n2632 VCC.n2296 2.37764
R6609 VCC.n2360 VCC.n2358 2.37764
R6610 VCC.n2911 VCC.n2909 2.37764
R6611 VCC.n3184 VCC.n2848 2.37764
R6612 VCC.n3741 VCC.n3405 2.37764
R6613 VCC.n3469 VCC.n3467 2.37764
R6614 VCC.n4020 VCC.n4018 2.37764
R6615 VCC.n4293 VCC.n3957 2.37764
R6616 VCC.n4850 VCC.n4514 2.37764
R6617 VCC.n4578 VCC.n4576 2.37764
R6618 VCC.n5129 VCC.n5127 2.37764
R6619 VCC.n5402 VCC.n5066 2.37764
R6620 VCC.n5958 VCC.n5622 2.37764
R6621 VCC.n5686 VCC.n5684 2.37764
R6622 VCC.n6236 VCC.n6234 2.37764
R6623 VCC.n6509 VCC.n6173 2.37764
R6624 VCC.n7065 VCC.n6729 2.37764
R6625 VCC.n6793 VCC.n6791 2.37764
R6626 VCC.n7343 VCC.n7341 2.37764
R6627 VCC.n7616 VCC.n7280 2.37764
R6628 VCC.n8172 VCC.n7836 2.37764
R6629 VCC.n7900 VCC.n7898 2.37764
R6630 VCC.n8536 VCC.n8387 2.37764
R6631 VCC.n208 VCC.n194 2.34304
R6632 VCC.n81 VCC.n79 2.34304
R6633 VCC.n123 VCC.n121 2.34304
R6634 VCC.n760 VCC.n746 2.34304
R6635 VCC.n633 VCC.n631 2.34304
R6636 VCC.n675 VCC.n673 2.34304
R6637 VCC.n1190 VCC.n1188 2.34304
R6638 VCC.n1232 VCC.n1230 2.34304
R6639 VCC.n1318 VCC.n1304 2.34304
R6640 VCC.n1869 VCC.n1855 2.34304
R6641 VCC.n1742 VCC.n1740 2.34304
R6642 VCC.n1784 VCC.n1782 2.34304
R6643 VCC.n2299 VCC.n2297 2.34304
R6644 VCC.n2341 VCC.n2339 2.34304
R6645 VCC.n2427 VCC.n2413 2.34304
R6646 VCC.n2978 VCC.n2964 2.34304
R6647 VCC.n2851 VCC.n2849 2.34304
R6648 VCC.n2893 VCC.n2891 2.34304
R6649 VCC.n3408 VCC.n3406 2.34304
R6650 VCC.n3450 VCC.n3448 2.34304
R6651 VCC.n3536 VCC.n3522 2.34304
R6652 VCC.n4087 VCC.n4073 2.34304
R6653 VCC.n3960 VCC.n3958 2.34304
R6654 VCC.n4002 VCC.n4000 2.34304
R6655 VCC.n4517 VCC.n4515 2.34304
R6656 VCC.n4559 VCC.n4557 2.34304
R6657 VCC.n4645 VCC.n4631 2.34304
R6658 VCC.n5196 VCC.n5182 2.34304
R6659 VCC.n5069 VCC.n5067 2.34304
R6660 VCC.n5111 VCC.n5109 2.34304
R6661 VCC.n5625 VCC.n5623 2.34304
R6662 VCC.n5667 VCC.n5665 2.34304
R6663 VCC.n5753 VCC.n5739 2.34304
R6664 VCC.n6303 VCC.n6289 2.34304
R6665 VCC.n6176 VCC.n6174 2.34304
R6666 VCC.n6218 VCC.n6216 2.34304
R6667 VCC.n6732 VCC.n6730 2.34304
R6668 VCC.n6774 VCC.n6772 2.34304
R6669 VCC.n6860 VCC.n6846 2.34304
R6670 VCC.n7410 VCC.n7396 2.34304
R6671 VCC.n7283 VCC.n7281 2.34304
R6672 VCC.n7325 VCC.n7323 2.34304
R6673 VCC.n7839 VCC.n7837 2.34304
R6674 VCC.n7881 VCC.n7879 2.34304
R6675 VCC.n7967 VCC.n7953 2.34304
R6676 VCC.n8390 VCC.n8388 2.34304
R6677 VCC.n8432 VCC.n8430 2.34304
R6678 VCC.n1662 VCC.n1107 2.29829
R6679 VCC.n3880 VCC.n3325 2.29829
R6680 VCC.n8682 VCC.n8681 2.29829
R6681 VCC.n8678 VCC.n8677 2.29829
R6682 VCC.n201 VCC.n183 2.28621
R6683 VCC.n326 VCC.n118 2.28621
R6684 VCC.n753 VCC.n735 2.28621
R6685 VCC.n878 VCC.n670 2.28621
R6686 VCC.n1435 VCC.n1227 2.28621
R6687 VCC.n1311 VCC.n1293 2.28621
R6688 VCC.n1862 VCC.n1844 2.28621
R6689 VCC.n1987 VCC.n1779 2.28621
R6690 VCC.n2544 VCC.n2336 2.28621
R6691 VCC.n2420 VCC.n2402 2.28621
R6692 VCC.n2971 VCC.n2953 2.28621
R6693 VCC.n3096 VCC.n2888 2.28621
R6694 VCC.n3653 VCC.n3445 2.28621
R6695 VCC.n3529 VCC.n3511 2.28621
R6696 VCC.n4080 VCC.n4062 2.28621
R6697 VCC.n4205 VCC.n3997 2.28621
R6698 VCC.n4762 VCC.n4554 2.28621
R6699 VCC.n4638 VCC.n4620 2.28621
R6700 VCC.n5189 VCC.n5171 2.28621
R6701 VCC.n5314 VCC.n5106 2.28621
R6702 VCC.n5870 VCC.n5662 2.28621
R6703 VCC.n5746 VCC.n5728 2.28621
R6704 VCC.n6296 VCC.n6278 2.28621
R6705 VCC.n6421 VCC.n6213 2.28621
R6706 VCC.n6977 VCC.n6769 2.28621
R6707 VCC.n6853 VCC.n6835 2.28621
R6708 VCC.n7403 VCC.n7385 2.28621
R6709 VCC.n7528 VCC.n7320 2.28621
R6710 VCC.n8084 VCC.n7876 2.28621
R6711 VCC.n7960 VCC.n7942 2.28621
R6712 VCC.n8448 VCC.n8427 2.28621
R6713 VCC.n130 VCC.n129 2.2505
R6714 VCC.n304 VCC.n133 2.2505
R6715 VCC.n277 VCC.n149 2.2505
R6716 VCC.n193 VCC.n190 2.2505
R6717 VCC.n186 VCC.n185 2.2505
R6718 VCC.n235 VCC.n234 2.2505
R6719 VCC.n69 VCC.n68 2.2505
R6720 VCC.n439 VCC.n72 2.2505
R6721 VCC.n404 VCC.n89 2.2505
R6722 VCC.n332 VCC.n319 2.2505
R6723 VCC.n116 VCC.n115 2.2505
R6724 VCC.n351 VCC.n349 2.2505
R6725 VCC.n539 VCC.n12 2.2505
R6726 VCC.n465 VCC.n59 2.2505
R6727 VCC.n488 VCC.n487 2.2505
R6728 VCC.n28 VCC.n26 2.2505
R6729 VCC.n533 VCC.n15 2.2505
R6730 VCC.n457 VCC.n64 2.2505
R6731 VCC.n682 VCC.n681 2.2505
R6732 VCC.n856 VCC.n685 2.2505
R6733 VCC.n829 VCC.n701 2.2505
R6734 VCC.n745 VCC.n742 2.2505
R6735 VCC.n738 VCC.n737 2.2505
R6736 VCC.n787 VCC.n786 2.2505
R6737 VCC.n621 VCC.n620 2.2505
R6738 VCC.n991 VCC.n624 2.2505
R6739 VCC.n956 VCC.n641 2.2505
R6740 VCC.n884 VCC.n871 2.2505
R6741 VCC.n668 VCC.n667 2.2505
R6742 VCC.n903 VCC.n901 2.2505
R6743 VCC.n1093 VCC.n1092 2.2505
R6744 VCC.n1085 VCC.n567 2.2505
R6745 VCC.n580 VCC.n578 2.2505
R6746 VCC.n1009 VCC.n616 2.2505
R6747 VCC.n1017 VCC.n611 2.2505
R6748 VCC.n1040 VCC.n1039 2.2505
R6749 VCC.n1639 VCC.n1638 2.2505
R6750 VCC.n1590 VCC.n1589 2.2505
R6751 VCC.n1120 VCC.n1118 2.2505
R6752 VCC.n1625 VCC.n1132 2.2505
R6753 VCC.n1575 VCC.n1574 2.2505
R6754 VCC.n1568 VCC.n1173 2.2505
R6755 VCC.n1178 VCC.n1177 2.2505
R6756 VCC.n1549 VCC.n1181 2.2505
R6757 VCC.n1513 VCC.n1198 2.2505
R6758 VCC.n1460 VCC.n1458 2.2505
R6759 VCC.n1225 VCC.n1224 2.2505
R6760 VCC.n1441 VCC.n1440 2.2505
R6761 VCC.n1240 VCC.n1239 2.2505
R6762 VCC.n1414 VCC.n1243 2.2505
R6763 VCC.n1387 VCC.n1259 2.2505
R6764 VCC.n1345 VCC.n1344 2.2505
R6765 VCC.n1296 VCC.n1295 2.2505
R6766 VCC.n1303 VCC.n1300 2.2505
R6767 VCC.n1791 VCC.n1790 2.2505
R6768 VCC.n1965 VCC.n1794 2.2505
R6769 VCC.n1938 VCC.n1810 2.2505
R6770 VCC.n1854 VCC.n1851 2.2505
R6771 VCC.n1847 VCC.n1846 2.2505
R6772 VCC.n1896 VCC.n1895 2.2505
R6773 VCC.n1730 VCC.n1729 2.2505
R6774 VCC.n2100 VCC.n1733 2.2505
R6775 VCC.n2065 VCC.n1750 2.2505
R6776 VCC.n1993 VCC.n1980 2.2505
R6777 VCC.n1777 VCC.n1776 2.2505
R6778 VCC.n2012 VCC.n2010 2.2505
R6779 VCC.n2202 VCC.n2201 2.2505
R6780 VCC.n2194 VCC.n1676 2.2505
R6781 VCC.n1689 VCC.n1687 2.2505
R6782 VCC.n2118 VCC.n1725 2.2505
R6783 VCC.n2126 VCC.n1720 2.2505
R6784 VCC.n2149 VCC.n2148 2.2505
R6785 VCC.n2748 VCC.n2747 2.2505
R6786 VCC.n2699 VCC.n2698 2.2505
R6787 VCC.n2229 VCC.n2227 2.2505
R6788 VCC.n2734 VCC.n2241 2.2505
R6789 VCC.n2684 VCC.n2683 2.2505
R6790 VCC.n2677 VCC.n2282 2.2505
R6791 VCC.n2287 VCC.n2286 2.2505
R6792 VCC.n2658 VCC.n2290 2.2505
R6793 VCC.n2622 VCC.n2307 2.2505
R6794 VCC.n2569 VCC.n2567 2.2505
R6795 VCC.n2334 VCC.n2333 2.2505
R6796 VCC.n2550 VCC.n2549 2.2505
R6797 VCC.n2349 VCC.n2348 2.2505
R6798 VCC.n2523 VCC.n2352 2.2505
R6799 VCC.n2496 VCC.n2368 2.2505
R6800 VCC.n2454 VCC.n2453 2.2505
R6801 VCC.n2405 VCC.n2404 2.2505
R6802 VCC.n2412 VCC.n2409 2.2505
R6803 VCC.n2900 VCC.n2899 2.2505
R6804 VCC.n3074 VCC.n2903 2.2505
R6805 VCC.n3047 VCC.n2919 2.2505
R6806 VCC.n2963 VCC.n2960 2.2505
R6807 VCC.n2956 VCC.n2955 2.2505
R6808 VCC.n3005 VCC.n3004 2.2505
R6809 VCC.n2839 VCC.n2838 2.2505
R6810 VCC.n3209 VCC.n2842 2.2505
R6811 VCC.n3174 VCC.n2859 2.2505
R6812 VCC.n3102 VCC.n3089 2.2505
R6813 VCC.n2886 VCC.n2885 2.2505
R6814 VCC.n3121 VCC.n3119 2.2505
R6815 VCC.n3311 VCC.n3310 2.2505
R6816 VCC.n3303 VCC.n2785 2.2505
R6817 VCC.n2798 VCC.n2796 2.2505
R6818 VCC.n3227 VCC.n2834 2.2505
R6819 VCC.n3235 VCC.n2829 2.2505
R6820 VCC.n3258 VCC.n3257 2.2505
R6821 VCC.n3857 VCC.n3856 2.2505
R6822 VCC.n3808 VCC.n3807 2.2505
R6823 VCC.n3338 VCC.n3336 2.2505
R6824 VCC.n3843 VCC.n3350 2.2505
R6825 VCC.n3793 VCC.n3792 2.2505
R6826 VCC.n3786 VCC.n3391 2.2505
R6827 VCC.n3396 VCC.n3395 2.2505
R6828 VCC.n3767 VCC.n3399 2.2505
R6829 VCC.n3731 VCC.n3416 2.2505
R6830 VCC.n3678 VCC.n3676 2.2505
R6831 VCC.n3443 VCC.n3442 2.2505
R6832 VCC.n3659 VCC.n3658 2.2505
R6833 VCC.n3458 VCC.n3457 2.2505
R6834 VCC.n3632 VCC.n3461 2.2505
R6835 VCC.n3605 VCC.n3477 2.2505
R6836 VCC.n3563 VCC.n3562 2.2505
R6837 VCC.n3514 VCC.n3513 2.2505
R6838 VCC.n3521 VCC.n3518 2.2505
R6839 VCC.n4009 VCC.n4008 2.2505
R6840 VCC.n4183 VCC.n4012 2.2505
R6841 VCC.n4156 VCC.n4028 2.2505
R6842 VCC.n4072 VCC.n4069 2.2505
R6843 VCC.n4065 VCC.n4064 2.2505
R6844 VCC.n4114 VCC.n4113 2.2505
R6845 VCC.n3948 VCC.n3947 2.2505
R6846 VCC.n4318 VCC.n3951 2.2505
R6847 VCC.n4283 VCC.n3968 2.2505
R6848 VCC.n4211 VCC.n4198 2.2505
R6849 VCC.n3995 VCC.n3994 2.2505
R6850 VCC.n4230 VCC.n4228 2.2505
R6851 VCC.n4420 VCC.n4419 2.2505
R6852 VCC.n4412 VCC.n3894 2.2505
R6853 VCC.n3907 VCC.n3905 2.2505
R6854 VCC.n4336 VCC.n3943 2.2505
R6855 VCC.n4344 VCC.n3938 2.2505
R6856 VCC.n4367 VCC.n4366 2.2505
R6857 VCC.n4966 VCC.n4965 2.2505
R6858 VCC.n4917 VCC.n4916 2.2505
R6859 VCC.n4447 VCC.n4445 2.2505
R6860 VCC.n4952 VCC.n4459 2.2505
R6861 VCC.n4902 VCC.n4901 2.2505
R6862 VCC.n4895 VCC.n4500 2.2505
R6863 VCC.n4505 VCC.n4504 2.2505
R6864 VCC.n4876 VCC.n4508 2.2505
R6865 VCC.n4840 VCC.n4525 2.2505
R6866 VCC.n4787 VCC.n4785 2.2505
R6867 VCC.n4552 VCC.n4551 2.2505
R6868 VCC.n4768 VCC.n4767 2.2505
R6869 VCC.n4567 VCC.n4566 2.2505
R6870 VCC.n4741 VCC.n4570 2.2505
R6871 VCC.n4714 VCC.n4586 2.2505
R6872 VCC.n4672 VCC.n4671 2.2505
R6873 VCC.n4623 VCC.n4622 2.2505
R6874 VCC.n4630 VCC.n4627 2.2505
R6875 VCC.n5118 VCC.n5117 2.2505
R6876 VCC.n5292 VCC.n5121 2.2505
R6877 VCC.n5265 VCC.n5137 2.2505
R6878 VCC.n5181 VCC.n5178 2.2505
R6879 VCC.n5174 VCC.n5173 2.2505
R6880 VCC.n5223 VCC.n5222 2.2505
R6881 VCC.n5057 VCC.n5056 2.2505
R6882 VCC.n5427 VCC.n5060 2.2505
R6883 VCC.n5392 VCC.n5077 2.2505
R6884 VCC.n5320 VCC.n5307 2.2505
R6885 VCC.n5104 VCC.n5103 2.2505
R6886 VCC.n5339 VCC.n5337 2.2505
R6887 VCC.n5529 VCC.n5528 2.2505
R6888 VCC.n5521 VCC.n5003 2.2505
R6889 VCC.n5016 VCC.n5014 2.2505
R6890 VCC.n5445 VCC.n5052 2.2505
R6891 VCC.n5453 VCC.n5047 2.2505
R6892 VCC.n5476 VCC.n5475 2.2505
R6893 VCC.n6074 VCC.n6073 2.2505
R6894 VCC.n6025 VCC.n6024 2.2505
R6895 VCC.n5555 VCC.n5553 2.2505
R6896 VCC.n6060 VCC.n5567 2.2505
R6897 VCC.n6010 VCC.n6009 2.2505
R6898 VCC.n6003 VCC.n5608 2.2505
R6899 VCC.n5613 VCC.n5612 2.2505
R6900 VCC.n5984 VCC.n5616 2.2505
R6901 VCC.n5948 VCC.n5633 2.2505
R6902 VCC.n5895 VCC.n5893 2.2505
R6903 VCC.n5660 VCC.n5659 2.2505
R6904 VCC.n5876 VCC.n5875 2.2505
R6905 VCC.n5675 VCC.n5674 2.2505
R6906 VCC.n5849 VCC.n5678 2.2505
R6907 VCC.n5822 VCC.n5694 2.2505
R6908 VCC.n5780 VCC.n5779 2.2505
R6909 VCC.n5731 VCC.n5730 2.2505
R6910 VCC.n5738 VCC.n5735 2.2505
R6911 VCC.n6225 VCC.n6224 2.2505
R6912 VCC.n6399 VCC.n6228 2.2505
R6913 VCC.n6372 VCC.n6244 2.2505
R6914 VCC.n6288 VCC.n6285 2.2505
R6915 VCC.n6281 VCC.n6280 2.2505
R6916 VCC.n6330 VCC.n6329 2.2505
R6917 VCC.n6164 VCC.n6163 2.2505
R6918 VCC.n6534 VCC.n6167 2.2505
R6919 VCC.n6499 VCC.n6184 2.2505
R6920 VCC.n6427 VCC.n6414 2.2505
R6921 VCC.n6211 VCC.n6210 2.2505
R6922 VCC.n6446 VCC.n6444 2.2505
R6923 VCC.n6636 VCC.n6635 2.2505
R6924 VCC.n6628 VCC.n6110 2.2505
R6925 VCC.n6123 VCC.n6121 2.2505
R6926 VCC.n6552 VCC.n6159 2.2505
R6927 VCC.n6560 VCC.n6154 2.2505
R6928 VCC.n6583 VCC.n6582 2.2505
R6929 VCC.n7181 VCC.n7180 2.2505
R6930 VCC.n7132 VCC.n7131 2.2505
R6931 VCC.n6662 VCC.n6660 2.2505
R6932 VCC.n7167 VCC.n6674 2.2505
R6933 VCC.n7117 VCC.n7116 2.2505
R6934 VCC.n7110 VCC.n6715 2.2505
R6935 VCC.n6720 VCC.n6719 2.2505
R6936 VCC.n7091 VCC.n6723 2.2505
R6937 VCC.n7055 VCC.n6740 2.2505
R6938 VCC.n7002 VCC.n7000 2.2505
R6939 VCC.n6767 VCC.n6766 2.2505
R6940 VCC.n6983 VCC.n6982 2.2505
R6941 VCC.n6782 VCC.n6781 2.2505
R6942 VCC.n6956 VCC.n6785 2.2505
R6943 VCC.n6929 VCC.n6801 2.2505
R6944 VCC.n6887 VCC.n6886 2.2505
R6945 VCC.n6838 VCC.n6837 2.2505
R6946 VCC.n6845 VCC.n6842 2.2505
R6947 VCC.n7332 VCC.n7331 2.2505
R6948 VCC.n7506 VCC.n7335 2.2505
R6949 VCC.n7479 VCC.n7351 2.2505
R6950 VCC.n7395 VCC.n7392 2.2505
R6951 VCC.n7388 VCC.n7387 2.2505
R6952 VCC.n7437 VCC.n7436 2.2505
R6953 VCC.n7271 VCC.n7270 2.2505
R6954 VCC.n7641 VCC.n7274 2.2505
R6955 VCC.n7606 VCC.n7291 2.2505
R6956 VCC.n7534 VCC.n7521 2.2505
R6957 VCC.n7318 VCC.n7317 2.2505
R6958 VCC.n7553 VCC.n7551 2.2505
R6959 VCC.n7743 VCC.n7742 2.2505
R6960 VCC.n7735 VCC.n7217 2.2505
R6961 VCC.n7230 VCC.n7228 2.2505
R6962 VCC.n7659 VCC.n7266 2.2505
R6963 VCC.n7667 VCC.n7261 2.2505
R6964 VCC.n7690 VCC.n7689 2.2505
R6965 VCC.n8288 VCC.n8287 2.2505
R6966 VCC.n8239 VCC.n8238 2.2505
R6967 VCC.n7769 VCC.n7767 2.2505
R6968 VCC.n8274 VCC.n7781 2.2505
R6969 VCC.n8224 VCC.n8223 2.2505
R6970 VCC.n8217 VCC.n7822 2.2505
R6971 VCC.n7827 VCC.n7826 2.2505
R6972 VCC.n8198 VCC.n7830 2.2505
R6973 VCC.n8162 VCC.n7847 2.2505
R6974 VCC.n8109 VCC.n8107 2.2505
R6975 VCC.n7874 VCC.n7873 2.2505
R6976 VCC.n8090 VCC.n8089 2.2505
R6977 VCC.n7889 VCC.n7888 2.2505
R6978 VCC.n8063 VCC.n7892 2.2505
R6979 VCC.n8036 VCC.n7908 2.2505
R6980 VCC.n7994 VCC.n7993 2.2505
R6981 VCC.n7945 VCC.n7944 2.2505
R6982 VCC.n7952 VCC.n7949 2.2505
R6983 VCC.n8378 VCC.n8377 2.2505
R6984 VCC.n8561 VCC.n8381 2.2505
R6985 VCC.n8526 VCC.n8398 2.2505
R6986 VCC.n8454 VCC.n8441 2.2505
R6987 VCC.n8425 VCC.n8424 2.2505
R6988 VCC.n8473 VCC.n8471 2.2505
R6989 VCC.n8663 VCC.n8662 2.2505
R6990 VCC.n8655 VCC.n8324 2.2505
R6991 VCC.n8337 VCC.n8335 2.2505
R6992 VCC.n8579 VCC.n8373 2.2505
R6993 VCC.n8587 VCC.n8368 2.2505
R6994 VCC.n8610 VCC.n8609 2.2505
R6995 VCC.n8677 VCC 2.24163
R6996 VCC.n2216 VCC.n1662 2.21741
R6997 VCC.n4434 VCC.n3880 2.21741
R6998 VCC.n8681 VCC.n8680 2.21741
R6999 VCC.n264 VCC.n263 2.10336
R7000 VCC.n386 VCC.n385 2.10336
R7001 VCC.n816 VCC.n815 2.10336
R7002 VCC.n938 VCC.n937 2.10336
R7003 VCC.n1495 VCC.n1494 2.10336
R7004 VCC.n1374 VCC.n1373 2.10336
R7005 VCC.n1925 VCC.n1924 2.10336
R7006 VCC.n2047 VCC.n2046 2.10336
R7007 VCC.n2604 VCC.n2603 2.10336
R7008 VCC.n2483 VCC.n2482 2.10336
R7009 VCC.n3034 VCC.n3033 2.10336
R7010 VCC.n3156 VCC.n3155 2.10336
R7011 VCC.n3713 VCC.n3712 2.10336
R7012 VCC.n3592 VCC.n3591 2.10336
R7013 VCC.n4143 VCC.n4142 2.10336
R7014 VCC.n4265 VCC.n4264 2.10336
R7015 VCC.n4822 VCC.n4821 2.10336
R7016 VCC.n4701 VCC.n4700 2.10336
R7017 VCC.n5252 VCC.n5251 2.10336
R7018 VCC.n5374 VCC.n5373 2.10336
R7019 VCC.n5930 VCC.n5929 2.10336
R7020 VCC.n5809 VCC.n5808 2.10336
R7021 VCC.n6359 VCC.n6358 2.10336
R7022 VCC.n6481 VCC.n6480 2.10336
R7023 VCC.n7037 VCC.n7036 2.10336
R7024 VCC.n6916 VCC.n6915 2.10336
R7025 VCC.n7466 VCC.n7465 2.10336
R7026 VCC.n7588 VCC.n7587 2.10336
R7027 VCC.n8144 VCC.n8143 2.10336
R7028 VCC.n8023 VCC.n8022 2.10336
R7029 VCC.n8508 VCC.n8507 2.10336
R7030 VCC.n264 VCC.n155 2.01193
R7031 VCC.n385 VCC.n384 2.01193
R7032 VCC.n816 VCC.n707 2.01193
R7033 VCC.n937 VCC.n936 2.01193
R7034 VCC.n1494 VCC.n1493 2.01193
R7035 VCC.n1374 VCC.n1265 2.01193
R7036 VCC.n1925 VCC.n1816 2.01193
R7037 VCC.n2046 VCC.n2045 2.01193
R7038 VCC.n2603 VCC.n2602 2.01193
R7039 VCC.n2483 VCC.n2374 2.01193
R7040 VCC.n3034 VCC.n2925 2.01193
R7041 VCC.n3155 VCC.n3154 2.01193
R7042 VCC.n3712 VCC.n3711 2.01193
R7043 VCC.n3592 VCC.n3483 2.01193
R7044 VCC.n4143 VCC.n4034 2.01193
R7045 VCC.n4264 VCC.n4263 2.01193
R7046 VCC.n4821 VCC.n4820 2.01193
R7047 VCC.n4701 VCC.n4592 2.01193
R7048 VCC.n5252 VCC.n5143 2.01193
R7049 VCC.n5373 VCC.n5372 2.01193
R7050 VCC.n5929 VCC.n5928 2.01193
R7051 VCC.n5809 VCC.n5700 2.01193
R7052 VCC.n6359 VCC.n6250 2.01193
R7053 VCC.n6480 VCC.n6479 2.01193
R7054 VCC.n7036 VCC.n7035 2.01193
R7055 VCC.n6916 VCC.n6807 2.01193
R7056 VCC.n7466 VCC.n7357 2.01193
R7057 VCC.n7587 VCC.n7586 2.01193
R7058 VCC.n8143 VCC.n8142 2.01193
R7059 VCC.n8023 VCC.n7914 2.01193
R7060 VCC.n8507 VCC.n8506 2.01193
R7061 VCC.n550 VCC.n549 2.00996
R7062 VCC.n1104 VCC.n1103 2.00996
R7063 VCC.n1658 VCC.n1657 2.00996
R7064 VCC.n2213 VCC.n2212 2.00996
R7065 VCC.n2767 VCC.n2766 2.00996
R7066 VCC.n3322 VCC.n3321 2.00996
R7067 VCC.n3876 VCC.n3875 2.00996
R7068 VCC.n4431 VCC.n4430 2.00996
R7069 VCC.n4985 VCC.n4984 2.00996
R7070 VCC.n5540 VCC.n5539 2.00996
R7071 VCC.n6093 VCC.n6092 2.00996
R7072 VCC.n6647 VCC.n6646 2.00996
R7073 VCC.n7200 VCC.n7199 2.00996
R7074 VCC.n7754 VCC.n7753 2.00996
R7075 VCC.n8307 VCC.n8306 2.00996
R7076 VCC.n8674 VCC.n8673 2.00996
R7077 VCC VCC.n2216 1.98947
R7078 VCC.n8680 VCC 1.98947
R7079 VCC.n451 VCC.n65 1.98102
R7080 VCC.n1003 VCC.n617 1.98102
R7081 VCC.n2112 VCC.n1726 1.98102
R7082 VCC.n3221 VCC.n2835 1.98102
R7083 VCC.n4330 VCC.n3944 1.98102
R7084 VCC.n5439 VCC.n5053 1.98102
R7085 VCC.n6546 VCC.n6160 1.98102
R7086 VCC.n7653 VCC.n7267 1.98102
R7087 VCC.n8573 VCC.n8374 1.98102
R7088 VCC.n1561 VCC.n1174 1.98071
R7089 VCC.n2670 VCC.n2283 1.98071
R7090 VCC.n3779 VCC.n3392 1.98071
R7091 VCC.n4888 VCC.n4501 1.98071
R7092 VCC.n5996 VCC.n5609 1.98071
R7093 VCC.n7103 VCC.n6716 1.98071
R7094 VCC.n8210 VCC.n7823 1.98071
R7095 VCC.n1107 VCC 1.87918
R7096 VCC.n3325 VCC 1.87918
R7097 VCC VCC.n8682 1.87918
R7098 VCC VCC.n8678 1.87918
R7099 VCC.n229 VCC.n228 1.82742
R7100 VCC.n268 VCC.n142 1.82742
R7101 VCC.n361 VCC.n360 1.82742
R7102 VCC.n396 VCC.n395 1.82742
R7103 VCC.n781 VCC.n780 1.82742
R7104 VCC.n820 VCC.n694 1.82742
R7105 VCC.n913 VCC.n912 1.82742
R7106 VCC.n948 VCC.n947 1.82742
R7107 VCC.n1470 VCC.n1469 1.82742
R7108 VCC.n1505 VCC.n1504 1.82742
R7109 VCC.n1339 VCC.n1338 1.82742
R7110 VCC.n1378 VCC.n1252 1.82742
R7111 VCC.n1890 VCC.n1889 1.82742
R7112 VCC.n1929 VCC.n1803 1.82742
R7113 VCC.n2022 VCC.n2021 1.82742
R7114 VCC.n2057 VCC.n2056 1.82742
R7115 VCC.n2579 VCC.n2578 1.82742
R7116 VCC.n2614 VCC.n2613 1.82742
R7117 VCC.n2448 VCC.n2447 1.82742
R7118 VCC.n2487 VCC.n2361 1.82742
R7119 VCC.n2999 VCC.n2998 1.82742
R7120 VCC.n3038 VCC.n2912 1.82742
R7121 VCC.n3131 VCC.n3130 1.82742
R7122 VCC.n3166 VCC.n3165 1.82742
R7123 VCC.n3688 VCC.n3687 1.82742
R7124 VCC.n3723 VCC.n3722 1.82742
R7125 VCC.n3557 VCC.n3556 1.82742
R7126 VCC.n3596 VCC.n3470 1.82742
R7127 VCC.n4108 VCC.n4107 1.82742
R7128 VCC.n4147 VCC.n4021 1.82742
R7129 VCC.n4240 VCC.n4239 1.82742
R7130 VCC.n4275 VCC.n4274 1.82742
R7131 VCC.n4797 VCC.n4796 1.82742
R7132 VCC.n4832 VCC.n4831 1.82742
R7133 VCC.n4666 VCC.n4665 1.82742
R7134 VCC.n4705 VCC.n4579 1.82742
R7135 VCC.n5217 VCC.n5216 1.82742
R7136 VCC.n5256 VCC.n5130 1.82742
R7137 VCC.n5349 VCC.n5348 1.82742
R7138 VCC.n5384 VCC.n5383 1.82742
R7139 VCC.n5905 VCC.n5904 1.82742
R7140 VCC.n5940 VCC.n5939 1.82742
R7141 VCC.n5774 VCC.n5773 1.82742
R7142 VCC.n5813 VCC.n5687 1.82742
R7143 VCC.n6324 VCC.n6323 1.82742
R7144 VCC.n6363 VCC.n6237 1.82742
R7145 VCC.n6456 VCC.n6455 1.82742
R7146 VCC.n6491 VCC.n6490 1.82742
R7147 VCC.n7012 VCC.n7011 1.82742
R7148 VCC.n7047 VCC.n7046 1.82742
R7149 VCC.n6881 VCC.n6880 1.82742
R7150 VCC.n6920 VCC.n6794 1.82742
R7151 VCC.n7431 VCC.n7430 1.82742
R7152 VCC.n7470 VCC.n7344 1.82742
R7153 VCC.n7563 VCC.n7562 1.82742
R7154 VCC.n7598 VCC.n7597 1.82742
R7155 VCC.n8119 VCC.n8118 1.82742
R7156 VCC.n8154 VCC.n8153 1.82742
R7157 VCC.n7988 VCC.n7987 1.82742
R7158 VCC.n8027 VCC.n7901 1.82742
R7159 VCC.n8483 VCC.n8482 1.82742
R7160 VCC.n8518 VCC.n8517 1.82742
R7161 VCC VCC.n4434 1.67697
R7162 VCC.n492 VCC.n42 1.62907
R7163 VCC.n524 VCC.n23 1.62907
R7164 VCC.n1044 VCC.n594 1.62907
R7165 VCC.n1076 VCC.n575 1.62907
R7166 VCC.n1586 VCC.n1162 1.62907
R7167 VCC.n1622 VCC.n1142 1.62907
R7168 VCC.n2153 VCC.n1703 1.62907
R7169 VCC.n2185 VCC.n1684 1.62907
R7170 VCC.n2695 VCC.n2271 1.62907
R7171 VCC.n2731 VCC.n2251 1.62907
R7172 VCC.n3262 VCC.n2812 1.62907
R7173 VCC.n3294 VCC.n2793 1.62907
R7174 VCC.n3804 VCC.n3380 1.62907
R7175 VCC.n3840 VCC.n3360 1.62907
R7176 VCC.n4371 VCC.n3921 1.62907
R7177 VCC.n4403 VCC.n3902 1.62907
R7178 VCC.n4913 VCC.n4489 1.62907
R7179 VCC.n4949 VCC.n4469 1.62907
R7180 VCC.n5480 VCC.n5030 1.62907
R7181 VCC.n5512 VCC.n5011 1.62907
R7182 VCC.n6021 VCC.n5597 1.62907
R7183 VCC.n6057 VCC.n5577 1.62907
R7184 VCC.n6587 VCC.n6137 1.62907
R7185 VCC.n6619 VCC.n6118 1.62907
R7186 VCC.n7128 VCC.n6704 1.62907
R7187 VCC.n7164 VCC.n6684 1.62907
R7188 VCC.n7694 VCC.n7244 1.62907
R7189 VCC.n7726 VCC.n7225 1.62907
R7190 VCC.n8235 VCC.n7811 1.62907
R7191 VCC.n8271 VCC.n7791 1.62907
R7192 VCC.n8614 VCC.n8351 1.62907
R7193 VCC.n8646 VCC.n8332 1.62907
R7194 VCC.n468 VCC.n57 1.55479
R7195 VCC.n1020 VCC.n609 1.55479
R7196 VCC.n1577 VCC.n1165 1.55479
R7197 VCC.n2129 VCC.n1718 1.55479
R7198 VCC.n2686 VCC.n2274 1.55479
R7199 VCC.n3238 VCC.n2827 1.55479
R7200 VCC.n3795 VCC.n3383 1.55479
R7201 VCC.n4347 VCC.n3936 1.55479
R7202 VCC.n4904 VCC.n4492 1.55479
R7203 VCC.n5456 VCC.n5045 1.55479
R7204 VCC.n6012 VCC.n5600 1.55479
R7205 VCC.n6563 VCC.n6152 1.55479
R7206 VCC.n7119 VCC.n6707 1.55479
R7207 VCC.n7670 VCC.n7259 1.55479
R7208 VCC.n8226 VCC.n7814 1.55479
R7209 VCC.n8590 VCC.n8366 1.55479
R7210 VCC.n253 VCC.n252 1.5005
R7211 VCC.n805 VCC.n804 1.5005
R7212 VCC.n1363 VCC.n1362 1.5005
R7213 VCC.n1914 VCC.n1913 1.5005
R7214 VCC.n2472 VCC.n2471 1.5005
R7215 VCC.n3023 VCC.n3022 1.5005
R7216 VCC.n3581 VCC.n3580 1.5005
R7217 VCC.n4132 VCC.n4131 1.5005
R7218 VCC.n4690 VCC.n4689 1.5005
R7219 VCC.n5241 VCC.n5240 1.5005
R7220 VCC.n5798 VCC.n5797 1.5005
R7221 VCC.n6348 VCC.n6347 1.5005
R7222 VCC.n6905 VCC.n6904 1.5005
R7223 VCC.n7455 VCC.n7454 1.5005
R7224 VCC.n8012 VCC.n8011 1.5005
R7225 VCC.n178 VCC.n169 1.46336
R7226 VCC.n270 VCC.n151 1.46336
R7227 VCC.n364 VCC.n106 1.46336
R7228 VCC.n392 VCC.n91 1.46336
R7229 VCC.n530 VCC.n7 1.46336
R7230 VCC.n730 VCC.n721 1.46336
R7231 VCC.n822 VCC.n703 1.46336
R7232 VCC.n916 VCC.n658 1.46336
R7233 VCC.n944 VCC.n643 1.46336
R7234 VCC.n1082 VCC.n561 1.46336
R7235 VCC.n1123 VCC.n1117 1.46336
R7236 VCC.n1473 VCC.n1215 1.46336
R7237 VCC.n1501 VCC.n1200 1.46336
R7238 VCC.n1288 VCC.n1279 1.46336
R7239 VCC.n1380 VCC.n1261 1.46336
R7240 VCC.n1839 VCC.n1830 1.46336
R7241 VCC.n1931 VCC.n1812 1.46336
R7242 VCC.n2025 VCC.n1767 1.46336
R7243 VCC.n2053 VCC.n1752 1.46336
R7244 VCC.n2191 VCC.n1670 1.46336
R7245 VCC.n2232 VCC.n2226 1.46336
R7246 VCC.n2582 VCC.n2324 1.46336
R7247 VCC.n2610 VCC.n2309 1.46336
R7248 VCC.n2397 VCC.n2388 1.46336
R7249 VCC.n2489 VCC.n2370 1.46336
R7250 VCC.n2948 VCC.n2939 1.46336
R7251 VCC.n3040 VCC.n2921 1.46336
R7252 VCC.n3134 VCC.n2876 1.46336
R7253 VCC.n3162 VCC.n2861 1.46336
R7254 VCC.n3300 VCC.n2779 1.46336
R7255 VCC.n3341 VCC.n3335 1.46336
R7256 VCC.n3691 VCC.n3433 1.46336
R7257 VCC.n3719 VCC.n3418 1.46336
R7258 VCC.n3506 VCC.n3497 1.46336
R7259 VCC.n3598 VCC.n3479 1.46336
R7260 VCC.n4057 VCC.n4048 1.46336
R7261 VCC.n4149 VCC.n4030 1.46336
R7262 VCC.n4243 VCC.n3985 1.46336
R7263 VCC.n4271 VCC.n3970 1.46336
R7264 VCC.n4409 VCC.n3888 1.46336
R7265 VCC.n4450 VCC.n4444 1.46336
R7266 VCC.n4800 VCC.n4542 1.46336
R7267 VCC.n4828 VCC.n4527 1.46336
R7268 VCC.n4615 VCC.n4606 1.46336
R7269 VCC.n4707 VCC.n4588 1.46336
R7270 VCC.n5166 VCC.n5157 1.46336
R7271 VCC.n5258 VCC.n5139 1.46336
R7272 VCC.n5352 VCC.n5094 1.46336
R7273 VCC.n5380 VCC.n5079 1.46336
R7274 VCC.n5518 VCC.n4997 1.46336
R7275 VCC.n5558 VCC.n5552 1.46336
R7276 VCC.n5908 VCC.n5650 1.46336
R7277 VCC.n5936 VCC.n5635 1.46336
R7278 VCC.n5723 VCC.n5714 1.46336
R7279 VCC.n5815 VCC.n5696 1.46336
R7280 VCC.n6273 VCC.n6264 1.46336
R7281 VCC.n6365 VCC.n6246 1.46336
R7282 VCC.n6459 VCC.n6201 1.46336
R7283 VCC.n6487 VCC.n6186 1.46336
R7284 VCC.n6625 VCC.n6104 1.46336
R7285 VCC.n6665 VCC.n6659 1.46336
R7286 VCC.n7015 VCC.n6757 1.46336
R7287 VCC.n7043 VCC.n6742 1.46336
R7288 VCC.n6830 VCC.n6821 1.46336
R7289 VCC.n6922 VCC.n6803 1.46336
R7290 VCC.n7380 VCC.n7371 1.46336
R7291 VCC.n7472 VCC.n7353 1.46336
R7292 VCC.n7566 VCC.n7308 1.46336
R7293 VCC.n7594 VCC.n7293 1.46336
R7294 VCC.n7732 VCC.n7211 1.46336
R7295 VCC.n7772 VCC.n7766 1.46336
R7296 VCC.n8122 VCC.n7864 1.46336
R7297 VCC.n8150 VCC.n7849 1.46336
R7298 VCC.n7937 VCC.n7928 1.46336
R7299 VCC.n8029 VCC.n7910 1.46336
R7300 VCC.n8486 VCC.n8415 1.46336
R7301 VCC.n8514 VCC.n8400 1.46336
R7302 VCC.n8652 VCC.n8318 1.46336
R7303 VCC.n476 VCC.n43 1.37193
R7304 VCC.n491 VCC.n39 1.37193
R7305 VCC.n498 VCC.n24 1.37193
R7306 VCC.n515 VCC.n25 1.37193
R7307 VCC.n1028 VCC.n595 1.37193
R7308 VCC.n1043 VCC.n591 1.37193
R7309 VCC.n1050 VCC.n576 1.37193
R7310 VCC.n1067 VCC.n577 1.37193
R7311 VCC.n1594 VCC.n1593 1.37193
R7312 VCC.n1160 VCC.n1145 1.37193
R7313 VCC.n1617 VCC.n1135 1.37193
R7314 VCC.n1141 VCC.n1140 1.37193
R7315 VCC.n2137 VCC.n1704 1.37193
R7316 VCC.n2152 VCC.n1700 1.37193
R7317 VCC.n2159 VCC.n1685 1.37193
R7318 VCC.n2176 VCC.n1686 1.37193
R7319 VCC.n2703 VCC.n2702 1.37193
R7320 VCC.n2269 VCC.n2254 1.37193
R7321 VCC.n2726 VCC.n2244 1.37193
R7322 VCC.n2250 VCC.n2249 1.37193
R7323 VCC.n3246 VCC.n2813 1.37193
R7324 VCC.n3261 VCC.n2809 1.37193
R7325 VCC.n3268 VCC.n2794 1.37193
R7326 VCC.n3285 VCC.n2795 1.37193
R7327 VCC.n3812 VCC.n3811 1.37193
R7328 VCC.n3378 VCC.n3363 1.37193
R7329 VCC.n3835 VCC.n3353 1.37193
R7330 VCC.n3359 VCC.n3358 1.37193
R7331 VCC.n4355 VCC.n3922 1.37193
R7332 VCC.n4370 VCC.n3918 1.37193
R7333 VCC.n4377 VCC.n3903 1.37193
R7334 VCC.n4394 VCC.n3904 1.37193
R7335 VCC.n4921 VCC.n4920 1.37193
R7336 VCC.n4487 VCC.n4472 1.37193
R7337 VCC.n4944 VCC.n4462 1.37193
R7338 VCC.n4468 VCC.n4467 1.37193
R7339 VCC.n5464 VCC.n5031 1.37193
R7340 VCC.n5479 VCC.n5027 1.37193
R7341 VCC.n5486 VCC.n5012 1.37193
R7342 VCC.n5503 VCC.n5013 1.37193
R7343 VCC.n6029 VCC.n6028 1.37193
R7344 VCC.n5595 VCC.n5580 1.37193
R7345 VCC.n6052 VCC.n5570 1.37193
R7346 VCC.n5576 VCC.n5575 1.37193
R7347 VCC.n6571 VCC.n6138 1.37193
R7348 VCC.n6586 VCC.n6134 1.37193
R7349 VCC.n6593 VCC.n6119 1.37193
R7350 VCC.n6610 VCC.n6120 1.37193
R7351 VCC.n7136 VCC.n7135 1.37193
R7352 VCC.n6702 VCC.n6687 1.37193
R7353 VCC.n7159 VCC.n6677 1.37193
R7354 VCC.n6683 VCC.n6682 1.37193
R7355 VCC.n7678 VCC.n7245 1.37193
R7356 VCC.n7693 VCC.n7241 1.37193
R7357 VCC.n7700 VCC.n7226 1.37193
R7358 VCC.n7717 VCC.n7227 1.37193
R7359 VCC.n8243 VCC.n8242 1.37193
R7360 VCC.n7809 VCC.n7794 1.37193
R7361 VCC.n8266 VCC.n7784 1.37193
R7362 VCC.n7790 VCC.n7789 1.37193
R7363 VCC.n8598 VCC.n8352 1.37193
R7364 VCC.n8613 VCC.n8348 1.37193
R7365 VCC.n8620 VCC.n8333 1.37193
R7366 VCC.n8637 VCC.n8334 1.37193
R7367 VCC.n224 VCC.n223 1.2805
R7368 VCC.n287 VCC.n286 1.2805
R7369 VCC.n341 VCC.n339 1.2805
R7370 VCC.n415 VCC.n413 1.2805
R7371 VCC.n776 VCC.n775 1.2805
R7372 VCC.n839 VCC.n838 1.2805
R7373 VCC.n893 VCC.n891 1.2805
R7374 VCC.n967 VCC.n965 1.2805
R7375 VCC.n1450 VCC.n1448 1.2805
R7376 VCC.n1524 VCC.n1522 1.2805
R7377 VCC.n1334 VCC.n1333 1.2805
R7378 VCC.n1397 VCC.n1396 1.2805
R7379 VCC.n1885 VCC.n1884 1.2805
R7380 VCC.n1948 VCC.n1947 1.2805
R7381 VCC.n2002 VCC.n2000 1.2805
R7382 VCC.n2076 VCC.n2074 1.2805
R7383 VCC.n2559 VCC.n2557 1.2805
R7384 VCC.n2633 VCC.n2631 1.2805
R7385 VCC.n2443 VCC.n2442 1.2805
R7386 VCC.n2506 VCC.n2505 1.2805
R7387 VCC.n2994 VCC.n2993 1.2805
R7388 VCC.n3057 VCC.n3056 1.2805
R7389 VCC.n3111 VCC.n3109 1.2805
R7390 VCC.n3185 VCC.n3183 1.2805
R7391 VCC.n3668 VCC.n3666 1.2805
R7392 VCC.n3742 VCC.n3740 1.2805
R7393 VCC.n3552 VCC.n3551 1.2805
R7394 VCC.n3615 VCC.n3614 1.2805
R7395 VCC.n4103 VCC.n4102 1.2805
R7396 VCC.n4166 VCC.n4165 1.2805
R7397 VCC.n4220 VCC.n4218 1.2805
R7398 VCC.n4294 VCC.n4292 1.2805
R7399 VCC.n4777 VCC.n4775 1.2805
R7400 VCC.n4851 VCC.n4849 1.2805
R7401 VCC.n4661 VCC.n4660 1.2805
R7402 VCC.n4724 VCC.n4723 1.2805
R7403 VCC.n5212 VCC.n5211 1.2805
R7404 VCC.n5275 VCC.n5274 1.2805
R7405 VCC.n5329 VCC.n5327 1.2805
R7406 VCC.n5403 VCC.n5401 1.2805
R7407 VCC.n5885 VCC.n5883 1.2805
R7408 VCC.n5959 VCC.n5957 1.2805
R7409 VCC.n5769 VCC.n5768 1.2805
R7410 VCC.n5832 VCC.n5831 1.2805
R7411 VCC.n6319 VCC.n6318 1.2805
R7412 VCC.n6382 VCC.n6381 1.2805
R7413 VCC.n6436 VCC.n6434 1.2805
R7414 VCC.n6510 VCC.n6508 1.2805
R7415 VCC.n6992 VCC.n6990 1.2805
R7416 VCC.n7066 VCC.n7064 1.2805
R7417 VCC.n6876 VCC.n6875 1.2805
R7418 VCC.n6939 VCC.n6938 1.2805
R7419 VCC.n7426 VCC.n7425 1.2805
R7420 VCC.n7489 VCC.n7488 1.2805
R7421 VCC.n7543 VCC.n7541 1.2805
R7422 VCC.n7617 VCC.n7615 1.2805
R7423 VCC.n8099 VCC.n8097 1.2805
R7424 VCC.n8173 VCC.n8171 1.2805
R7425 VCC.n7983 VCC.n7982 1.2805
R7426 VCC.n8046 VCC.n8045 1.2805
R7427 VCC.n8463 VCC.n8461 1.2805
R7428 VCC.n8537 VCC.n8535 1.2805
R7429 VCC.n475 VCC.n54 1.18907
R7430 VCC.n529 VCC.n20 1.18907
R7431 VCC.n1027 VCC.n606 1.18907
R7432 VCC.n1081 VCC.n572 1.18907
R7433 VCC.n1578 VCC.n1159 1.18907
R7434 VCC.n1649 VCC.n1116 1.18907
R7435 VCC.n2136 VCC.n1715 1.18907
R7436 VCC.n2190 VCC.n1681 1.18907
R7437 VCC.n2687 VCC.n2268 1.18907
R7438 VCC.n2758 VCC.n2225 1.18907
R7439 VCC.n3245 VCC.n2824 1.18907
R7440 VCC.n3299 VCC.n2790 1.18907
R7441 VCC.n3796 VCC.n3377 1.18907
R7442 VCC.n3867 VCC.n3334 1.18907
R7443 VCC.n4354 VCC.n3933 1.18907
R7444 VCC.n4408 VCC.n3899 1.18907
R7445 VCC.n4905 VCC.n4486 1.18907
R7446 VCC.n4976 VCC.n4443 1.18907
R7447 VCC.n5463 VCC.n5042 1.18907
R7448 VCC.n5517 VCC.n5008 1.18907
R7449 VCC.n6013 VCC.n5594 1.18907
R7450 VCC.n6084 VCC.n5551 1.18907
R7451 VCC.n6570 VCC.n6149 1.18907
R7452 VCC.n6624 VCC.n6115 1.18907
R7453 VCC.n7120 VCC.n6701 1.18907
R7454 VCC.n7191 VCC.n6658 1.18907
R7455 VCC.n7677 VCC.n7256 1.18907
R7456 VCC.n7731 VCC.n7222 1.18907
R7457 VCC.n8227 VCC.n7808 1.18907
R7458 VCC.n8298 VCC.n7765 1.18907
R7459 VCC.n8597 VCC.n8363 1.18907
R7460 VCC.n8651 VCC.n8329 1.18907
R7461 VCC.n1 VCC.n0 1.13717
R7462 VCC.n189 VCC.n188 1.13717
R7463 VCC.n187 VCC.n173 1.13717
R7464 VCC.n244 VCC.n243 1.13717
R7465 VCC.n164 VCC.n147 1.13717
R7466 VCC.n132 VCC.n131 1.13717
R7467 VCC.n128 VCC.n127 1.13717
R7468 VCC.n316 VCC.n126 1.13717
R7469 VCC.n346 VCC.n345 1.13717
R7470 VCC.n370 VCC.n369 1.13717
R7471 VCC.n373 VCC.n87 1.13717
R7472 VCC.n71 VCC.n70 1.13717
R7473 VCC.n67 VCC.n66 1.13717
R7474 VCC.n63 VCC.n62 1.13717
R7475 VCC.n61 VCC.n49 1.13717
R7476 VCC.n484 VCC.n483 1.13717
R7477 VCC.n34 VCC.n30 1.13717
R7478 VCC.n14 VCC.n13 1.13717
R7479 VCC.n741 VCC.n740 1.13717
R7480 VCC.n739 VCC.n725 1.13717
R7481 VCC.n796 VCC.n795 1.13717
R7482 VCC.n716 VCC.n699 1.13717
R7483 VCC.n684 VCC.n683 1.13717
R7484 VCC.n680 VCC.n679 1.13717
R7485 VCC.n868 VCC.n678 1.13717
R7486 VCC.n898 VCC.n897 1.13717
R7487 VCC.n922 VCC.n921 1.13717
R7488 VCC.n925 VCC.n639 1.13717
R7489 VCC.n623 VCC.n622 1.13717
R7490 VCC.n619 VCC.n618 1.13717
R7491 VCC.n615 VCC.n614 1.13717
R7492 VCC.n613 VCC.n601 1.13717
R7493 VCC.n1036 VCC.n1035 1.13717
R7494 VCC.n586 VCC.n582 1.13717
R7495 VCC.n566 VCC.n565 1.13717
R7496 VCC.n555 VCC.n554 1.13717
R7497 VCC.n1299 VCC.n1298 1.13717
R7498 VCC.n1297 VCC.n1283 1.13717
R7499 VCC.n1354 VCC.n1353 1.13717
R7500 VCC.n1274 VCC.n1257 1.13717
R7501 VCC.n1242 VCC.n1241 1.13717
R7502 VCC.n1238 VCC.n1237 1.13717
R7503 VCC.n1426 VCC.n1236 1.13717
R7504 VCC.n1170 VCC.n1154 1.13717
R7505 VCC.n1602 VCC.n1601 1.13717
R7506 VCC.n1609 VCC.n1130 1.13717
R7507 VCC.n1127 VCC.n1126 1.13717
R7508 VCC.n1109 VCC.n1108 1.13717
R7509 VCC.n1172 VCC.n1171 1.13717
R7510 VCC.n1455 VCC.n1454 1.13717
R7511 VCC.n1479 VCC.n1478 1.13717
R7512 VCC.n1482 VCC.n1196 1.13717
R7513 VCC.n1180 VCC.n1179 1.13717
R7514 VCC.n1176 VCC.n1175 1.13717
R7515 VCC.n1850 VCC.n1849 1.13717
R7516 VCC.n1848 VCC.n1834 1.13717
R7517 VCC.n1905 VCC.n1904 1.13717
R7518 VCC.n1825 VCC.n1808 1.13717
R7519 VCC.n1793 VCC.n1792 1.13717
R7520 VCC.n1789 VCC.n1788 1.13717
R7521 VCC.n1977 VCC.n1787 1.13717
R7522 VCC.n2007 VCC.n2006 1.13717
R7523 VCC.n2031 VCC.n2030 1.13717
R7524 VCC.n2034 VCC.n1748 1.13717
R7525 VCC.n1732 VCC.n1731 1.13717
R7526 VCC.n1728 VCC.n1727 1.13717
R7527 VCC.n1724 VCC.n1723 1.13717
R7528 VCC.n1722 VCC.n1710 1.13717
R7529 VCC.n2145 VCC.n2144 1.13717
R7530 VCC.n1695 VCC.n1691 1.13717
R7531 VCC.n1675 VCC.n1674 1.13717
R7532 VCC.n1664 VCC.n1663 1.13717
R7533 VCC.n2408 VCC.n2407 1.13717
R7534 VCC.n2406 VCC.n2392 1.13717
R7535 VCC.n2463 VCC.n2462 1.13717
R7536 VCC.n2383 VCC.n2366 1.13717
R7537 VCC.n2351 VCC.n2350 1.13717
R7538 VCC.n2347 VCC.n2346 1.13717
R7539 VCC.n2535 VCC.n2345 1.13717
R7540 VCC.n2279 VCC.n2263 1.13717
R7541 VCC.n2711 VCC.n2710 1.13717
R7542 VCC.n2718 VCC.n2239 1.13717
R7543 VCC.n2236 VCC.n2235 1.13717
R7544 VCC.n2218 VCC.n2217 1.13717
R7545 VCC.n2281 VCC.n2280 1.13717
R7546 VCC.n2564 VCC.n2563 1.13717
R7547 VCC.n2588 VCC.n2587 1.13717
R7548 VCC.n2591 VCC.n2305 1.13717
R7549 VCC.n2289 VCC.n2288 1.13717
R7550 VCC.n2285 VCC.n2284 1.13717
R7551 VCC.n2959 VCC.n2958 1.13717
R7552 VCC.n2957 VCC.n2943 1.13717
R7553 VCC.n3014 VCC.n3013 1.13717
R7554 VCC.n2934 VCC.n2917 1.13717
R7555 VCC.n2902 VCC.n2901 1.13717
R7556 VCC.n2898 VCC.n2897 1.13717
R7557 VCC.n3086 VCC.n2896 1.13717
R7558 VCC.n3116 VCC.n3115 1.13717
R7559 VCC.n3140 VCC.n3139 1.13717
R7560 VCC.n3143 VCC.n2857 1.13717
R7561 VCC.n2841 VCC.n2840 1.13717
R7562 VCC.n2837 VCC.n2836 1.13717
R7563 VCC.n2833 VCC.n2832 1.13717
R7564 VCC.n2831 VCC.n2819 1.13717
R7565 VCC.n3254 VCC.n3253 1.13717
R7566 VCC.n2804 VCC.n2800 1.13717
R7567 VCC.n2784 VCC.n2783 1.13717
R7568 VCC.n2773 VCC.n2772 1.13717
R7569 VCC.n3517 VCC.n3516 1.13717
R7570 VCC.n3515 VCC.n3501 1.13717
R7571 VCC.n3572 VCC.n3571 1.13717
R7572 VCC.n3492 VCC.n3475 1.13717
R7573 VCC.n3460 VCC.n3459 1.13717
R7574 VCC.n3456 VCC.n3455 1.13717
R7575 VCC.n3644 VCC.n3454 1.13717
R7576 VCC.n3388 VCC.n3372 1.13717
R7577 VCC.n3820 VCC.n3819 1.13717
R7578 VCC.n3827 VCC.n3348 1.13717
R7579 VCC.n3345 VCC.n3344 1.13717
R7580 VCC.n3327 VCC.n3326 1.13717
R7581 VCC.n3390 VCC.n3389 1.13717
R7582 VCC.n3673 VCC.n3672 1.13717
R7583 VCC.n3697 VCC.n3696 1.13717
R7584 VCC.n3700 VCC.n3414 1.13717
R7585 VCC.n3398 VCC.n3397 1.13717
R7586 VCC.n3394 VCC.n3393 1.13717
R7587 VCC.n4068 VCC.n4067 1.13717
R7588 VCC.n4066 VCC.n4052 1.13717
R7589 VCC.n4123 VCC.n4122 1.13717
R7590 VCC.n4043 VCC.n4026 1.13717
R7591 VCC.n4011 VCC.n4010 1.13717
R7592 VCC.n4007 VCC.n4006 1.13717
R7593 VCC.n4195 VCC.n4005 1.13717
R7594 VCC.n4225 VCC.n4224 1.13717
R7595 VCC.n4249 VCC.n4248 1.13717
R7596 VCC.n4252 VCC.n3966 1.13717
R7597 VCC.n3950 VCC.n3949 1.13717
R7598 VCC.n3946 VCC.n3945 1.13717
R7599 VCC.n3942 VCC.n3941 1.13717
R7600 VCC.n3940 VCC.n3928 1.13717
R7601 VCC.n4363 VCC.n4362 1.13717
R7602 VCC.n3913 VCC.n3909 1.13717
R7603 VCC.n3893 VCC.n3892 1.13717
R7604 VCC.n3882 VCC.n3881 1.13717
R7605 VCC.n4626 VCC.n4625 1.13717
R7606 VCC.n4624 VCC.n4610 1.13717
R7607 VCC.n4681 VCC.n4680 1.13717
R7608 VCC.n4601 VCC.n4584 1.13717
R7609 VCC.n4569 VCC.n4568 1.13717
R7610 VCC.n4565 VCC.n4564 1.13717
R7611 VCC.n4753 VCC.n4563 1.13717
R7612 VCC.n4497 VCC.n4481 1.13717
R7613 VCC.n4929 VCC.n4928 1.13717
R7614 VCC.n4936 VCC.n4457 1.13717
R7615 VCC.n4454 VCC.n4453 1.13717
R7616 VCC.n4436 VCC.n4435 1.13717
R7617 VCC.n4499 VCC.n4498 1.13717
R7618 VCC.n4782 VCC.n4781 1.13717
R7619 VCC.n4806 VCC.n4805 1.13717
R7620 VCC.n4809 VCC.n4523 1.13717
R7621 VCC.n4507 VCC.n4506 1.13717
R7622 VCC.n4503 VCC.n4502 1.13717
R7623 VCC.n5177 VCC.n5176 1.13717
R7624 VCC.n5175 VCC.n5161 1.13717
R7625 VCC.n5232 VCC.n5231 1.13717
R7626 VCC.n5152 VCC.n5135 1.13717
R7627 VCC.n5120 VCC.n5119 1.13717
R7628 VCC.n5116 VCC.n5115 1.13717
R7629 VCC.n5304 VCC.n5114 1.13717
R7630 VCC.n5334 VCC.n5333 1.13717
R7631 VCC.n5358 VCC.n5357 1.13717
R7632 VCC.n5361 VCC.n5075 1.13717
R7633 VCC.n5059 VCC.n5058 1.13717
R7634 VCC.n5055 VCC.n5054 1.13717
R7635 VCC.n5051 VCC.n5050 1.13717
R7636 VCC.n5049 VCC.n5037 1.13717
R7637 VCC.n5472 VCC.n5471 1.13717
R7638 VCC.n5022 VCC.n5018 1.13717
R7639 VCC.n5002 VCC.n5001 1.13717
R7640 VCC.n4991 VCC.n4990 1.13717
R7641 VCC.n5734 VCC.n5733 1.13717
R7642 VCC.n5732 VCC.n5718 1.13717
R7643 VCC.n5789 VCC.n5788 1.13717
R7644 VCC.n5709 VCC.n5692 1.13717
R7645 VCC.n5677 VCC.n5676 1.13717
R7646 VCC.n5673 VCC.n5672 1.13717
R7647 VCC.n5861 VCC.n5671 1.13717
R7648 VCC.n5605 VCC.n5589 1.13717
R7649 VCC.n6037 VCC.n6036 1.13717
R7650 VCC.n6044 VCC.n5565 1.13717
R7651 VCC.n5562 VCC.n5561 1.13717
R7652 VCC.n5544 VCC.n5543 1.13717
R7653 VCC.n5607 VCC.n5606 1.13717
R7654 VCC.n5890 VCC.n5889 1.13717
R7655 VCC.n5914 VCC.n5913 1.13717
R7656 VCC.n5917 VCC.n5631 1.13717
R7657 VCC.n5615 VCC.n5614 1.13717
R7658 VCC.n5611 VCC.n5610 1.13717
R7659 VCC.n6284 VCC.n6283 1.13717
R7660 VCC.n6282 VCC.n6268 1.13717
R7661 VCC.n6339 VCC.n6338 1.13717
R7662 VCC.n6259 VCC.n6242 1.13717
R7663 VCC.n6227 VCC.n6226 1.13717
R7664 VCC.n6223 VCC.n6222 1.13717
R7665 VCC.n6411 VCC.n6221 1.13717
R7666 VCC.n6441 VCC.n6440 1.13717
R7667 VCC.n6465 VCC.n6464 1.13717
R7668 VCC.n6468 VCC.n6182 1.13717
R7669 VCC.n6166 VCC.n6165 1.13717
R7670 VCC.n6162 VCC.n6161 1.13717
R7671 VCC.n6158 VCC.n6157 1.13717
R7672 VCC.n6156 VCC.n6144 1.13717
R7673 VCC.n6579 VCC.n6578 1.13717
R7674 VCC.n6129 VCC.n6125 1.13717
R7675 VCC.n6109 VCC.n6108 1.13717
R7676 VCC.n6098 VCC.n6097 1.13717
R7677 VCC.n6841 VCC.n6840 1.13717
R7678 VCC.n6839 VCC.n6825 1.13717
R7679 VCC.n6896 VCC.n6895 1.13717
R7680 VCC.n6816 VCC.n6799 1.13717
R7681 VCC.n6784 VCC.n6783 1.13717
R7682 VCC.n6780 VCC.n6779 1.13717
R7683 VCC.n6968 VCC.n6778 1.13717
R7684 VCC.n6712 VCC.n6696 1.13717
R7685 VCC.n7144 VCC.n7143 1.13717
R7686 VCC.n7151 VCC.n6672 1.13717
R7687 VCC.n6669 VCC.n6668 1.13717
R7688 VCC.n6651 VCC.n6650 1.13717
R7689 VCC.n6714 VCC.n6713 1.13717
R7690 VCC.n6997 VCC.n6996 1.13717
R7691 VCC.n7021 VCC.n7020 1.13717
R7692 VCC.n7024 VCC.n6738 1.13717
R7693 VCC.n6722 VCC.n6721 1.13717
R7694 VCC.n6718 VCC.n6717 1.13717
R7695 VCC.n7391 VCC.n7390 1.13717
R7696 VCC.n7389 VCC.n7375 1.13717
R7697 VCC.n7446 VCC.n7445 1.13717
R7698 VCC.n7366 VCC.n7349 1.13717
R7699 VCC.n7334 VCC.n7333 1.13717
R7700 VCC.n7330 VCC.n7329 1.13717
R7701 VCC.n7518 VCC.n7328 1.13717
R7702 VCC.n7548 VCC.n7547 1.13717
R7703 VCC.n7572 VCC.n7571 1.13717
R7704 VCC.n7575 VCC.n7289 1.13717
R7705 VCC.n7273 VCC.n7272 1.13717
R7706 VCC.n7269 VCC.n7268 1.13717
R7707 VCC.n7265 VCC.n7264 1.13717
R7708 VCC.n7263 VCC.n7251 1.13717
R7709 VCC.n7686 VCC.n7685 1.13717
R7710 VCC.n7236 VCC.n7232 1.13717
R7711 VCC.n7216 VCC.n7215 1.13717
R7712 VCC.n7205 VCC.n7204 1.13717
R7713 VCC.n7948 VCC.n7947 1.13717
R7714 VCC.n7946 VCC.n7932 1.13717
R7715 VCC.n8003 VCC.n8002 1.13717
R7716 VCC.n7923 VCC.n7906 1.13717
R7717 VCC.n7891 VCC.n7890 1.13717
R7718 VCC.n7887 VCC.n7886 1.13717
R7719 VCC.n8075 VCC.n7885 1.13717
R7720 VCC.n7819 VCC.n7803 1.13717
R7721 VCC.n8251 VCC.n8250 1.13717
R7722 VCC.n8258 VCC.n7779 1.13717
R7723 VCC.n7776 VCC.n7775 1.13717
R7724 VCC.n7758 VCC.n7757 1.13717
R7725 VCC.n7821 VCC.n7820 1.13717
R7726 VCC.n8104 VCC.n8103 1.13717
R7727 VCC.n8128 VCC.n8127 1.13717
R7728 VCC.n8131 VCC.n7845 1.13717
R7729 VCC.n7829 VCC.n7828 1.13717
R7730 VCC.n7825 VCC.n7824 1.13717
R7731 VCC.n8438 VCC.n8435 1.13717
R7732 VCC.n8468 VCC.n8467 1.13717
R7733 VCC.n8492 VCC.n8491 1.13717
R7734 VCC.n8495 VCC.n8396 1.13717
R7735 VCC.n8380 VCC.n8379 1.13717
R7736 VCC.n8376 VCC.n8375 1.13717
R7737 VCC.n8372 VCC.n8371 1.13717
R7738 VCC.n8370 VCC.n8358 1.13717
R7739 VCC.n8606 VCC.n8605 1.13717
R7740 VCC.n8343 VCC.n8339 1.13717
R7741 VCC.n8323 VCC.n8322 1.13717
R7742 VCC.n8312 VCC.n8311 1.13717
R7743 VCC.n376 VCC.n101 1.1255
R7744 VCC.n500 VCC.n37 1.1255
R7745 VCC.n928 VCC.n653 1.1255
R7746 VCC.n1052 VCC.n589 1.1255
R7747 VCC.n1615 VCC.n1147 1.1255
R7748 VCC.n1485 VCC.n1210 1.1255
R7749 VCC.n2037 VCC.n1762 1.1255
R7750 VCC.n2161 VCC.n1698 1.1255
R7751 VCC.n2724 VCC.n2256 1.1255
R7752 VCC.n2594 VCC.n2319 1.1255
R7753 VCC.n3146 VCC.n2871 1.1255
R7754 VCC.n3270 VCC.n2807 1.1255
R7755 VCC.n3833 VCC.n3365 1.1255
R7756 VCC.n3703 VCC.n3428 1.1255
R7757 VCC.n4255 VCC.n3980 1.1255
R7758 VCC.n4379 VCC.n3916 1.1255
R7759 VCC.n4942 VCC.n4474 1.1255
R7760 VCC.n4812 VCC.n4537 1.1255
R7761 VCC.n5364 VCC.n5089 1.1255
R7762 VCC.n5488 VCC.n5025 1.1255
R7763 VCC.n6050 VCC.n5582 1.1255
R7764 VCC.n5920 VCC.n5645 1.1255
R7765 VCC.n6471 VCC.n6196 1.1255
R7766 VCC.n6595 VCC.n6132 1.1255
R7767 VCC.n7157 VCC.n6689 1.1255
R7768 VCC.n7027 VCC.n6752 1.1255
R7769 VCC.n7578 VCC.n7303 1.1255
R7770 VCC.n7702 VCC.n7239 1.1255
R7771 VCC.n8264 VCC.n7796 1.1255
R7772 VCC.n8134 VCC.n7859 1.1255
R7773 VCC.n8498 VCC.n8410 1.1255
R7774 VCC.n8622 VCC.n8346 1.1255
R7775 VCC.n213 VCC.n207 1.00621
R7776 VCC.n201 VCC.n195 1.00621
R7777 VCC.n160 VCC.n159 1.00621
R7778 VCC.n333 VCC.n124 1.00621
R7779 VCC.n326 VCC.n325 1.00621
R7780 VCC.n391 VCC.n95 1.00621
R7781 VCC.n422 VCC.n421 1.00621
R7782 VCC.n545 VCC.n3 1.00621
R7783 VCC.n765 VCC.n759 1.00621
R7784 VCC.n753 VCC.n747 1.00621
R7785 VCC.n712 VCC.n711 1.00621
R7786 VCC.n885 VCC.n676 1.00621
R7787 VCC.n878 VCC.n877 1.00621
R7788 VCC.n943 VCC.n647 1.00621
R7789 VCC.n974 VCC.n973 1.00621
R7790 VCC.n1099 VCC.n557 1.00621
R7791 VCC.n1532 VCC.n1531 1.00621
R7792 VCC.n1656 VCC.n1112 1.00621
R7793 VCC.n1442 VCC.n1233 1.00621
R7794 VCC.n1435 VCC.n1434 1.00621
R7795 VCC.n1500 VCC.n1204 1.00621
R7796 VCC.n1323 VCC.n1317 1.00621
R7797 VCC.n1311 VCC.n1305 1.00621
R7798 VCC.n1270 VCC.n1269 1.00621
R7799 VCC.n1874 VCC.n1868 1.00621
R7800 VCC.n1862 VCC.n1856 1.00621
R7801 VCC.n1821 VCC.n1820 1.00621
R7802 VCC.n1994 VCC.n1785 1.00621
R7803 VCC.n1987 VCC.n1986 1.00621
R7804 VCC.n2052 VCC.n1756 1.00621
R7805 VCC.n2083 VCC.n2082 1.00621
R7806 VCC.n2208 VCC.n1666 1.00621
R7807 VCC.n2641 VCC.n2640 1.00621
R7808 VCC.n2765 VCC.n2221 1.00621
R7809 VCC.n2551 VCC.n2342 1.00621
R7810 VCC.n2544 VCC.n2543 1.00621
R7811 VCC.n2609 VCC.n2313 1.00621
R7812 VCC.n2432 VCC.n2426 1.00621
R7813 VCC.n2420 VCC.n2414 1.00621
R7814 VCC.n2379 VCC.n2378 1.00621
R7815 VCC.n2983 VCC.n2977 1.00621
R7816 VCC.n2971 VCC.n2965 1.00621
R7817 VCC.n2930 VCC.n2929 1.00621
R7818 VCC.n3103 VCC.n2894 1.00621
R7819 VCC.n3096 VCC.n3095 1.00621
R7820 VCC.n3161 VCC.n2865 1.00621
R7821 VCC.n3192 VCC.n3191 1.00621
R7822 VCC.n3317 VCC.n2775 1.00621
R7823 VCC.n3750 VCC.n3749 1.00621
R7824 VCC.n3874 VCC.n3330 1.00621
R7825 VCC.n3660 VCC.n3451 1.00621
R7826 VCC.n3653 VCC.n3652 1.00621
R7827 VCC.n3718 VCC.n3422 1.00621
R7828 VCC.n3541 VCC.n3535 1.00621
R7829 VCC.n3529 VCC.n3523 1.00621
R7830 VCC.n3488 VCC.n3487 1.00621
R7831 VCC.n4092 VCC.n4086 1.00621
R7832 VCC.n4080 VCC.n4074 1.00621
R7833 VCC.n4039 VCC.n4038 1.00621
R7834 VCC.n4212 VCC.n4003 1.00621
R7835 VCC.n4205 VCC.n4204 1.00621
R7836 VCC.n4270 VCC.n3974 1.00621
R7837 VCC.n4301 VCC.n4300 1.00621
R7838 VCC.n4426 VCC.n3884 1.00621
R7839 VCC.n4859 VCC.n4858 1.00621
R7840 VCC.n4983 VCC.n4439 1.00621
R7841 VCC.n4769 VCC.n4560 1.00621
R7842 VCC.n4762 VCC.n4761 1.00621
R7843 VCC.n4827 VCC.n4531 1.00621
R7844 VCC.n4650 VCC.n4644 1.00621
R7845 VCC.n4638 VCC.n4632 1.00621
R7846 VCC.n4597 VCC.n4596 1.00621
R7847 VCC.n5201 VCC.n5195 1.00621
R7848 VCC.n5189 VCC.n5183 1.00621
R7849 VCC.n5148 VCC.n5147 1.00621
R7850 VCC.n5321 VCC.n5112 1.00621
R7851 VCC.n5314 VCC.n5313 1.00621
R7852 VCC.n5379 VCC.n5083 1.00621
R7853 VCC.n5410 VCC.n5409 1.00621
R7854 VCC.n5535 VCC.n4993 1.00621
R7855 VCC.n5967 VCC.n5966 1.00621
R7856 VCC.n6091 VCC.n5547 1.00621
R7857 VCC.n5877 VCC.n5668 1.00621
R7858 VCC.n5870 VCC.n5869 1.00621
R7859 VCC.n5935 VCC.n5639 1.00621
R7860 VCC.n5758 VCC.n5752 1.00621
R7861 VCC.n5746 VCC.n5740 1.00621
R7862 VCC.n5705 VCC.n5704 1.00621
R7863 VCC.n6308 VCC.n6302 1.00621
R7864 VCC.n6296 VCC.n6290 1.00621
R7865 VCC.n6255 VCC.n6254 1.00621
R7866 VCC.n6428 VCC.n6219 1.00621
R7867 VCC.n6421 VCC.n6420 1.00621
R7868 VCC.n6486 VCC.n6190 1.00621
R7869 VCC.n6517 VCC.n6516 1.00621
R7870 VCC.n6642 VCC.n6100 1.00621
R7871 VCC.n7074 VCC.n7073 1.00621
R7872 VCC.n7198 VCC.n6654 1.00621
R7873 VCC.n6984 VCC.n6775 1.00621
R7874 VCC.n6977 VCC.n6976 1.00621
R7875 VCC.n7042 VCC.n6746 1.00621
R7876 VCC.n6865 VCC.n6859 1.00621
R7877 VCC.n6853 VCC.n6847 1.00621
R7878 VCC.n6812 VCC.n6811 1.00621
R7879 VCC.n7415 VCC.n7409 1.00621
R7880 VCC.n7403 VCC.n7397 1.00621
R7881 VCC.n7362 VCC.n7361 1.00621
R7882 VCC.n7535 VCC.n7326 1.00621
R7883 VCC.n7528 VCC.n7527 1.00621
R7884 VCC.n7593 VCC.n7297 1.00621
R7885 VCC.n7624 VCC.n7623 1.00621
R7886 VCC.n7749 VCC.n7207 1.00621
R7887 VCC.n8181 VCC.n8180 1.00621
R7888 VCC.n8305 VCC.n7761 1.00621
R7889 VCC.n8091 VCC.n7882 1.00621
R7890 VCC.n8084 VCC.n8083 1.00621
R7891 VCC.n8149 VCC.n7853 1.00621
R7892 VCC.n7972 VCC.n7966 1.00621
R7893 VCC.n7960 VCC.n7954 1.00621
R7894 VCC.n7919 VCC.n7918 1.00621
R7895 VCC.n8455 VCC.n8433 1.00621
R7896 VCC.n8448 VCC.n8447 1.00621
R7897 VCC.n8513 VCC.n8404 1.00621
R7898 VCC.n8544 VCC.n8543 1.00621
R7899 VCC.n8669 VCC.n8314 1.00621
R7900 VCC.n230 VCC.n180 0.9505
R7901 VCC.n269 VCC.n143 0.9505
R7902 VCC.n359 VCC.n107 0.9505
R7903 VCC.n397 VCC.n92 0.9505
R7904 VCC.n782 VCC.n732 0.9505
R7905 VCC.n821 VCC.n695 0.9505
R7906 VCC.n911 VCC.n659 0.9505
R7907 VCC.n949 VCC.n644 0.9505
R7908 VCC.n1468 VCC.n1216 0.9505
R7909 VCC.n1506 VCC.n1201 0.9505
R7910 VCC.n1340 VCC.n1290 0.9505
R7911 VCC.n1379 VCC.n1253 0.9505
R7912 VCC.n1891 VCC.n1841 0.9505
R7913 VCC.n1930 VCC.n1804 0.9505
R7914 VCC.n2020 VCC.n1768 0.9505
R7915 VCC.n2058 VCC.n1753 0.9505
R7916 VCC.n2577 VCC.n2325 0.9505
R7917 VCC.n2615 VCC.n2310 0.9505
R7918 VCC.n2449 VCC.n2399 0.9505
R7919 VCC.n2488 VCC.n2362 0.9505
R7920 VCC.n3000 VCC.n2950 0.9505
R7921 VCC.n3039 VCC.n2913 0.9505
R7922 VCC.n3129 VCC.n2877 0.9505
R7923 VCC.n3167 VCC.n2862 0.9505
R7924 VCC.n3686 VCC.n3434 0.9505
R7925 VCC.n3724 VCC.n3419 0.9505
R7926 VCC.n3558 VCC.n3508 0.9505
R7927 VCC.n3597 VCC.n3471 0.9505
R7928 VCC.n4109 VCC.n4059 0.9505
R7929 VCC.n4148 VCC.n4022 0.9505
R7930 VCC.n4238 VCC.n3986 0.9505
R7931 VCC.n4276 VCC.n3971 0.9505
R7932 VCC.n4795 VCC.n4543 0.9505
R7933 VCC.n4833 VCC.n4528 0.9505
R7934 VCC.n4667 VCC.n4617 0.9505
R7935 VCC.n4706 VCC.n4580 0.9505
R7936 VCC.n5218 VCC.n5168 0.9505
R7937 VCC.n5257 VCC.n5131 0.9505
R7938 VCC.n5347 VCC.n5095 0.9505
R7939 VCC.n5385 VCC.n5080 0.9505
R7940 VCC.n5903 VCC.n5651 0.9505
R7941 VCC.n5941 VCC.n5636 0.9505
R7942 VCC.n5775 VCC.n5725 0.9505
R7943 VCC.n5814 VCC.n5688 0.9505
R7944 VCC.n6325 VCC.n6275 0.9505
R7945 VCC.n6364 VCC.n6238 0.9505
R7946 VCC.n6454 VCC.n6202 0.9505
R7947 VCC.n6492 VCC.n6187 0.9505
R7948 VCC.n7010 VCC.n6758 0.9505
R7949 VCC.n7048 VCC.n6743 0.9505
R7950 VCC.n6882 VCC.n6832 0.9505
R7951 VCC.n6921 VCC.n6795 0.9505
R7952 VCC.n7432 VCC.n7382 0.9505
R7953 VCC.n7471 VCC.n7345 0.9505
R7954 VCC.n7561 VCC.n7309 0.9505
R7955 VCC.n7599 VCC.n7294 0.9505
R7956 VCC.n8117 VCC.n7865 0.9505
R7957 VCC.n8155 VCC.n7850 0.9505
R7958 VCC.n7989 VCC.n7939 0.9505
R7959 VCC.n8028 VCC.n7902 0.9505
R7960 VCC.n8481 VCC.n8416 0.9505
R7961 VCC.n8519 VCC.n8401 0.9505
R7962 VCC.n248 VCC.n247 0.914786
R7963 VCC.n263 VCC.n156 0.914786
R7964 VCC.n297 VCC.n139 0.914786
R7965 VCC.n296 VCC.n295 0.914786
R7966 VCC.n366 VCC.n365 0.914786
R7967 VCC.n384 VCC.n97 0.914786
R7968 VCC.n432 VCC.n78 0.914786
R7969 VCC.n431 VCC.n430 0.914786
R7970 VCC.n800 VCC.n799 0.914786
R7971 VCC.n815 VCC.n708 0.914786
R7972 VCC.n849 VCC.n691 0.914786
R7973 VCC.n848 VCC.n847 0.914786
R7974 VCC.n918 VCC.n917 0.914786
R7975 VCC.n936 VCC.n649 0.914786
R7976 VCC.n984 VCC.n630 0.914786
R7977 VCC.n983 VCC.n982 0.914786
R7978 VCC.n1475 VCC.n1474 0.914786
R7979 VCC.n1493 VCC.n1206 0.914786
R7980 VCC.n1542 VCC.n1187 0.914786
R7981 VCC.n1541 VCC.n1540 0.914786
R7982 VCC.n1358 VCC.n1357 0.914786
R7983 VCC.n1373 VCC.n1266 0.914786
R7984 VCC.n1407 VCC.n1249 0.914786
R7985 VCC.n1406 VCC.n1405 0.914786
R7986 VCC.n1909 VCC.n1908 0.914786
R7987 VCC.n1924 VCC.n1817 0.914786
R7988 VCC.n1958 VCC.n1800 0.914786
R7989 VCC.n1957 VCC.n1956 0.914786
R7990 VCC.n2027 VCC.n2026 0.914786
R7991 VCC.n2045 VCC.n1758 0.914786
R7992 VCC.n2093 VCC.n1739 0.914786
R7993 VCC.n2092 VCC.n2091 0.914786
R7994 VCC.n2584 VCC.n2583 0.914786
R7995 VCC.n2602 VCC.n2315 0.914786
R7996 VCC.n2651 VCC.n2296 0.914786
R7997 VCC.n2650 VCC.n2649 0.914786
R7998 VCC.n2467 VCC.n2466 0.914786
R7999 VCC.n2482 VCC.n2375 0.914786
R8000 VCC.n2516 VCC.n2358 0.914786
R8001 VCC.n2515 VCC.n2514 0.914786
R8002 VCC.n3018 VCC.n3017 0.914786
R8003 VCC.n3033 VCC.n2926 0.914786
R8004 VCC.n3067 VCC.n2909 0.914786
R8005 VCC.n3066 VCC.n3065 0.914786
R8006 VCC.n3136 VCC.n3135 0.914786
R8007 VCC.n3154 VCC.n2867 0.914786
R8008 VCC.n3202 VCC.n2848 0.914786
R8009 VCC.n3201 VCC.n3200 0.914786
R8010 VCC.n3693 VCC.n3692 0.914786
R8011 VCC.n3711 VCC.n3424 0.914786
R8012 VCC.n3760 VCC.n3405 0.914786
R8013 VCC.n3759 VCC.n3758 0.914786
R8014 VCC.n3576 VCC.n3575 0.914786
R8015 VCC.n3591 VCC.n3484 0.914786
R8016 VCC.n3625 VCC.n3467 0.914786
R8017 VCC.n3624 VCC.n3623 0.914786
R8018 VCC.n4127 VCC.n4126 0.914786
R8019 VCC.n4142 VCC.n4035 0.914786
R8020 VCC.n4176 VCC.n4018 0.914786
R8021 VCC.n4175 VCC.n4174 0.914786
R8022 VCC.n4245 VCC.n4244 0.914786
R8023 VCC.n4263 VCC.n3976 0.914786
R8024 VCC.n4311 VCC.n3957 0.914786
R8025 VCC.n4310 VCC.n4309 0.914786
R8026 VCC.n4802 VCC.n4801 0.914786
R8027 VCC.n4820 VCC.n4533 0.914786
R8028 VCC.n4869 VCC.n4514 0.914786
R8029 VCC.n4868 VCC.n4867 0.914786
R8030 VCC.n4685 VCC.n4684 0.914786
R8031 VCC.n4700 VCC.n4593 0.914786
R8032 VCC.n4734 VCC.n4576 0.914786
R8033 VCC.n4733 VCC.n4732 0.914786
R8034 VCC.n5236 VCC.n5235 0.914786
R8035 VCC.n5251 VCC.n5144 0.914786
R8036 VCC.n5285 VCC.n5127 0.914786
R8037 VCC.n5284 VCC.n5283 0.914786
R8038 VCC.n5354 VCC.n5353 0.914786
R8039 VCC.n5372 VCC.n5085 0.914786
R8040 VCC.n5420 VCC.n5066 0.914786
R8041 VCC.n5419 VCC.n5418 0.914786
R8042 VCC.n5910 VCC.n5909 0.914786
R8043 VCC.n5928 VCC.n5641 0.914786
R8044 VCC.n5977 VCC.n5622 0.914786
R8045 VCC.n5976 VCC.n5975 0.914786
R8046 VCC.n5793 VCC.n5792 0.914786
R8047 VCC.n5808 VCC.n5701 0.914786
R8048 VCC.n5842 VCC.n5684 0.914786
R8049 VCC.n5841 VCC.n5840 0.914786
R8050 VCC.n6343 VCC.n6342 0.914786
R8051 VCC.n6358 VCC.n6251 0.914786
R8052 VCC.n6392 VCC.n6234 0.914786
R8053 VCC.n6391 VCC.n6390 0.914786
R8054 VCC.n6461 VCC.n6460 0.914786
R8055 VCC.n6479 VCC.n6192 0.914786
R8056 VCC.n6527 VCC.n6173 0.914786
R8057 VCC.n6526 VCC.n6525 0.914786
R8058 VCC.n7017 VCC.n7016 0.914786
R8059 VCC.n7035 VCC.n6748 0.914786
R8060 VCC.n7084 VCC.n6729 0.914786
R8061 VCC.n7083 VCC.n7082 0.914786
R8062 VCC.n6900 VCC.n6899 0.914786
R8063 VCC.n6915 VCC.n6808 0.914786
R8064 VCC.n6949 VCC.n6791 0.914786
R8065 VCC.n6948 VCC.n6947 0.914786
R8066 VCC.n7450 VCC.n7449 0.914786
R8067 VCC.n7465 VCC.n7358 0.914786
R8068 VCC.n7499 VCC.n7341 0.914786
R8069 VCC.n7498 VCC.n7497 0.914786
R8070 VCC.n7568 VCC.n7567 0.914786
R8071 VCC.n7586 VCC.n7299 0.914786
R8072 VCC.n7634 VCC.n7280 0.914786
R8073 VCC.n7633 VCC.n7632 0.914786
R8074 VCC.n8124 VCC.n8123 0.914786
R8075 VCC.n8142 VCC.n7855 0.914786
R8076 VCC.n8191 VCC.n7836 0.914786
R8077 VCC.n8190 VCC.n8189 0.914786
R8078 VCC.n8007 VCC.n8006 0.914786
R8079 VCC.n8022 VCC.n7915 0.914786
R8080 VCC.n8056 VCC.n7898 0.914786
R8081 VCC.n8055 VCC.n8054 0.914786
R8082 VCC.n8488 VCC.n8487 0.914786
R8083 VCC.n8506 VCC.n8406 0.914786
R8084 VCC.n8554 VCC.n8387 0.914786
R8085 VCC.n8553 VCC.n8552 0.914786
R8086 VCC.n223 VCC.n184 0.823357
R8087 VCC.n232 VCC.n177 0.823357
R8088 VCC.n249 VCC.n155 0.823357
R8089 VCC.n285 VCC.n144 0.823357
R8090 VCC.n341 VCC.n340 0.823357
R8091 VCC.n357 VCC.n110 0.823357
R8092 VCC.n387 VCC.n386 0.823357
R8093 VCC.n412 VCC.n84 0.823357
R8094 VCC.n775 VCC.n736 0.823357
R8095 VCC.n784 VCC.n729 0.823357
R8096 VCC.n801 VCC.n707 0.823357
R8097 VCC.n837 VCC.n696 0.823357
R8098 VCC.n893 VCC.n892 0.823357
R8099 VCC.n909 VCC.n662 0.823357
R8100 VCC.n939 VCC.n938 0.823357
R8101 VCC.n964 VCC.n636 0.823357
R8102 VCC.n1450 VCC.n1449 0.823357
R8103 VCC.n1466 VCC.n1219 0.823357
R8104 VCC.n1496 VCC.n1495 0.823357
R8105 VCC.n1521 VCC.n1193 0.823357
R8106 VCC.n1333 VCC.n1294 0.823357
R8107 VCC.n1342 VCC.n1287 0.823357
R8108 VCC.n1359 VCC.n1265 0.823357
R8109 VCC.n1395 VCC.n1254 0.823357
R8110 VCC.n1884 VCC.n1845 0.823357
R8111 VCC.n1893 VCC.n1838 0.823357
R8112 VCC.n1910 VCC.n1816 0.823357
R8113 VCC.n1946 VCC.n1805 0.823357
R8114 VCC.n2002 VCC.n2001 0.823357
R8115 VCC.n2018 VCC.n1771 0.823357
R8116 VCC.n2048 VCC.n2047 0.823357
R8117 VCC.n2073 VCC.n1745 0.823357
R8118 VCC.n2559 VCC.n2558 0.823357
R8119 VCC.n2575 VCC.n2328 0.823357
R8120 VCC.n2605 VCC.n2604 0.823357
R8121 VCC.n2630 VCC.n2302 0.823357
R8122 VCC.n2442 VCC.n2403 0.823357
R8123 VCC.n2451 VCC.n2396 0.823357
R8124 VCC.n2468 VCC.n2374 0.823357
R8125 VCC.n2504 VCC.n2363 0.823357
R8126 VCC.n2993 VCC.n2954 0.823357
R8127 VCC.n3002 VCC.n2947 0.823357
R8128 VCC.n3019 VCC.n2925 0.823357
R8129 VCC.n3055 VCC.n2914 0.823357
R8130 VCC.n3111 VCC.n3110 0.823357
R8131 VCC.n3127 VCC.n2880 0.823357
R8132 VCC.n3157 VCC.n3156 0.823357
R8133 VCC.n3182 VCC.n2854 0.823357
R8134 VCC.n3668 VCC.n3667 0.823357
R8135 VCC.n3684 VCC.n3437 0.823357
R8136 VCC.n3714 VCC.n3713 0.823357
R8137 VCC.n3739 VCC.n3411 0.823357
R8138 VCC.n3551 VCC.n3512 0.823357
R8139 VCC.n3560 VCC.n3505 0.823357
R8140 VCC.n3577 VCC.n3483 0.823357
R8141 VCC.n3613 VCC.n3472 0.823357
R8142 VCC.n4102 VCC.n4063 0.823357
R8143 VCC.n4111 VCC.n4056 0.823357
R8144 VCC.n4128 VCC.n4034 0.823357
R8145 VCC.n4164 VCC.n4023 0.823357
R8146 VCC.n4220 VCC.n4219 0.823357
R8147 VCC.n4236 VCC.n3989 0.823357
R8148 VCC.n4266 VCC.n4265 0.823357
R8149 VCC.n4291 VCC.n3963 0.823357
R8150 VCC.n4777 VCC.n4776 0.823357
R8151 VCC.n4793 VCC.n4546 0.823357
R8152 VCC.n4823 VCC.n4822 0.823357
R8153 VCC.n4848 VCC.n4520 0.823357
R8154 VCC.n4660 VCC.n4621 0.823357
R8155 VCC.n4669 VCC.n4614 0.823357
R8156 VCC.n4686 VCC.n4592 0.823357
R8157 VCC.n4722 VCC.n4581 0.823357
R8158 VCC.n5211 VCC.n5172 0.823357
R8159 VCC.n5220 VCC.n5165 0.823357
R8160 VCC.n5237 VCC.n5143 0.823357
R8161 VCC.n5273 VCC.n5132 0.823357
R8162 VCC.n5329 VCC.n5328 0.823357
R8163 VCC.n5345 VCC.n5098 0.823357
R8164 VCC.n5375 VCC.n5374 0.823357
R8165 VCC.n5400 VCC.n5072 0.823357
R8166 VCC.n5885 VCC.n5884 0.823357
R8167 VCC.n5901 VCC.n5654 0.823357
R8168 VCC.n5931 VCC.n5930 0.823357
R8169 VCC.n5956 VCC.n5628 0.823357
R8170 VCC.n5768 VCC.n5729 0.823357
R8171 VCC.n5777 VCC.n5722 0.823357
R8172 VCC.n5794 VCC.n5700 0.823357
R8173 VCC.n5830 VCC.n5689 0.823357
R8174 VCC.n6318 VCC.n6279 0.823357
R8175 VCC.n6327 VCC.n6272 0.823357
R8176 VCC.n6344 VCC.n6250 0.823357
R8177 VCC.n6380 VCC.n6239 0.823357
R8178 VCC.n6436 VCC.n6435 0.823357
R8179 VCC.n6452 VCC.n6205 0.823357
R8180 VCC.n6482 VCC.n6481 0.823357
R8181 VCC.n6507 VCC.n6179 0.823357
R8182 VCC.n6992 VCC.n6991 0.823357
R8183 VCC.n7008 VCC.n6761 0.823357
R8184 VCC.n7038 VCC.n7037 0.823357
R8185 VCC.n7063 VCC.n6735 0.823357
R8186 VCC.n6875 VCC.n6836 0.823357
R8187 VCC.n6884 VCC.n6829 0.823357
R8188 VCC.n6901 VCC.n6807 0.823357
R8189 VCC.n6937 VCC.n6796 0.823357
R8190 VCC.n7425 VCC.n7386 0.823357
R8191 VCC.n7434 VCC.n7379 0.823357
R8192 VCC.n7451 VCC.n7357 0.823357
R8193 VCC.n7487 VCC.n7346 0.823357
R8194 VCC.n7543 VCC.n7542 0.823357
R8195 VCC.n7559 VCC.n7312 0.823357
R8196 VCC.n7589 VCC.n7588 0.823357
R8197 VCC.n7614 VCC.n7286 0.823357
R8198 VCC.n8099 VCC.n8098 0.823357
R8199 VCC.n8115 VCC.n7868 0.823357
R8200 VCC.n8145 VCC.n8144 0.823357
R8201 VCC.n8170 VCC.n7842 0.823357
R8202 VCC.n7982 VCC.n7943 0.823357
R8203 VCC.n7991 VCC.n7936 0.823357
R8204 VCC.n8008 VCC.n7914 0.823357
R8205 VCC.n8044 VCC.n7903 0.823357
R8206 VCC.n8463 VCC.n8462 0.823357
R8207 VCC.n8479 VCC.n8419 0.823357
R8208 VCC.n8509 VCC.n8508 0.823357
R8209 VCC.n8534 VCC.n8393 0.823357
R8210 VCC.n184 VCC.n177 0.731929
R8211 VCC.n272 VCC.n144 0.731929
R8212 VCC.n287 VCC.n285 0.731929
R8213 VCC.n340 VCC.n110 0.731929
R8214 VCC.n399 VCC.n84 0.731929
R8215 VCC.n413 VCC.n412 0.731929
R8216 VCC.n736 VCC.n729 0.731929
R8217 VCC.n824 VCC.n696 0.731929
R8218 VCC.n839 VCC.n837 0.731929
R8219 VCC.n892 VCC.n662 0.731929
R8220 VCC.n951 VCC.n636 0.731929
R8221 VCC.n965 VCC.n964 0.731929
R8222 VCC.n1449 VCC.n1219 0.731929
R8223 VCC.n1508 VCC.n1193 0.731929
R8224 VCC.n1522 VCC.n1521 0.731929
R8225 VCC.n1294 VCC.n1287 0.731929
R8226 VCC.n1382 VCC.n1254 0.731929
R8227 VCC.n1397 VCC.n1395 0.731929
R8228 VCC.n1845 VCC.n1838 0.731929
R8229 VCC.n1933 VCC.n1805 0.731929
R8230 VCC.n1948 VCC.n1946 0.731929
R8231 VCC.n2001 VCC.n1771 0.731929
R8232 VCC.n2060 VCC.n1745 0.731929
R8233 VCC.n2074 VCC.n2073 0.731929
R8234 VCC.n2558 VCC.n2328 0.731929
R8235 VCC.n2617 VCC.n2302 0.731929
R8236 VCC.n2631 VCC.n2630 0.731929
R8237 VCC.n2403 VCC.n2396 0.731929
R8238 VCC.n2491 VCC.n2363 0.731929
R8239 VCC.n2506 VCC.n2504 0.731929
R8240 VCC.n2954 VCC.n2947 0.731929
R8241 VCC.n3042 VCC.n2914 0.731929
R8242 VCC.n3057 VCC.n3055 0.731929
R8243 VCC.n3110 VCC.n2880 0.731929
R8244 VCC.n3169 VCC.n2854 0.731929
R8245 VCC.n3183 VCC.n3182 0.731929
R8246 VCC.n3667 VCC.n3437 0.731929
R8247 VCC.n3726 VCC.n3411 0.731929
R8248 VCC.n3740 VCC.n3739 0.731929
R8249 VCC.n3512 VCC.n3505 0.731929
R8250 VCC.n3600 VCC.n3472 0.731929
R8251 VCC.n3615 VCC.n3613 0.731929
R8252 VCC.n4063 VCC.n4056 0.731929
R8253 VCC.n4151 VCC.n4023 0.731929
R8254 VCC.n4166 VCC.n4164 0.731929
R8255 VCC.n4219 VCC.n3989 0.731929
R8256 VCC.n4278 VCC.n3963 0.731929
R8257 VCC.n4292 VCC.n4291 0.731929
R8258 VCC.n4776 VCC.n4546 0.731929
R8259 VCC.n4835 VCC.n4520 0.731929
R8260 VCC.n4849 VCC.n4848 0.731929
R8261 VCC.n4621 VCC.n4614 0.731929
R8262 VCC.n4709 VCC.n4581 0.731929
R8263 VCC.n4724 VCC.n4722 0.731929
R8264 VCC.n5172 VCC.n5165 0.731929
R8265 VCC.n5260 VCC.n5132 0.731929
R8266 VCC.n5275 VCC.n5273 0.731929
R8267 VCC.n5328 VCC.n5098 0.731929
R8268 VCC.n5387 VCC.n5072 0.731929
R8269 VCC.n5401 VCC.n5400 0.731929
R8270 VCC.n5884 VCC.n5654 0.731929
R8271 VCC.n5943 VCC.n5628 0.731929
R8272 VCC.n5957 VCC.n5956 0.731929
R8273 VCC.n5729 VCC.n5722 0.731929
R8274 VCC.n5817 VCC.n5689 0.731929
R8275 VCC.n5832 VCC.n5830 0.731929
R8276 VCC.n6279 VCC.n6272 0.731929
R8277 VCC.n6367 VCC.n6239 0.731929
R8278 VCC.n6382 VCC.n6380 0.731929
R8279 VCC.n6435 VCC.n6205 0.731929
R8280 VCC.n6494 VCC.n6179 0.731929
R8281 VCC.n6508 VCC.n6507 0.731929
R8282 VCC.n6991 VCC.n6761 0.731929
R8283 VCC.n7050 VCC.n6735 0.731929
R8284 VCC.n7064 VCC.n7063 0.731929
R8285 VCC.n6836 VCC.n6829 0.731929
R8286 VCC.n6924 VCC.n6796 0.731929
R8287 VCC.n6939 VCC.n6937 0.731929
R8288 VCC.n7386 VCC.n7379 0.731929
R8289 VCC.n7474 VCC.n7346 0.731929
R8290 VCC.n7489 VCC.n7487 0.731929
R8291 VCC.n7542 VCC.n7312 0.731929
R8292 VCC.n7601 VCC.n7286 0.731929
R8293 VCC.n7615 VCC.n7614 0.731929
R8294 VCC.n8098 VCC.n7868 0.731929
R8295 VCC.n8157 VCC.n7842 0.731929
R8296 VCC.n8171 VCC.n8170 0.731929
R8297 VCC.n7943 VCC.n7936 0.731929
R8298 VCC.n8031 VCC.n7903 0.731929
R8299 VCC.n8046 VCC.n8044 0.731929
R8300 VCC.n8462 VCC.n8419 0.731929
R8301 VCC.n8521 VCC.n8393 0.731929
R8302 VCC.n8535 VCC.n8534 0.731929
R8303 VCC.n247 VCC.n169 0.6405
R8304 VCC.n297 VCC.n296 0.6405
R8305 VCC.n366 VCC.n364 0.6405
R8306 VCC.n432 VCC.n431 0.6405
R8307 VCC.n799 VCC.n721 0.6405
R8308 VCC.n849 VCC.n848 0.6405
R8309 VCC.n918 VCC.n916 0.6405
R8310 VCC.n984 VCC.n983 0.6405
R8311 VCC.n1475 VCC.n1473 0.6405
R8312 VCC.n1542 VCC.n1541 0.6405
R8313 VCC.n1357 VCC.n1279 0.6405
R8314 VCC.n1407 VCC.n1406 0.6405
R8315 VCC.n1908 VCC.n1830 0.6405
R8316 VCC.n1958 VCC.n1957 0.6405
R8317 VCC.n2027 VCC.n2025 0.6405
R8318 VCC.n2093 VCC.n2092 0.6405
R8319 VCC.n2584 VCC.n2582 0.6405
R8320 VCC.n2651 VCC.n2650 0.6405
R8321 VCC.n2466 VCC.n2388 0.6405
R8322 VCC.n2516 VCC.n2515 0.6405
R8323 VCC.n3017 VCC.n2939 0.6405
R8324 VCC.n3067 VCC.n3066 0.6405
R8325 VCC.n3136 VCC.n3134 0.6405
R8326 VCC.n3202 VCC.n3201 0.6405
R8327 VCC.n3693 VCC.n3691 0.6405
R8328 VCC.n3760 VCC.n3759 0.6405
R8329 VCC.n3575 VCC.n3497 0.6405
R8330 VCC.n3625 VCC.n3624 0.6405
R8331 VCC.n4126 VCC.n4048 0.6405
R8332 VCC.n4176 VCC.n4175 0.6405
R8333 VCC.n4245 VCC.n4243 0.6405
R8334 VCC.n4311 VCC.n4310 0.6405
R8335 VCC.n4802 VCC.n4800 0.6405
R8336 VCC.n4869 VCC.n4868 0.6405
R8337 VCC.n4684 VCC.n4606 0.6405
R8338 VCC.n4734 VCC.n4733 0.6405
R8339 VCC.n5235 VCC.n5157 0.6405
R8340 VCC.n5285 VCC.n5284 0.6405
R8341 VCC.n5354 VCC.n5352 0.6405
R8342 VCC.n5420 VCC.n5419 0.6405
R8343 VCC.n5910 VCC.n5908 0.6405
R8344 VCC.n5977 VCC.n5976 0.6405
R8345 VCC.n5792 VCC.n5714 0.6405
R8346 VCC.n5842 VCC.n5841 0.6405
R8347 VCC.n6342 VCC.n6264 0.6405
R8348 VCC.n6392 VCC.n6391 0.6405
R8349 VCC.n6461 VCC.n6459 0.6405
R8350 VCC.n6527 VCC.n6526 0.6405
R8351 VCC.n7017 VCC.n7015 0.6405
R8352 VCC.n7084 VCC.n7083 0.6405
R8353 VCC.n6899 VCC.n6821 0.6405
R8354 VCC.n6949 VCC.n6948 0.6405
R8355 VCC.n7449 VCC.n7371 0.6405
R8356 VCC.n7499 VCC.n7498 0.6405
R8357 VCC.n7568 VCC.n7566 0.6405
R8358 VCC.n7634 VCC.n7633 0.6405
R8359 VCC.n8124 VCC.n8122 0.6405
R8360 VCC.n8191 VCC.n8190 0.6405
R8361 VCC.n8006 VCC.n7928 0.6405
R8362 VCC.n8056 VCC.n8055 0.6405
R8363 VCC.n8488 VCC.n8486 0.6405
R8364 VCC.n8554 VCC.n8553 0.6405
R8365 VCC.n4989 VCC 0.621824
R8366 VCC.n207 VCC.n195 0.549071
R8367 VCC.n159 VCC.n151 0.549071
R8368 VCC.n325 VCC.n124 0.549071
R8369 VCC.n392 VCC.n391 0.549071
R8370 VCC.n759 VCC.n747 0.549071
R8371 VCC.n711 VCC.n703 0.549071
R8372 VCC.n877 VCC.n676 0.549071
R8373 VCC.n944 VCC.n943 0.549071
R8374 VCC.n1434 VCC.n1233 0.549071
R8375 VCC.n1501 VCC.n1500 0.549071
R8376 VCC.n1317 VCC.n1305 0.549071
R8377 VCC.n1269 VCC.n1261 0.549071
R8378 VCC.n1868 VCC.n1856 0.549071
R8379 VCC.n1820 VCC.n1812 0.549071
R8380 VCC.n1986 VCC.n1785 0.549071
R8381 VCC.n2053 VCC.n2052 0.549071
R8382 VCC.n2543 VCC.n2342 0.549071
R8383 VCC.n2610 VCC.n2609 0.549071
R8384 VCC.n2426 VCC.n2414 0.549071
R8385 VCC.n2378 VCC.n2370 0.549071
R8386 VCC.n2977 VCC.n2965 0.549071
R8387 VCC.n2929 VCC.n2921 0.549071
R8388 VCC.n3095 VCC.n2894 0.549071
R8389 VCC.n3162 VCC.n3161 0.549071
R8390 VCC.n3652 VCC.n3451 0.549071
R8391 VCC.n3719 VCC.n3718 0.549071
R8392 VCC.n3535 VCC.n3523 0.549071
R8393 VCC.n3487 VCC.n3479 0.549071
R8394 VCC.n4086 VCC.n4074 0.549071
R8395 VCC.n4038 VCC.n4030 0.549071
R8396 VCC.n4204 VCC.n4003 0.549071
R8397 VCC.n4271 VCC.n4270 0.549071
R8398 VCC.n4761 VCC.n4560 0.549071
R8399 VCC.n4828 VCC.n4827 0.549071
R8400 VCC.n4644 VCC.n4632 0.549071
R8401 VCC.n4596 VCC.n4588 0.549071
R8402 VCC.n5195 VCC.n5183 0.549071
R8403 VCC.n5147 VCC.n5139 0.549071
R8404 VCC.n5313 VCC.n5112 0.549071
R8405 VCC.n5380 VCC.n5379 0.549071
R8406 VCC.n5869 VCC.n5668 0.549071
R8407 VCC.n5936 VCC.n5935 0.549071
R8408 VCC.n5752 VCC.n5740 0.549071
R8409 VCC.n5704 VCC.n5696 0.549071
R8410 VCC.n6302 VCC.n6290 0.549071
R8411 VCC.n6254 VCC.n6246 0.549071
R8412 VCC.n6420 VCC.n6219 0.549071
R8413 VCC.n6487 VCC.n6486 0.549071
R8414 VCC.n6976 VCC.n6775 0.549071
R8415 VCC.n7043 VCC.n7042 0.549071
R8416 VCC.n6859 VCC.n6847 0.549071
R8417 VCC.n6811 VCC.n6803 0.549071
R8418 VCC.n7409 VCC.n7397 0.549071
R8419 VCC.n7361 VCC.n7353 0.549071
R8420 VCC.n7527 VCC.n7326 0.549071
R8421 VCC.n7594 VCC.n7593 0.549071
R8422 VCC.n8083 VCC.n7882 0.549071
R8423 VCC.n8150 VCC.n8149 0.549071
R8424 VCC.n7966 VCC.n7954 0.549071
R8425 VCC.n7918 VCC.n7910 0.549071
R8426 VCC.n8447 VCC.n8433 0.549071
R8427 VCC.n8514 VCC.n8513 0.549071
R8428 VCC.n449 VCC 0.535293
R8429 VCC.n1001 VCC 0.535293
R8430 VCC.n1559 VCC 0.535293
R8431 VCC.n2110 VCC 0.535293
R8432 VCC.n2668 VCC 0.535293
R8433 VCC.n3219 VCC 0.535293
R8434 VCC.n3777 VCC 0.535293
R8435 VCC.n4328 VCC 0.535293
R8436 VCC.n4886 VCC 0.535293
R8437 VCC.n5437 VCC 0.535293
R8438 VCC.n5994 VCC 0.535293
R8439 VCC.n6544 VCC 0.535293
R8440 VCC.n7101 VCC 0.535293
R8441 VCC.n7651 VCC 0.535293
R8442 VCC.n8208 VCC 0.535293
R8443 VCC.n8571 VCC 0.535293
R8444 VCC.n549 VCC.n3 0.507747
R8445 VCC.n1103 VCC.n557 0.507747
R8446 VCC.n1657 VCC.n1656 0.507747
R8447 VCC.n2212 VCC.n1666 0.507747
R8448 VCC.n2766 VCC.n2765 0.507747
R8449 VCC.n3321 VCC.n2775 0.507747
R8450 VCC.n3875 VCC.n3874 0.507747
R8451 VCC.n4430 VCC.n3884 0.507747
R8452 VCC.n4984 VCC.n4983 0.507747
R8453 VCC.n5539 VCC.n4993 0.507747
R8454 VCC.n6092 VCC.n6091 0.507747
R8455 VCC.n6646 VCC.n6100 0.507747
R8456 VCC.n7199 VCC.n7198 0.507747
R8457 VCC.n7753 VCC.n7207 0.507747
R8458 VCC.n8306 VCC.n8305 0.507747
R8459 VCC.n8673 VCC.n8314 0.507747
R8460 VCC.n1532 VCC.n1174 0.465127
R8461 VCC.n2641 VCC.n2283 0.465127
R8462 VCC.n3750 VCC.n3392 0.465127
R8463 VCC.n4859 VCC.n4501 0.465127
R8464 VCC.n5967 VCC.n5609 0.465127
R8465 VCC.n7074 VCC.n6716 0.465127
R8466 VCC.n8181 VCC.n7823 0.465127
R8467 VCC.n422 VCC.n65 0.465115
R8468 VCC.n974 VCC.n617 0.465115
R8469 VCC.n2083 VCC.n1726 0.465115
R8470 VCC.n3192 VCC.n2835 0.465115
R8471 VCC.n4301 VCC.n3944 0.465115
R8472 VCC.n5410 VCC.n5053 0.465115
R8473 VCC.n6517 VCC.n6160 0.465115
R8474 VCC.n7624 VCC.n7267 0.465115
R8475 VCC.n8544 VCC.n8374 0.465115
R8476 VCC.n249 VCC.n248 0.366214
R8477 VCC.n468 VCC.n54 0.366214
R8478 VCC.n531 VCC.n529 0.366214
R8479 VCC.n801 VCC.n800 0.366214
R8480 VCC.n1020 VCC.n606 0.366214
R8481 VCC.n1083 VCC.n1081 0.366214
R8482 VCC.n1578 VCC.n1577 0.366214
R8483 VCC.n1649 VCC.n1648 0.366214
R8484 VCC.n1359 VCC.n1358 0.366214
R8485 VCC.n1910 VCC.n1909 0.366214
R8486 VCC.n2129 VCC.n1715 0.366214
R8487 VCC.n2192 VCC.n2190 0.366214
R8488 VCC.n2687 VCC.n2686 0.366214
R8489 VCC.n2758 VCC.n2757 0.366214
R8490 VCC.n2468 VCC.n2467 0.366214
R8491 VCC.n3019 VCC.n3018 0.366214
R8492 VCC.n3238 VCC.n2824 0.366214
R8493 VCC.n3301 VCC.n3299 0.366214
R8494 VCC.n3796 VCC.n3795 0.366214
R8495 VCC.n3867 VCC.n3866 0.366214
R8496 VCC.n3577 VCC.n3576 0.366214
R8497 VCC.n4128 VCC.n4127 0.366214
R8498 VCC.n4347 VCC.n3933 0.366214
R8499 VCC.n4410 VCC.n4408 0.366214
R8500 VCC.n4905 VCC.n4904 0.366214
R8501 VCC.n4976 VCC.n4975 0.366214
R8502 VCC.n4686 VCC.n4685 0.366214
R8503 VCC.n5237 VCC.n5236 0.366214
R8504 VCC.n5456 VCC.n5042 0.366214
R8505 VCC.n5519 VCC.n5517 0.366214
R8506 VCC.n6013 VCC.n6012 0.366214
R8507 VCC.n6084 VCC.n6083 0.366214
R8508 VCC.n5794 VCC.n5793 0.366214
R8509 VCC.n6344 VCC.n6343 0.366214
R8510 VCC.n6563 VCC.n6149 0.366214
R8511 VCC.n6626 VCC.n6624 0.366214
R8512 VCC.n7120 VCC.n7119 0.366214
R8513 VCC.n7191 VCC.n7190 0.366214
R8514 VCC.n6901 VCC.n6900 0.366214
R8515 VCC.n7451 VCC.n7450 0.366214
R8516 VCC.n7670 VCC.n7256 0.366214
R8517 VCC.n7733 VCC.n7731 0.366214
R8518 VCC.n8227 VCC.n8226 0.366214
R8519 VCC.n8298 VCC.n8297 0.366214
R8520 VCC.n8008 VCC.n8007 0.366214
R8521 VCC.n8590 VCC.n8363 0.366214
R8522 VCC.n8653 VCC.n8651 0.366214
R8523 VCC VCC.n553 0.338784
R8524 VCC VCC.n2771 0.338735
R8525 VCC VCC.n4989 0.338735
R8526 VCC.n8679 VCC 0.338735
R8527 VCC.n2771 VCC 0.309324
R8528 VCC VCC.n8679 0.309324
R8529 VCC VCC.n552 0.300964
R8530 VCC VCC.n1106 0.300964
R8531 VCC VCC.n1660 0.300964
R8532 VCC VCC.n2215 0.300964
R8533 VCC VCC.n2769 0.300964
R8534 VCC VCC.n3324 0.300964
R8535 VCC VCC.n3878 0.300964
R8536 VCC VCC.n4433 0.300964
R8537 VCC VCC.n4987 0.300964
R8538 VCC VCC.n5542 0.300964
R8539 VCC VCC.n6095 0.300964
R8540 VCC VCC.n6649 0.300964
R8541 VCC VCC.n7202 0.300964
R8542 VCC VCC.n7756 0.300964
R8543 VCC VCC.n8309 0.300964
R8544 VCC VCC.n8676 0.300964
R8545 VCC.n191 VCC 0.294921
R8546 VCC.n743 VCC 0.294921
R8547 VCC.n1301 VCC 0.294921
R8548 VCC.n1852 VCC 0.294921
R8549 VCC.n2410 VCC 0.294921
R8550 VCC.n2961 VCC 0.294921
R8551 VCC.n3519 VCC 0.294921
R8552 VCC.n4070 VCC 0.294921
R8553 VCC.n4628 VCC 0.294921
R8554 VCC.n5179 VCC 0.294921
R8555 VCC.n5736 VCC 0.294921
R8556 VCC.n6286 VCC 0.294921
R8557 VCC.n6843 VCC 0.294921
R8558 VCC.n7393 VCC 0.294921
R8559 VCC.n7950 VCC 0.294921
R8560 VCC.n8437 VCC 0.294921
R8561 VCC.n315 VCC 0.287536
R8562 VCC.n867 VCC 0.287536
R8563 VCC.n1425 VCC 0.287536
R8564 VCC.n1976 VCC 0.287536
R8565 VCC.n2534 VCC 0.287536
R8566 VCC.n3085 VCC 0.287536
R8567 VCC.n3643 VCC 0.287536
R8568 VCC.n4194 VCC 0.287536
R8569 VCC.n4752 VCC 0.287536
R8570 VCC.n5303 VCC 0.287536
R8571 VCC.n5860 VCC 0.287536
R8572 VCC.n6410 VCC 0.287536
R8573 VCC.n6967 VCC 0.287536
R8574 VCC.n7517 VCC 0.287536
R8575 VCC.n8074 VCC 0.287536
R8576 VCC.n224 VCC.n183 0.274786
R8577 VCC.n286 VCC.n141 0.274786
R8578 VCC.n339 VCC.n118 0.274786
R8579 VCC.n365 VCC.n97 0.274786
R8580 VCC.n387 VCC.n95 0.274786
R8581 VCC.n415 VCC.n414 0.274786
R8582 VCC.n776 VCC.n735 0.274786
R8583 VCC.n838 VCC.n693 0.274786
R8584 VCC.n891 VCC.n670 0.274786
R8585 VCC.n917 VCC.n649 0.274786
R8586 VCC.n939 VCC.n647 0.274786
R8587 VCC.n967 VCC.n966 0.274786
R8588 VCC.n1448 VCC.n1227 0.274786
R8589 VCC.n1474 VCC.n1206 0.274786
R8590 VCC.n1496 VCC.n1204 0.274786
R8591 VCC.n1524 VCC.n1523 0.274786
R8592 VCC.n1334 VCC.n1293 0.274786
R8593 VCC.n1396 VCC.n1251 0.274786
R8594 VCC.n1885 VCC.n1844 0.274786
R8595 VCC.n1947 VCC.n1802 0.274786
R8596 VCC.n2000 VCC.n1779 0.274786
R8597 VCC.n2026 VCC.n1758 0.274786
R8598 VCC.n2048 VCC.n1756 0.274786
R8599 VCC.n2076 VCC.n2075 0.274786
R8600 VCC.n2557 VCC.n2336 0.274786
R8601 VCC.n2583 VCC.n2315 0.274786
R8602 VCC.n2605 VCC.n2313 0.274786
R8603 VCC.n2633 VCC.n2632 0.274786
R8604 VCC.n2443 VCC.n2402 0.274786
R8605 VCC.n2505 VCC.n2360 0.274786
R8606 VCC.n2994 VCC.n2953 0.274786
R8607 VCC.n3056 VCC.n2911 0.274786
R8608 VCC.n3109 VCC.n2888 0.274786
R8609 VCC.n3135 VCC.n2867 0.274786
R8610 VCC.n3157 VCC.n2865 0.274786
R8611 VCC.n3185 VCC.n3184 0.274786
R8612 VCC.n3666 VCC.n3445 0.274786
R8613 VCC.n3692 VCC.n3424 0.274786
R8614 VCC.n3714 VCC.n3422 0.274786
R8615 VCC.n3742 VCC.n3741 0.274786
R8616 VCC.n3552 VCC.n3511 0.274786
R8617 VCC.n3614 VCC.n3469 0.274786
R8618 VCC.n4103 VCC.n4062 0.274786
R8619 VCC.n4165 VCC.n4020 0.274786
R8620 VCC.n4218 VCC.n3997 0.274786
R8621 VCC.n4244 VCC.n3976 0.274786
R8622 VCC.n4266 VCC.n3974 0.274786
R8623 VCC.n4294 VCC.n4293 0.274786
R8624 VCC.n4775 VCC.n4554 0.274786
R8625 VCC.n4801 VCC.n4533 0.274786
R8626 VCC.n4823 VCC.n4531 0.274786
R8627 VCC.n4851 VCC.n4850 0.274786
R8628 VCC.n4661 VCC.n4620 0.274786
R8629 VCC.n4723 VCC.n4578 0.274786
R8630 VCC.n5212 VCC.n5171 0.274786
R8631 VCC.n5274 VCC.n5129 0.274786
R8632 VCC.n5327 VCC.n5106 0.274786
R8633 VCC.n5353 VCC.n5085 0.274786
R8634 VCC.n5375 VCC.n5083 0.274786
R8635 VCC.n5403 VCC.n5402 0.274786
R8636 VCC.n5883 VCC.n5662 0.274786
R8637 VCC.n5909 VCC.n5641 0.274786
R8638 VCC.n5931 VCC.n5639 0.274786
R8639 VCC.n5959 VCC.n5958 0.274786
R8640 VCC.n5769 VCC.n5728 0.274786
R8641 VCC.n5831 VCC.n5686 0.274786
R8642 VCC.n6319 VCC.n6278 0.274786
R8643 VCC.n6381 VCC.n6236 0.274786
R8644 VCC.n6434 VCC.n6213 0.274786
R8645 VCC.n6460 VCC.n6192 0.274786
R8646 VCC.n6482 VCC.n6190 0.274786
R8647 VCC.n6510 VCC.n6509 0.274786
R8648 VCC.n6990 VCC.n6769 0.274786
R8649 VCC.n7016 VCC.n6748 0.274786
R8650 VCC.n7038 VCC.n6746 0.274786
R8651 VCC.n7066 VCC.n7065 0.274786
R8652 VCC.n6876 VCC.n6835 0.274786
R8653 VCC.n6938 VCC.n6793 0.274786
R8654 VCC.n7426 VCC.n7385 0.274786
R8655 VCC.n7488 VCC.n7343 0.274786
R8656 VCC.n7541 VCC.n7320 0.274786
R8657 VCC.n7567 VCC.n7299 0.274786
R8658 VCC.n7589 VCC.n7297 0.274786
R8659 VCC.n7617 VCC.n7616 0.274786
R8660 VCC.n8097 VCC.n7876 0.274786
R8661 VCC.n8123 VCC.n7855 0.274786
R8662 VCC.n8145 VCC.n7853 0.274786
R8663 VCC.n8173 VCC.n8172 0.274786
R8664 VCC.n7983 VCC.n7942 0.274786
R8665 VCC.n8045 VCC.n7900 0.274786
R8666 VCC.n8461 VCC.n8427 0.274786
R8667 VCC.n8487 VCC.n8406 0.274786
R8668 VCC.n8509 VCC.n8404 0.274786
R8669 VCC.n8537 VCC.n8536 0.274786
R8670 VCC VCC.n313 0.213679
R8671 VCC VCC.n865 0.213679
R8672 VCC VCC.n1423 0.213679
R8673 VCC VCC.n1974 0.213679
R8674 VCC VCC.n2532 0.213679
R8675 VCC VCC.n3083 0.213679
R8676 VCC VCC.n3641 0.213679
R8677 VCC VCC.n4192 0.213679
R8678 VCC VCC.n4750 0.213679
R8679 VCC VCC.n5301 0.213679
R8680 VCC VCC.n5858 0.213679
R8681 VCC VCC.n6408 0.213679
R8682 VCC VCC.n6965 0.213679
R8683 VCC VCC.n7515 0.213679
R8684 VCC VCC.n8072 0.213679
R8685 VCC.n160 VCC.n156 0.183357
R8686 VCC.n490 VCC.n43 0.183357
R8687 VCC.n491 VCC.n490 0.183357
R8688 VCC.n523 VCC.n24 0.183357
R8689 VCC.n523 VCC.n25 0.183357
R8690 VCC.n712 VCC.n708 0.183357
R8691 VCC.n1042 VCC.n595 0.183357
R8692 VCC.n1043 VCC.n1042 0.183357
R8693 VCC.n1075 VCC.n576 0.183357
R8694 VCC.n1075 VCC.n577 0.183357
R8695 VCC.n1593 VCC.n1587 0.183357
R8696 VCC.n1587 VCC.n1160 0.183357
R8697 VCC.n1623 VCC.n1135 0.183357
R8698 VCC.n1623 VCC.n1141 0.183357
R8699 VCC.n1270 VCC.n1266 0.183357
R8700 VCC.n1821 VCC.n1817 0.183357
R8701 VCC.n2151 VCC.n1704 0.183357
R8702 VCC.n2152 VCC.n2151 0.183357
R8703 VCC.n2184 VCC.n1685 0.183357
R8704 VCC.n2184 VCC.n1686 0.183357
R8705 VCC.n2702 VCC.n2696 0.183357
R8706 VCC.n2696 VCC.n2269 0.183357
R8707 VCC.n2732 VCC.n2244 0.183357
R8708 VCC.n2732 VCC.n2250 0.183357
R8709 VCC.n2379 VCC.n2375 0.183357
R8710 VCC.n2930 VCC.n2926 0.183357
R8711 VCC.n3260 VCC.n2813 0.183357
R8712 VCC.n3261 VCC.n3260 0.183357
R8713 VCC.n3293 VCC.n2794 0.183357
R8714 VCC.n3293 VCC.n2795 0.183357
R8715 VCC.n3811 VCC.n3805 0.183357
R8716 VCC.n3805 VCC.n3378 0.183357
R8717 VCC.n3841 VCC.n3353 0.183357
R8718 VCC.n3841 VCC.n3359 0.183357
R8719 VCC.n3488 VCC.n3484 0.183357
R8720 VCC.n4039 VCC.n4035 0.183357
R8721 VCC.n4369 VCC.n3922 0.183357
R8722 VCC.n4370 VCC.n4369 0.183357
R8723 VCC.n4402 VCC.n3903 0.183357
R8724 VCC.n4402 VCC.n3904 0.183357
R8725 VCC.n4920 VCC.n4914 0.183357
R8726 VCC.n4914 VCC.n4487 0.183357
R8727 VCC.n4950 VCC.n4462 0.183357
R8728 VCC.n4950 VCC.n4468 0.183357
R8729 VCC.n4597 VCC.n4593 0.183357
R8730 VCC.n5148 VCC.n5144 0.183357
R8731 VCC.n5478 VCC.n5031 0.183357
R8732 VCC.n5479 VCC.n5478 0.183357
R8733 VCC.n5511 VCC.n5012 0.183357
R8734 VCC.n5511 VCC.n5013 0.183357
R8735 VCC.n6028 VCC.n6022 0.183357
R8736 VCC.n6022 VCC.n5595 0.183357
R8737 VCC.n6058 VCC.n5570 0.183357
R8738 VCC.n6058 VCC.n5576 0.183357
R8739 VCC.n5705 VCC.n5701 0.183357
R8740 VCC.n6255 VCC.n6251 0.183357
R8741 VCC.n6585 VCC.n6138 0.183357
R8742 VCC.n6586 VCC.n6585 0.183357
R8743 VCC.n6618 VCC.n6119 0.183357
R8744 VCC.n6618 VCC.n6120 0.183357
R8745 VCC.n7135 VCC.n7129 0.183357
R8746 VCC.n7129 VCC.n6702 0.183357
R8747 VCC.n7165 VCC.n6677 0.183357
R8748 VCC.n7165 VCC.n6683 0.183357
R8749 VCC.n6812 VCC.n6808 0.183357
R8750 VCC.n7362 VCC.n7358 0.183357
R8751 VCC.n7692 VCC.n7245 0.183357
R8752 VCC.n7693 VCC.n7692 0.183357
R8753 VCC.n7725 VCC.n7226 0.183357
R8754 VCC.n7725 VCC.n7227 0.183357
R8755 VCC.n8242 VCC.n8236 0.183357
R8756 VCC.n8236 VCC.n7809 0.183357
R8757 VCC.n8272 VCC.n7784 0.183357
R8758 VCC.n8272 VCC.n7790 0.183357
R8759 VCC.n7919 VCC.n7915 0.183357
R8760 VCC.n8612 VCC.n8352 0.183357
R8761 VCC.n8613 VCC.n8612 0.183357
R8762 VCC.n8645 VCC.n8333 0.183357
R8763 VCC.n8645 VCC.n8334 0.183357
R8764 VCC VCC.n448 0.114307
R8765 VCC VCC.n1000 0.114307
R8766 VCC VCC.n1558 0.114307
R8767 VCC VCC.n2109 0.114307
R8768 VCC VCC.n2667 0.114307
R8769 VCC VCC.n3218 0.114307
R8770 VCC VCC.n3776 0.114307
R8771 VCC VCC.n4327 0.114307
R8772 VCC VCC.n4885 0.114307
R8773 VCC VCC.n5436 0.114307
R8774 VCC VCC.n5993 0.114307
R8775 VCC VCC.n6543 0.114307
R8776 VCC VCC.n7100 0.114307
R8777 VCC VCC.n7650 0.114307
R8778 VCC VCC.n8207 0.114307
R8779 VCC VCC.n8570 0.114307
R8780 VCC.n231 VCC.n178 0.0919286
R8781 VCC.n271 VCC.n270 0.0919286
R8782 VCC.n358 VCC.n106 0.0919286
R8783 VCC.n398 VCC.n91 0.0919286
R8784 VCC.n531 VCC.n530 0.0919286
R8785 VCC.n544 VCC.n7 0.0919286
R8786 VCC.n783 VCC.n730 0.0919286
R8787 VCC.n823 VCC.n822 0.0919286
R8788 VCC.n910 VCC.n658 0.0919286
R8789 VCC.n950 VCC.n643 0.0919286
R8790 VCC.n1083 VCC.n1082 0.0919286
R8791 VCC.n1098 VCC.n561 0.0919286
R8792 VCC.n1648 VCC.n1117 0.0919286
R8793 VCC.n1124 VCC.n1123 0.0919286
R8794 VCC.n1467 VCC.n1215 0.0919286
R8795 VCC.n1507 VCC.n1200 0.0919286
R8796 VCC.n1341 VCC.n1288 0.0919286
R8797 VCC.n1381 VCC.n1380 0.0919286
R8798 VCC.n1892 VCC.n1839 0.0919286
R8799 VCC.n1932 VCC.n1931 0.0919286
R8800 VCC.n2019 VCC.n1767 0.0919286
R8801 VCC.n2059 VCC.n1752 0.0919286
R8802 VCC.n2192 VCC.n2191 0.0919286
R8803 VCC.n2207 VCC.n1670 0.0919286
R8804 VCC.n2757 VCC.n2226 0.0919286
R8805 VCC.n2233 VCC.n2232 0.0919286
R8806 VCC.n2576 VCC.n2324 0.0919286
R8807 VCC.n2616 VCC.n2309 0.0919286
R8808 VCC.n2450 VCC.n2397 0.0919286
R8809 VCC.n2490 VCC.n2489 0.0919286
R8810 VCC.n3001 VCC.n2948 0.0919286
R8811 VCC.n3041 VCC.n3040 0.0919286
R8812 VCC.n3128 VCC.n2876 0.0919286
R8813 VCC.n3168 VCC.n2861 0.0919286
R8814 VCC.n3301 VCC.n3300 0.0919286
R8815 VCC.n3316 VCC.n2779 0.0919286
R8816 VCC.n3866 VCC.n3335 0.0919286
R8817 VCC.n3342 VCC.n3341 0.0919286
R8818 VCC.n3685 VCC.n3433 0.0919286
R8819 VCC.n3725 VCC.n3418 0.0919286
R8820 VCC.n3559 VCC.n3506 0.0919286
R8821 VCC.n3599 VCC.n3598 0.0919286
R8822 VCC.n4110 VCC.n4057 0.0919286
R8823 VCC.n4150 VCC.n4149 0.0919286
R8824 VCC.n4237 VCC.n3985 0.0919286
R8825 VCC.n4277 VCC.n3970 0.0919286
R8826 VCC.n4410 VCC.n4409 0.0919286
R8827 VCC.n4425 VCC.n3888 0.0919286
R8828 VCC.n4975 VCC.n4444 0.0919286
R8829 VCC.n4451 VCC.n4450 0.0919286
R8830 VCC.n4794 VCC.n4542 0.0919286
R8831 VCC.n4834 VCC.n4527 0.0919286
R8832 VCC.n4668 VCC.n4615 0.0919286
R8833 VCC.n4708 VCC.n4707 0.0919286
R8834 VCC.n5219 VCC.n5166 0.0919286
R8835 VCC.n5259 VCC.n5258 0.0919286
R8836 VCC.n5346 VCC.n5094 0.0919286
R8837 VCC.n5386 VCC.n5079 0.0919286
R8838 VCC.n5519 VCC.n5518 0.0919286
R8839 VCC.n5534 VCC.n4997 0.0919286
R8840 VCC.n6083 VCC.n5552 0.0919286
R8841 VCC.n5559 VCC.n5558 0.0919286
R8842 VCC.n5902 VCC.n5650 0.0919286
R8843 VCC.n5942 VCC.n5635 0.0919286
R8844 VCC.n5776 VCC.n5723 0.0919286
R8845 VCC.n5816 VCC.n5815 0.0919286
R8846 VCC.n6326 VCC.n6273 0.0919286
R8847 VCC.n6366 VCC.n6365 0.0919286
R8848 VCC.n6453 VCC.n6201 0.0919286
R8849 VCC.n6493 VCC.n6186 0.0919286
R8850 VCC.n6626 VCC.n6625 0.0919286
R8851 VCC.n6641 VCC.n6104 0.0919286
R8852 VCC.n7190 VCC.n6659 0.0919286
R8853 VCC.n6666 VCC.n6665 0.0919286
R8854 VCC.n7009 VCC.n6757 0.0919286
R8855 VCC.n7049 VCC.n6742 0.0919286
R8856 VCC.n6883 VCC.n6830 0.0919286
R8857 VCC.n6923 VCC.n6922 0.0919286
R8858 VCC.n7433 VCC.n7380 0.0919286
R8859 VCC.n7473 VCC.n7472 0.0919286
R8860 VCC.n7560 VCC.n7308 0.0919286
R8861 VCC.n7600 VCC.n7293 0.0919286
R8862 VCC.n7733 VCC.n7732 0.0919286
R8863 VCC.n7748 VCC.n7211 0.0919286
R8864 VCC.n8297 VCC.n7766 0.0919286
R8865 VCC.n7773 VCC.n7772 0.0919286
R8866 VCC.n8116 VCC.n7864 0.0919286
R8867 VCC.n8156 VCC.n7849 0.0919286
R8868 VCC.n7990 VCC.n7937 0.0919286
R8869 VCC.n8030 VCC.n8029 0.0919286
R8870 VCC.n8480 VCC.n8415 0.0919286
R8871 VCC.n8520 VCC.n8400 0.0919286
R8872 VCC.n8653 VCC.n8652 0.0919286
R8873 VCC.n8668 VCC.n8318 0.0919286
R8874 VCC.n1107 VCC 0.0247197
R8875 VCC.n2216 VCC 0.0247197
R8876 VCC.n3325 VCC 0.0247197
R8877 VCC.n4434 VCC 0.0247197
R8878 VCC.n8682 VCC 0.0247197
R8879 VCC.n8680 VCC 0.0247197
R8880 VCC.n8678 VCC 0.0247197
R8881 VCC.n553 VCC 0.0246714
R8882 VCC.n1661 VCC 0.0246714
R8883 VCC.n2770 VCC 0.0246714
R8884 VCC.n3879 VCC 0.0246714
R8885 VCC.n4988 VCC 0.0246714
R8886 VCC.n6096 VCC 0.0246714
R8887 VCC.n7203 VCC 0.0246714
R8888 VCC.n8310 VCC 0.0246714
R8889 VCC.n218 VCC.n217 0.024
R8890 VCC.n308 VCC.n307 0.024
R8891 VCC.n317 VCC.n114 0.024
R8892 VCC.n443 VCC.n442 0.024
R8893 VCC.n461 VCC.n460 0.024
R8894 VCC.n537 VCC.n536 0.024
R8895 VCC.n770 VCC.n769 0.024
R8896 VCC.n860 VCC.n859 0.024
R8897 VCC.n869 VCC.n666 0.024
R8898 VCC.n995 VCC.n994 0.024
R8899 VCC.n1013 VCC.n1012 0.024
R8900 VCC.n1089 VCC.n1088 0.024
R8901 VCC.n1328 VCC.n1327 0.024
R8902 VCC.n1418 VCC.n1417 0.024
R8903 VCC.n1427 VCC.n1223 0.024
R8904 VCC.n1553 VCC.n1552 0.024
R8905 VCC.n1572 VCC.n1571 0.024
R8906 VCC.n1636 VCC.n1635 0.024
R8907 VCC.n1879 VCC.n1878 0.024
R8908 VCC.n1969 VCC.n1968 0.024
R8909 VCC.n1978 VCC.n1775 0.024
R8910 VCC.n2104 VCC.n2103 0.024
R8911 VCC.n2122 VCC.n2121 0.024
R8912 VCC.n2198 VCC.n2197 0.024
R8913 VCC.n2437 VCC.n2436 0.024
R8914 VCC.n2527 VCC.n2526 0.024
R8915 VCC.n2536 VCC.n2332 0.024
R8916 VCC.n2662 VCC.n2661 0.024
R8917 VCC.n2681 VCC.n2680 0.024
R8918 VCC.n2745 VCC.n2744 0.024
R8919 VCC.n2988 VCC.n2987 0.024
R8920 VCC.n3078 VCC.n3077 0.024
R8921 VCC.n3087 VCC.n2884 0.024
R8922 VCC.n3213 VCC.n3212 0.024
R8923 VCC.n3231 VCC.n3230 0.024
R8924 VCC.n3307 VCC.n3306 0.024
R8925 VCC.n3546 VCC.n3545 0.024
R8926 VCC.n3636 VCC.n3635 0.024
R8927 VCC.n3645 VCC.n3441 0.024
R8928 VCC.n3771 VCC.n3770 0.024
R8929 VCC.n3790 VCC.n3789 0.024
R8930 VCC.n3854 VCC.n3853 0.024
R8931 VCC.n4097 VCC.n4096 0.024
R8932 VCC.n4187 VCC.n4186 0.024
R8933 VCC.n4196 VCC.n3993 0.024
R8934 VCC.n4322 VCC.n4321 0.024
R8935 VCC.n4340 VCC.n4339 0.024
R8936 VCC.n4416 VCC.n4415 0.024
R8937 VCC.n4655 VCC.n4654 0.024
R8938 VCC.n4745 VCC.n4744 0.024
R8939 VCC.n4754 VCC.n4550 0.024
R8940 VCC.n4880 VCC.n4879 0.024
R8941 VCC.n4899 VCC.n4898 0.024
R8942 VCC.n4963 VCC.n4962 0.024
R8943 VCC.n5206 VCC.n5205 0.024
R8944 VCC.n5296 VCC.n5295 0.024
R8945 VCC.n5305 VCC.n5102 0.024
R8946 VCC.n5431 VCC.n5430 0.024
R8947 VCC.n5449 VCC.n5448 0.024
R8948 VCC.n5525 VCC.n5524 0.024
R8949 VCC.n5763 VCC.n5762 0.024
R8950 VCC.n5853 VCC.n5852 0.024
R8951 VCC.n5862 VCC.n5658 0.024
R8952 VCC.n5988 VCC.n5987 0.024
R8953 VCC.n6007 VCC.n6006 0.024
R8954 VCC.n6071 VCC.n6070 0.024
R8955 VCC.n6313 VCC.n6312 0.024
R8956 VCC.n6403 VCC.n6402 0.024
R8957 VCC.n6412 VCC.n6209 0.024
R8958 VCC.n6538 VCC.n6537 0.024
R8959 VCC.n6556 VCC.n6555 0.024
R8960 VCC.n6632 VCC.n6631 0.024
R8961 VCC.n6870 VCC.n6869 0.024
R8962 VCC.n6960 VCC.n6959 0.024
R8963 VCC.n6969 VCC.n6765 0.024
R8964 VCC.n7095 VCC.n7094 0.024
R8965 VCC.n7114 VCC.n7113 0.024
R8966 VCC.n7178 VCC.n7177 0.024
R8967 VCC.n7420 VCC.n7419 0.024
R8968 VCC.n7510 VCC.n7509 0.024
R8969 VCC.n7519 VCC.n7316 0.024
R8970 VCC.n7645 VCC.n7644 0.024
R8971 VCC.n7663 VCC.n7662 0.024
R8972 VCC.n7739 VCC.n7738 0.024
R8973 VCC.n7977 VCC.n7976 0.024
R8974 VCC.n8067 VCC.n8066 0.024
R8975 VCC.n8076 VCC.n7872 0.024
R8976 VCC.n8202 VCC.n8201 0.024
R8977 VCC.n8221 VCC.n8220 0.024
R8978 VCC.n8285 VCC.n8284 0.024
R8979 VCC.n8439 VCC.n8423 0.024
R8980 VCC.n8565 VCC.n8564 0.024
R8981 VCC.n8583 VCC.n8582 0.024
R8982 VCC.n8659 VCC.n8658 0.024
R8983 VCC.n47 VCC.n38 0.0228214
R8984 VCC.n509 VCC.n508 0.0228214
R8985 VCC.n517 VCC.n16 0.0228214
R8986 VCC.n599 VCC.n590 0.0228214
R8987 VCC.n1061 VCC.n1060 0.0228214
R8988 VCC.n1069 VCC.n568 0.0228214
R8989 VCC.n1605 VCC.n1604 0.0228214
R8990 VCC.n1148 VCC.n1133 0.0228214
R8991 VCC.n1632 VCC.n1128 0.0228214
R8992 VCC.n1708 VCC.n1699 0.0228214
R8993 VCC.n2170 VCC.n2169 0.0228214
R8994 VCC.n2178 VCC.n1677 0.0228214
R8995 VCC.n2714 VCC.n2713 0.0228214
R8996 VCC.n2257 VCC.n2242 0.0228214
R8997 VCC.n2741 VCC.n2237 0.0228214
R8998 VCC.n2817 VCC.n2808 0.0228214
R8999 VCC.n3279 VCC.n3278 0.0228214
R9000 VCC.n3287 VCC.n2786 0.0228214
R9001 VCC.n3823 VCC.n3822 0.0228214
R9002 VCC.n3366 VCC.n3351 0.0228214
R9003 VCC.n3850 VCC.n3346 0.0228214
R9004 VCC.n3926 VCC.n3917 0.0228214
R9005 VCC.n4388 VCC.n4387 0.0228214
R9006 VCC.n4396 VCC.n3895 0.0228214
R9007 VCC.n4932 VCC.n4931 0.0228214
R9008 VCC.n4475 VCC.n4460 0.0228214
R9009 VCC.n4959 VCC.n4455 0.0228214
R9010 VCC.n5035 VCC.n5026 0.0228214
R9011 VCC.n5497 VCC.n5496 0.0228214
R9012 VCC.n5505 VCC.n5004 0.0228214
R9013 VCC.n6040 VCC.n6039 0.0228214
R9014 VCC.n5583 VCC.n5568 0.0228214
R9015 VCC.n6067 VCC.n5563 0.0228214
R9016 VCC.n6142 VCC.n6133 0.0228214
R9017 VCC.n6604 VCC.n6603 0.0228214
R9018 VCC.n6612 VCC.n6111 0.0228214
R9019 VCC.n7147 VCC.n7146 0.0228214
R9020 VCC.n6690 VCC.n6675 0.0228214
R9021 VCC.n7174 VCC.n6670 0.0228214
R9022 VCC.n7249 VCC.n7240 0.0228214
R9023 VCC.n7711 VCC.n7710 0.0228214
R9024 VCC.n7719 VCC.n7218 0.0228214
R9025 VCC.n8254 VCC.n8253 0.0228214
R9026 VCC.n7797 VCC.n7782 0.0228214
R9027 VCC.n8281 VCC.n7777 0.0228214
R9028 VCC.n8356 VCC.n8347 0.0228214
R9029 VCC.n8631 VCC.n8630 0.0228214
R9030 VCC.n8639 VCC.n8325 0.0228214
R9031 VCC.n553 VCC 0.0199714
R9032 VCC.n1661 VCC 0.0199714
R9033 VCC.n2770 VCC 0.0199714
R9034 VCC.n3879 VCC 0.0199714
R9035 VCC.n4988 VCC 0.0199714
R9036 VCC.n6096 VCC 0.0199714
R9037 VCC.n7203 VCC 0.0199714
R9038 VCC.n8310 VCC 0.0199714
R9039 VCC.n253 VCC.n157 0.0174643
R9040 VCC.n252 VCC.n163 0.0174643
R9041 VCC.n376 VCC.n99 0.0174643
R9042 VCC.n377 VCC.n376 0.0174643
R9043 VCC.n381 VCC.n101 0.0174643
R9044 VCC.n378 VCC.n101 0.0174643
R9045 VCC.n501 VCC.n500 0.0174643
R9046 VCC.n500 VCC.n32 0.0174643
R9047 VCC.n502 VCC.n37 0.0174643
R9048 VCC.n37 VCC.n33 0.0174643
R9049 VCC.n805 VCC.n709 0.0174643
R9050 VCC.n804 VCC.n715 0.0174643
R9051 VCC.n928 VCC.n651 0.0174643
R9052 VCC.n929 VCC.n928 0.0174643
R9053 VCC.n933 VCC.n653 0.0174643
R9054 VCC.n930 VCC.n653 0.0174643
R9055 VCC.n1053 VCC.n1052 0.0174643
R9056 VCC.n1052 VCC.n584 0.0174643
R9057 VCC.n1054 VCC.n589 0.0174643
R9058 VCC.n589 VCC.n585 0.0174643
R9059 VCC.n1615 VCC.n1146 0.0174643
R9060 VCC.n1615 VCC.n1614 0.0174643
R9061 VCC.n1607 VCC.n1147 0.0174643
R9062 VCC.n1613 VCC.n1147 0.0174643
R9063 VCC.n1485 VCC.n1208 0.0174643
R9064 VCC.n1486 VCC.n1485 0.0174643
R9065 VCC.n1490 VCC.n1210 0.0174643
R9066 VCC.n1487 VCC.n1210 0.0174643
R9067 VCC.n1363 VCC.n1267 0.0174643
R9068 VCC.n1362 VCC.n1273 0.0174643
R9069 VCC.n1914 VCC.n1818 0.0174643
R9070 VCC.n1913 VCC.n1824 0.0174643
R9071 VCC.n2037 VCC.n1760 0.0174643
R9072 VCC.n2038 VCC.n2037 0.0174643
R9073 VCC.n2042 VCC.n1762 0.0174643
R9074 VCC.n2039 VCC.n1762 0.0174643
R9075 VCC.n2162 VCC.n2161 0.0174643
R9076 VCC.n2161 VCC.n1693 0.0174643
R9077 VCC.n2163 VCC.n1698 0.0174643
R9078 VCC.n1698 VCC.n1694 0.0174643
R9079 VCC.n2724 VCC.n2255 0.0174643
R9080 VCC.n2724 VCC.n2723 0.0174643
R9081 VCC.n2716 VCC.n2256 0.0174643
R9082 VCC.n2722 VCC.n2256 0.0174643
R9083 VCC.n2594 VCC.n2317 0.0174643
R9084 VCC.n2595 VCC.n2594 0.0174643
R9085 VCC.n2599 VCC.n2319 0.0174643
R9086 VCC.n2596 VCC.n2319 0.0174643
R9087 VCC.n2472 VCC.n2376 0.0174643
R9088 VCC.n2471 VCC.n2382 0.0174643
R9089 VCC.n3023 VCC.n2927 0.0174643
R9090 VCC.n3022 VCC.n2933 0.0174643
R9091 VCC.n3146 VCC.n2869 0.0174643
R9092 VCC.n3147 VCC.n3146 0.0174643
R9093 VCC.n3151 VCC.n2871 0.0174643
R9094 VCC.n3148 VCC.n2871 0.0174643
R9095 VCC.n3271 VCC.n3270 0.0174643
R9096 VCC.n3270 VCC.n2802 0.0174643
R9097 VCC.n3272 VCC.n2807 0.0174643
R9098 VCC.n2807 VCC.n2803 0.0174643
R9099 VCC.n3833 VCC.n3364 0.0174643
R9100 VCC.n3833 VCC.n3832 0.0174643
R9101 VCC.n3825 VCC.n3365 0.0174643
R9102 VCC.n3831 VCC.n3365 0.0174643
R9103 VCC.n3703 VCC.n3426 0.0174643
R9104 VCC.n3704 VCC.n3703 0.0174643
R9105 VCC.n3708 VCC.n3428 0.0174643
R9106 VCC.n3705 VCC.n3428 0.0174643
R9107 VCC.n3581 VCC.n3485 0.0174643
R9108 VCC.n3580 VCC.n3491 0.0174643
R9109 VCC.n4132 VCC.n4036 0.0174643
R9110 VCC.n4131 VCC.n4042 0.0174643
R9111 VCC.n4255 VCC.n3978 0.0174643
R9112 VCC.n4256 VCC.n4255 0.0174643
R9113 VCC.n4260 VCC.n3980 0.0174643
R9114 VCC.n4257 VCC.n3980 0.0174643
R9115 VCC.n4380 VCC.n4379 0.0174643
R9116 VCC.n4379 VCC.n3911 0.0174643
R9117 VCC.n4381 VCC.n3916 0.0174643
R9118 VCC.n3916 VCC.n3912 0.0174643
R9119 VCC.n4942 VCC.n4473 0.0174643
R9120 VCC.n4942 VCC.n4941 0.0174643
R9121 VCC.n4934 VCC.n4474 0.0174643
R9122 VCC.n4940 VCC.n4474 0.0174643
R9123 VCC.n4812 VCC.n4535 0.0174643
R9124 VCC.n4813 VCC.n4812 0.0174643
R9125 VCC.n4817 VCC.n4537 0.0174643
R9126 VCC.n4814 VCC.n4537 0.0174643
R9127 VCC.n4690 VCC.n4594 0.0174643
R9128 VCC.n4689 VCC.n4600 0.0174643
R9129 VCC.n5241 VCC.n5145 0.0174643
R9130 VCC.n5240 VCC.n5151 0.0174643
R9131 VCC.n5364 VCC.n5087 0.0174643
R9132 VCC.n5365 VCC.n5364 0.0174643
R9133 VCC.n5369 VCC.n5089 0.0174643
R9134 VCC.n5366 VCC.n5089 0.0174643
R9135 VCC.n5489 VCC.n5488 0.0174643
R9136 VCC.n5488 VCC.n5020 0.0174643
R9137 VCC.n5490 VCC.n5025 0.0174643
R9138 VCC.n5025 VCC.n5021 0.0174643
R9139 VCC.n6050 VCC.n5581 0.0174643
R9140 VCC.n6050 VCC.n6049 0.0174643
R9141 VCC.n6042 VCC.n5582 0.0174643
R9142 VCC.n6048 VCC.n5582 0.0174643
R9143 VCC.n5920 VCC.n5643 0.0174643
R9144 VCC.n5921 VCC.n5920 0.0174643
R9145 VCC.n5925 VCC.n5645 0.0174643
R9146 VCC.n5922 VCC.n5645 0.0174643
R9147 VCC.n5798 VCC.n5702 0.0174643
R9148 VCC.n5797 VCC.n5708 0.0174643
R9149 VCC.n6348 VCC.n6252 0.0174643
R9150 VCC.n6347 VCC.n6258 0.0174643
R9151 VCC.n6471 VCC.n6194 0.0174643
R9152 VCC.n6472 VCC.n6471 0.0174643
R9153 VCC.n6476 VCC.n6196 0.0174643
R9154 VCC.n6473 VCC.n6196 0.0174643
R9155 VCC.n6596 VCC.n6595 0.0174643
R9156 VCC.n6595 VCC.n6127 0.0174643
R9157 VCC.n6597 VCC.n6132 0.0174643
R9158 VCC.n6132 VCC.n6128 0.0174643
R9159 VCC.n7157 VCC.n6688 0.0174643
R9160 VCC.n7157 VCC.n7156 0.0174643
R9161 VCC.n7149 VCC.n6689 0.0174643
R9162 VCC.n7155 VCC.n6689 0.0174643
R9163 VCC.n7027 VCC.n6750 0.0174643
R9164 VCC.n7028 VCC.n7027 0.0174643
R9165 VCC.n7032 VCC.n6752 0.0174643
R9166 VCC.n7029 VCC.n6752 0.0174643
R9167 VCC.n6905 VCC.n6809 0.0174643
R9168 VCC.n6904 VCC.n6815 0.0174643
R9169 VCC.n7455 VCC.n7359 0.0174643
R9170 VCC.n7454 VCC.n7365 0.0174643
R9171 VCC.n7578 VCC.n7301 0.0174643
R9172 VCC.n7579 VCC.n7578 0.0174643
R9173 VCC.n7583 VCC.n7303 0.0174643
R9174 VCC.n7580 VCC.n7303 0.0174643
R9175 VCC.n7703 VCC.n7702 0.0174643
R9176 VCC.n7702 VCC.n7234 0.0174643
R9177 VCC.n7704 VCC.n7239 0.0174643
R9178 VCC.n7239 VCC.n7235 0.0174643
R9179 VCC.n8264 VCC.n7795 0.0174643
R9180 VCC.n8264 VCC.n8263 0.0174643
R9181 VCC.n8256 VCC.n7796 0.0174643
R9182 VCC.n8262 VCC.n7796 0.0174643
R9183 VCC.n8134 VCC.n7857 0.0174643
R9184 VCC.n8135 VCC.n8134 0.0174643
R9185 VCC.n8139 VCC.n7859 0.0174643
R9186 VCC.n8136 VCC.n7859 0.0174643
R9187 VCC.n8012 VCC.n7916 0.0174643
R9188 VCC.n8011 VCC.n7922 0.0174643
R9189 VCC.n8498 VCC.n8408 0.0174643
R9190 VCC.n8499 VCC.n8498 0.0174643
R9191 VCC.n8503 VCC.n8410 0.0174643
R9192 VCC.n8500 VCC.n8410 0.0174643
R9193 VCC.n8623 VCC.n8622 0.0174643
R9194 VCC.n8622 VCC.n8341 0.0174643
R9195 VCC.n8624 VCC.n8346 0.0174643
R9196 VCC.n8346 VCC.n8342 0.0174643
R9197 VCC.n238 VCC.n233 0.0165714
R9198 VCC.n255 VCC.n254 0.0165714
R9199 VCC.n204 VCC.n197 0.0165714
R9200 VCC.n240 VCC.n239 0.0165714
R9201 VCC.n256 VCC.n167 0.0165714
R9202 VCC.n282 VCC.n146 0.0165714
R9203 VCC.n301 VCC.n300 0.0165714
R9204 VCC.n401 VCC.n400 0.0165714
R9205 VCC.n329 VCC.n321 0.0165714
R9206 VCC.n354 VCC.n348 0.0165714
R9207 VCC.n409 VCC.n86 0.0165714
R9208 VCC.n436 VCC.n435 0.0165714
R9209 VCC.n454 VCC.n60 0.0165714
R9210 VCC.n514 VCC.n29 0.0165714
R9211 VCC.n541 VCC.n10 0.0165714
R9212 VCC.n790 VCC.n785 0.0165714
R9213 VCC.n807 VCC.n806 0.0165714
R9214 VCC.n756 VCC.n749 0.0165714
R9215 VCC.n792 VCC.n791 0.0165714
R9216 VCC.n808 VCC.n719 0.0165714
R9217 VCC.n834 VCC.n698 0.0165714
R9218 VCC.n853 VCC.n852 0.0165714
R9219 VCC.n953 VCC.n952 0.0165714
R9220 VCC.n881 VCC.n873 0.0165714
R9221 VCC.n906 VCC.n900 0.0165714
R9222 VCC.n961 VCC.n638 0.0165714
R9223 VCC.n988 VCC.n987 0.0165714
R9224 VCC.n1006 VCC.n612 0.0165714
R9225 VCC.n1066 VCC.n581 0.0165714
R9226 VCC.n1095 VCC.n564 0.0165714
R9227 VCC.n1565 VCC.n1564 0.0165714
R9228 VCC.n1631 VCC.n1630 0.0165714
R9229 VCC.n1644 VCC.n1643 0.0165714
R9230 VCC.n1510 VCC.n1509 0.0165714
R9231 VCC.n1438 VCC.n1429 0.0165714
R9232 VCC.n1463 VCC.n1457 0.0165714
R9233 VCC.n1518 VCC.n1195 0.0165714
R9234 VCC.n1546 VCC.n1545 0.0165714
R9235 VCC.n1348 VCC.n1343 0.0165714
R9236 VCC.n1365 VCC.n1364 0.0165714
R9237 VCC.n1314 VCC.n1307 0.0165714
R9238 VCC.n1350 VCC.n1349 0.0165714
R9239 VCC.n1366 VCC.n1277 0.0165714
R9240 VCC.n1392 VCC.n1256 0.0165714
R9241 VCC.n1411 VCC.n1410 0.0165714
R9242 VCC.n1899 VCC.n1894 0.0165714
R9243 VCC.n1916 VCC.n1915 0.0165714
R9244 VCC.n1865 VCC.n1858 0.0165714
R9245 VCC.n1901 VCC.n1900 0.0165714
R9246 VCC.n1917 VCC.n1828 0.0165714
R9247 VCC.n1943 VCC.n1807 0.0165714
R9248 VCC.n1962 VCC.n1961 0.0165714
R9249 VCC.n2062 VCC.n2061 0.0165714
R9250 VCC.n1990 VCC.n1982 0.0165714
R9251 VCC.n2015 VCC.n2009 0.0165714
R9252 VCC.n2070 VCC.n1747 0.0165714
R9253 VCC.n2097 VCC.n2096 0.0165714
R9254 VCC.n2115 VCC.n1721 0.0165714
R9255 VCC.n2175 VCC.n1690 0.0165714
R9256 VCC.n2204 VCC.n1673 0.0165714
R9257 VCC.n2674 VCC.n2673 0.0165714
R9258 VCC.n2740 VCC.n2739 0.0165714
R9259 VCC.n2753 VCC.n2752 0.0165714
R9260 VCC.n2619 VCC.n2618 0.0165714
R9261 VCC.n2547 VCC.n2538 0.0165714
R9262 VCC.n2572 VCC.n2566 0.0165714
R9263 VCC.n2627 VCC.n2304 0.0165714
R9264 VCC.n2655 VCC.n2654 0.0165714
R9265 VCC.n2457 VCC.n2452 0.0165714
R9266 VCC.n2474 VCC.n2473 0.0165714
R9267 VCC.n2423 VCC.n2416 0.0165714
R9268 VCC.n2459 VCC.n2458 0.0165714
R9269 VCC.n2475 VCC.n2386 0.0165714
R9270 VCC.n2501 VCC.n2365 0.0165714
R9271 VCC.n2520 VCC.n2519 0.0165714
R9272 VCC.n3008 VCC.n3003 0.0165714
R9273 VCC.n3025 VCC.n3024 0.0165714
R9274 VCC.n2974 VCC.n2967 0.0165714
R9275 VCC.n3010 VCC.n3009 0.0165714
R9276 VCC.n3026 VCC.n2937 0.0165714
R9277 VCC.n3052 VCC.n2916 0.0165714
R9278 VCC.n3071 VCC.n3070 0.0165714
R9279 VCC.n3171 VCC.n3170 0.0165714
R9280 VCC.n3099 VCC.n3091 0.0165714
R9281 VCC.n3124 VCC.n3118 0.0165714
R9282 VCC.n3179 VCC.n2856 0.0165714
R9283 VCC.n3206 VCC.n3205 0.0165714
R9284 VCC.n3224 VCC.n2830 0.0165714
R9285 VCC.n3284 VCC.n2799 0.0165714
R9286 VCC.n3313 VCC.n2782 0.0165714
R9287 VCC.n3783 VCC.n3782 0.0165714
R9288 VCC.n3849 VCC.n3848 0.0165714
R9289 VCC.n3862 VCC.n3861 0.0165714
R9290 VCC.n3728 VCC.n3727 0.0165714
R9291 VCC.n3656 VCC.n3647 0.0165714
R9292 VCC.n3681 VCC.n3675 0.0165714
R9293 VCC.n3736 VCC.n3413 0.0165714
R9294 VCC.n3764 VCC.n3763 0.0165714
R9295 VCC.n3566 VCC.n3561 0.0165714
R9296 VCC.n3583 VCC.n3582 0.0165714
R9297 VCC.n3532 VCC.n3525 0.0165714
R9298 VCC.n3568 VCC.n3567 0.0165714
R9299 VCC.n3584 VCC.n3495 0.0165714
R9300 VCC.n3610 VCC.n3474 0.0165714
R9301 VCC.n3629 VCC.n3628 0.0165714
R9302 VCC.n4117 VCC.n4112 0.0165714
R9303 VCC.n4134 VCC.n4133 0.0165714
R9304 VCC.n4083 VCC.n4076 0.0165714
R9305 VCC.n4119 VCC.n4118 0.0165714
R9306 VCC.n4135 VCC.n4046 0.0165714
R9307 VCC.n4161 VCC.n4025 0.0165714
R9308 VCC.n4180 VCC.n4179 0.0165714
R9309 VCC.n4280 VCC.n4279 0.0165714
R9310 VCC.n4208 VCC.n4200 0.0165714
R9311 VCC.n4233 VCC.n4227 0.0165714
R9312 VCC.n4288 VCC.n3965 0.0165714
R9313 VCC.n4315 VCC.n4314 0.0165714
R9314 VCC.n4333 VCC.n3939 0.0165714
R9315 VCC.n4393 VCC.n3908 0.0165714
R9316 VCC.n4422 VCC.n3891 0.0165714
R9317 VCC.n4892 VCC.n4891 0.0165714
R9318 VCC.n4958 VCC.n4957 0.0165714
R9319 VCC.n4971 VCC.n4970 0.0165714
R9320 VCC.n4837 VCC.n4836 0.0165714
R9321 VCC.n4765 VCC.n4756 0.0165714
R9322 VCC.n4790 VCC.n4784 0.0165714
R9323 VCC.n4845 VCC.n4522 0.0165714
R9324 VCC.n4873 VCC.n4872 0.0165714
R9325 VCC.n4675 VCC.n4670 0.0165714
R9326 VCC.n4692 VCC.n4691 0.0165714
R9327 VCC.n4641 VCC.n4634 0.0165714
R9328 VCC.n4677 VCC.n4676 0.0165714
R9329 VCC.n4693 VCC.n4604 0.0165714
R9330 VCC.n4719 VCC.n4583 0.0165714
R9331 VCC.n4738 VCC.n4737 0.0165714
R9332 VCC.n5226 VCC.n5221 0.0165714
R9333 VCC.n5243 VCC.n5242 0.0165714
R9334 VCC.n5192 VCC.n5185 0.0165714
R9335 VCC.n5228 VCC.n5227 0.0165714
R9336 VCC.n5244 VCC.n5155 0.0165714
R9337 VCC.n5270 VCC.n5134 0.0165714
R9338 VCC.n5289 VCC.n5288 0.0165714
R9339 VCC.n5389 VCC.n5388 0.0165714
R9340 VCC.n5317 VCC.n5309 0.0165714
R9341 VCC.n5342 VCC.n5336 0.0165714
R9342 VCC.n5397 VCC.n5074 0.0165714
R9343 VCC.n5424 VCC.n5423 0.0165714
R9344 VCC.n5442 VCC.n5048 0.0165714
R9345 VCC.n5502 VCC.n5017 0.0165714
R9346 VCC.n5531 VCC.n5000 0.0165714
R9347 VCC.n6000 VCC.n5999 0.0165714
R9348 VCC.n6066 VCC.n6065 0.0165714
R9349 VCC.n6079 VCC.n6078 0.0165714
R9350 VCC.n5945 VCC.n5944 0.0165714
R9351 VCC.n5873 VCC.n5864 0.0165714
R9352 VCC.n5898 VCC.n5892 0.0165714
R9353 VCC.n5953 VCC.n5630 0.0165714
R9354 VCC.n5981 VCC.n5980 0.0165714
R9355 VCC.n5783 VCC.n5778 0.0165714
R9356 VCC.n5800 VCC.n5799 0.0165714
R9357 VCC.n5749 VCC.n5742 0.0165714
R9358 VCC.n5785 VCC.n5784 0.0165714
R9359 VCC.n5801 VCC.n5712 0.0165714
R9360 VCC.n5827 VCC.n5691 0.0165714
R9361 VCC.n5846 VCC.n5845 0.0165714
R9362 VCC.n6333 VCC.n6328 0.0165714
R9363 VCC.n6350 VCC.n6349 0.0165714
R9364 VCC.n6299 VCC.n6292 0.0165714
R9365 VCC.n6335 VCC.n6334 0.0165714
R9366 VCC.n6351 VCC.n6262 0.0165714
R9367 VCC.n6377 VCC.n6241 0.0165714
R9368 VCC.n6396 VCC.n6395 0.0165714
R9369 VCC.n6496 VCC.n6495 0.0165714
R9370 VCC.n6424 VCC.n6416 0.0165714
R9371 VCC.n6449 VCC.n6443 0.0165714
R9372 VCC.n6504 VCC.n6181 0.0165714
R9373 VCC.n6531 VCC.n6530 0.0165714
R9374 VCC.n6549 VCC.n6155 0.0165714
R9375 VCC.n6609 VCC.n6124 0.0165714
R9376 VCC.n6638 VCC.n6107 0.0165714
R9377 VCC.n7107 VCC.n7106 0.0165714
R9378 VCC.n7173 VCC.n7172 0.0165714
R9379 VCC.n7186 VCC.n7185 0.0165714
R9380 VCC.n7052 VCC.n7051 0.0165714
R9381 VCC.n6980 VCC.n6971 0.0165714
R9382 VCC.n7005 VCC.n6999 0.0165714
R9383 VCC.n7060 VCC.n6737 0.0165714
R9384 VCC.n7088 VCC.n7087 0.0165714
R9385 VCC.n6890 VCC.n6885 0.0165714
R9386 VCC.n6907 VCC.n6906 0.0165714
R9387 VCC.n6856 VCC.n6849 0.0165714
R9388 VCC.n6892 VCC.n6891 0.0165714
R9389 VCC.n6908 VCC.n6819 0.0165714
R9390 VCC.n6934 VCC.n6798 0.0165714
R9391 VCC.n6953 VCC.n6952 0.0165714
R9392 VCC.n7440 VCC.n7435 0.0165714
R9393 VCC.n7457 VCC.n7456 0.0165714
R9394 VCC.n7406 VCC.n7399 0.0165714
R9395 VCC.n7442 VCC.n7441 0.0165714
R9396 VCC.n7458 VCC.n7369 0.0165714
R9397 VCC.n7484 VCC.n7348 0.0165714
R9398 VCC.n7503 VCC.n7502 0.0165714
R9399 VCC.n7603 VCC.n7602 0.0165714
R9400 VCC.n7531 VCC.n7523 0.0165714
R9401 VCC.n7556 VCC.n7550 0.0165714
R9402 VCC.n7611 VCC.n7288 0.0165714
R9403 VCC.n7638 VCC.n7637 0.0165714
R9404 VCC.n7656 VCC.n7262 0.0165714
R9405 VCC.n7716 VCC.n7231 0.0165714
R9406 VCC.n7745 VCC.n7214 0.0165714
R9407 VCC.n8214 VCC.n8213 0.0165714
R9408 VCC.n8280 VCC.n8279 0.0165714
R9409 VCC.n8293 VCC.n8292 0.0165714
R9410 VCC.n8159 VCC.n8158 0.0165714
R9411 VCC.n8087 VCC.n8078 0.0165714
R9412 VCC.n8112 VCC.n8106 0.0165714
R9413 VCC.n8167 VCC.n7844 0.0165714
R9414 VCC.n8195 VCC.n8194 0.0165714
R9415 VCC.n7997 VCC.n7992 0.0165714
R9416 VCC.n8014 VCC.n8013 0.0165714
R9417 VCC.n7963 VCC.n7956 0.0165714
R9418 VCC.n7999 VCC.n7998 0.0165714
R9419 VCC.n8015 VCC.n7926 0.0165714
R9420 VCC.n8041 VCC.n7905 0.0165714
R9421 VCC.n8060 VCC.n8059 0.0165714
R9422 VCC.n8523 VCC.n8522 0.0165714
R9423 VCC.n8451 VCC.n8443 0.0165714
R9424 VCC.n8476 VCC.n8470 0.0165714
R9425 VCC.n8531 VCC.n8395 0.0165714
R9426 VCC.n8558 VCC.n8557 0.0165714
R9427 VCC.n8576 VCC.n8369 0.0165714
R9428 VCC.n8636 VCC.n8338 0.0165714
R9429 VCC.n8665 VCC.n8321 0.0165714
R9430 VCC.n274 VCC.n273 0.0156786
R9431 VCC.n240 VCC.n174 0.0156786
R9432 VCC.n356 VCC.n355 0.0156786
R9433 VCC.n410 VCC.n409 0.0156786
R9434 VCC.n480 VCC.n50 0.0156786
R9435 VCC.n826 VCC.n825 0.0156786
R9436 VCC.n792 VCC.n726 0.0156786
R9437 VCC.n908 VCC.n907 0.0156786
R9438 VCC.n962 VCC.n961 0.0156786
R9439 VCC.n1032 VCC.n602 0.0156786
R9440 VCC.n1598 VCC.n1155 0.0156786
R9441 VCC.n1465 VCC.n1464 0.0156786
R9442 VCC.n1519 VCC.n1518 0.0156786
R9443 VCC.n1384 VCC.n1383 0.0156786
R9444 VCC.n1350 VCC.n1284 0.0156786
R9445 VCC.n1935 VCC.n1934 0.0156786
R9446 VCC.n1901 VCC.n1835 0.0156786
R9447 VCC.n2017 VCC.n2016 0.0156786
R9448 VCC.n2071 VCC.n2070 0.0156786
R9449 VCC.n2141 VCC.n1711 0.0156786
R9450 VCC.n2707 VCC.n2264 0.0156786
R9451 VCC.n2574 VCC.n2573 0.0156786
R9452 VCC.n2628 VCC.n2627 0.0156786
R9453 VCC.n2493 VCC.n2492 0.0156786
R9454 VCC.n2459 VCC.n2393 0.0156786
R9455 VCC.n3044 VCC.n3043 0.0156786
R9456 VCC.n3010 VCC.n2944 0.0156786
R9457 VCC.n3126 VCC.n3125 0.0156786
R9458 VCC.n3180 VCC.n3179 0.0156786
R9459 VCC.n3250 VCC.n2820 0.0156786
R9460 VCC.n3816 VCC.n3373 0.0156786
R9461 VCC.n3683 VCC.n3682 0.0156786
R9462 VCC.n3737 VCC.n3736 0.0156786
R9463 VCC.n3602 VCC.n3601 0.0156786
R9464 VCC.n3568 VCC.n3502 0.0156786
R9465 VCC.n4153 VCC.n4152 0.0156786
R9466 VCC.n4119 VCC.n4053 0.0156786
R9467 VCC.n4235 VCC.n4234 0.0156786
R9468 VCC.n4289 VCC.n4288 0.0156786
R9469 VCC.n4359 VCC.n3929 0.0156786
R9470 VCC.n4925 VCC.n4482 0.0156786
R9471 VCC.n4792 VCC.n4791 0.0156786
R9472 VCC.n4846 VCC.n4845 0.0156786
R9473 VCC.n4711 VCC.n4710 0.0156786
R9474 VCC.n4677 VCC.n4611 0.0156786
R9475 VCC.n5262 VCC.n5261 0.0156786
R9476 VCC.n5228 VCC.n5162 0.0156786
R9477 VCC.n5344 VCC.n5343 0.0156786
R9478 VCC.n5398 VCC.n5397 0.0156786
R9479 VCC.n5468 VCC.n5038 0.0156786
R9480 VCC.n6033 VCC.n5590 0.0156786
R9481 VCC.n5900 VCC.n5899 0.0156786
R9482 VCC.n5954 VCC.n5953 0.0156786
R9483 VCC.n5819 VCC.n5818 0.0156786
R9484 VCC.n5785 VCC.n5719 0.0156786
R9485 VCC.n6369 VCC.n6368 0.0156786
R9486 VCC.n6335 VCC.n6269 0.0156786
R9487 VCC.n6451 VCC.n6450 0.0156786
R9488 VCC.n6505 VCC.n6504 0.0156786
R9489 VCC.n6575 VCC.n6145 0.0156786
R9490 VCC.n7140 VCC.n6697 0.0156786
R9491 VCC.n7007 VCC.n7006 0.0156786
R9492 VCC.n7061 VCC.n7060 0.0156786
R9493 VCC.n6926 VCC.n6925 0.0156786
R9494 VCC.n6892 VCC.n6826 0.0156786
R9495 VCC.n7476 VCC.n7475 0.0156786
R9496 VCC.n7442 VCC.n7376 0.0156786
R9497 VCC.n7558 VCC.n7557 0.0156786
R9498 VCC.n7612 VCC.n7611 0.0156786
R9499 VCC.n7682 VCC.n7252 0.0156786
R9500 VCC.n8247 VCC.n7804 0.0156786
R9501 VCC.n8114 VCC.n8113 0.0156786
R9502 VCC.n8168 VCC.n8167 0.0156786
R9503 VCC.n8033 VCC.n8032 0.0156786
R9504 VCC.n7999 VCC.n7933 0.0156786
R9505 VCC.n8478 VCC.n8477 0.0156786
R9506 VCC.n8532 VCC.n8531 0.0156786
R9507 VCC.n8602 VCC.n8359 0.0156786
R9508 VCC.n242 VCC.n241 0.0152714
R9509 VCC.n281 VCC.n280 0.0152714
R9510 VCC.n347 VCC.n102 0.0152714
R9511 VCC.n408 VCC.n407 0.0152714
R9512 VCC.n485 VCC.n481 0.0152714
R9513 VCC.n513 VCC.n512 0.0152714
R9514 VCC.n794 VCC.n793 0.0152714
R9515 VCC.n833 VCC.n832 0.0152714
R9516 VCC.n899 VCC.n654 0.0152714
R9517 VCC.n960 VCC.n959 0.0152714
R9518 VCC.n1037 VCC.n1033 0.0152714
R9519 VCC.n1065 VCC.n1064 0.0152714
R9520 VCC.n1352 VCC.n1351 0.0152714
R9521 VCC.n1391 VCC.n1390 0.0152714
R9522 VCC.n1456 VCC.n1211 0.0152714
R9523 VCC.n1517 VCC.n1516 0.0152714
R9524 VCC.n1600 VCC.n1599 0.0152714
R9525 VCC.n1629 VCC.n1628 0.0152714
R9526 VCC.n1903 VCC.n1902 0.0152714
R9527 VCC.n1942 VCC.n1941 0.0152714
R9528 VCC.n2008 VCC.n1763 0.0152714
R9529 VCC.n2069 VCC.n2068 0.0152714
R9530 VCC.n2146 VCC.n2142 0.0152714
R9531 VCC.n2174 VCC.n2173 0.0152714
R9532 VCC.n2461 VCC.n2460 0.0152714
R9533 VCC.n2500 VCC.n2499 0.0152714
R9534 VCC.n2565 VCC.n2320 0.0152714
R9535 VCC.n2626 VCC.n2625 0.0152714
R9536 VCC.n2709 VCC.n2708 0.0152714
R9537 VCC.n2738 VCC.n2737 0.0152714
R9538 VCC.n3012 VCC.n3011 0.0152714
R9539 VCC.n3051 VCC.n3050 0.0152714
R9540 VCC.n3117 VCC.n2872 0.0152714
R9541 VCC.n3178 VCC.n3177 0.0152714
R9542 VCC.n3255 VCC.n3251 0.0152714
R9543 VCC.n3283 VCC.n3282 0.0152714
R9544 VCC.n3570 VCC.n3569 0.0152714
R9545 VCC.n3609 VCC.n3608 0.0152714
R9546 VCC.n3674 VCC.n3429 0.0152714
R9547 VCC.n3735 VCC.n3734 0.0152714
R9548 VCC.n3818 VCC.n3817 0.0152714
R9549 VCC.n3847 VCC.n3846 0.0152714
R9550 VCC.n4121 VCC.n4120 0.0152714
R9551 VCC.n4160 VCC.n4159 0.0152714
R9552 VCC.n4226 VCC.n3981 0.0152714
R9553 VCC.n4287 VCC.n4286 0.0152714
R9554 VCC.n4364 VCC.n4360 0.0152714
R9555 VCC.n4392 VCC.n4391 0.0152714
R9556 VCC.n4679 VCC.n4678 0.0152714
R9557 VCC.n4718 VCC.n4717 0.0152714
R9558 VCC.n4783 VCC.n4538 0.0152714
R9559 VCC.n4844 VCC.n4843 0.0152714
R9560 VCC.n4927 VCC.n4926 0.0152714
R9561 VCC.n4956 VCC.n4955 0.0152714
R9562 VCC.n5230 VCC.n5229 0.0152714
R9563 VCC.n5269 VCC.n5268 0.0152714
R9564 VCC.n5335 VCC.n5090 0.0152714
R9565 VCC.n5396 VCC.n5395 0.0152714
R9566 VCC.n5473 VCC.n5469 0.0152714
R9567 VCC.n5501 VCC.n5500 0.0152714
R9568 VCC.n5787 VCC.n5786 0.0152714
R9569 VCC.n5826 VCC.n5825 0.0152714
R9570 VCC.n5891 VCC.n5646 0.0152714
R9571 VCC.n5952 VCC.n5951 0.0152714
R9572 VCC.n6035 VCC.n6034 0.0152714
R9573 VCC.n6064 VCC.n6063 0.0152714
R9574 VCC.n6337 VCC.n6336 0.0152714
R9575 VCC.n6376 VCC.n6375 0.0152714
R9576 VCC.n6442 VCC.n6197 0.0152714
R9577 VCC.n6503 VCC.n6502 0.0152714
R9578 VCC.n6580 VCC.n6576 0.0152714
R9579 VCC.n6608 VCC.n6607 0.0152714
R9580 VCC.n6894 VCC.n6893 0.0152714
R9581 VCC.n6933 VCC.n6932 0.0152714
R9582 VCC.n6998 VCC.n6753 0.0152714
R9583 VCC.n7059 VCC.n7058 0.0152714
R9584 VCC.n7142 VCC.n7141 0.0152714
R9585 VCC.n7171 VCC.n7170 0.0152714
R9586 VCC.n7444 VCC.n7443 0.0152714
R9587 VCC.n7483 VCC.n7482 0.0152714
R9588 VCC.n7549 VCC.n7304 0.0152714
R9589 VCC.n7610 VCC.n7609 0.0152714
R9590 VCC.n7687 VCC.n7683 0.0152714
R9591 VCC.n7715 VCC.n7714 0.0152714
R9592 VCC.n8001 VCC.n8000 0.0152714
R9593 VCC.n8040 VCC.n8039 0.0152714
R9594 VCC.n8105 VCC.n7860 0.0152714
R9595 VCC.n8166 VCC.n8165 0.0152714
R9596 VCC.n8249 VCC.n8248 0.0152714
R9597 VCC.n8278 VCC.n8277 0.0152714
R9598 VCC.n8469 VCC.n8411 0.0152714
R9599 VCC.n8530 VCC.n8529 0.0152714
R9600 VCC.n8607 VCC.n8603 0.0152714
R9601 VCC.n8635 VCC.n8634 0.0152714
R9602 VCC.n283 VCC.n282 0.0147857
R9603 VCC.n348 VCC.n113 0.0147857
R9604 VCC.n462 VCC.n52 0.0147857
R9605 VCC.n835 VCC.n834 0.0147857
R9606 VCC.n900 VCC.n665 0.0147857
R9607 VCC.n1014 VCC.n604 0.0147857
R9608 VCC.n1168 VCC.n1157 0.0147857
R9609 VCC.n1457 VCC.n1222 0.0147857
R9610 VCC.n1393 VCC.n1392 0.0147857
R9611 VCC.n1944 VCC.n1943 0.0147857
R9612 VCC.n2009 VCC.n1774 0.0147857
R9613 VCC.n2123 VCC.n1713 0.0147857
R9614 VCC.n2277 VCC.n2266 0.0147857
R9615 VCC.n2566 VCC.n2331 0.0147857
R9616 VCC.n2502 VCC.n2501 0.0147857
R9617 VCC.n3053 VCC.n3052 0.0147857
R9618 VCC.n3118 VCC.n2883 0.0147857
R9619 VCC.n3232 VCC.n2822 0.0147857
R9620 VCC.n3386 VCC.n3375 0.0147857
R9621 VCC.n3675 VCC.n3440 0.0147857
R9622 VCC.n3611 VCC.n3610 0.0147857
R9623 VCC.n4162 VCC.n4161 0.0147857
R9624 VCC.n4227 VCC.n3992 0.0147857
R9625 VCC.n4341 VCC.n3931 0.0147857
R9626 VCC.n4495 VCC.n4484 0.0147857
R9627 VCC.n4784 VCC.n4549 0.0147857
R9628 VCC.n4720 VCC.n4719 0.0147857
R9629 VCC.n5271 VCC.n5270 0.0147857
R9630 VCC.n5336 VCC.n5101 0.0147857
R9631 VCC.n5450 VCC.n5040 0.0147857
R9632 VCC.n5603 VCC.n5592 0.0147857
R9633 VCC.n5892 VCC.n5657 0.0147857
R9634 VCC.n5828 VCC.n5827 0.0147857
R9635 VCC.n6378 VCC.n6377 0.0147857
R9636 VCC.n6443 VCC.n6208 0.0147857
R9637 VCC.n6557 VCC.n6147 0.0147857
R9638 VCC.n6710 VCC.n6699 0.0147857
R9639 VCC.n6999 VCC.n6764 0.0147857
R9640 VCC.n6935 VCC.n6934 0.0147857
R9641 VCC.n7485 VCC.n7484 0.0147857
R9642 VCC.n7550 VCC.n7315 0.0147857
R9643 VCC.n7664 VCC.n7254 0.0147857
R9644 VCC.n7817 VCC.n7806 0.0147857
R9645 VCC.n8106 VCC.n7871 0.0147857
R9646 VCC.n8042 VCC.n8041 0.0147857
R9647 VCC.n8470 VCC.n8422 0.0147857
R9648 VCC.n8584 VCC.n8361 0.0147857
R9649 VCC.n258 VCC.n257 0.0132571
R9650 VCC.n380 VCC.n379 0.0132571
R9651 VCC.n504 VCC.n503 0.0132571
R9652 VCC.n810 VCC.n809 0.0132571
R9653 VCC.n932 VCC.n931 0.0132571
R9654 VCC.n1056 VCC.n1055 0.0132571
R9655 VCC.n1368 VCC.n1367 0.0132571
R9656 VCC.n1489 VCC.n1488 0.0132571
R9657 VCC.n1612 VCC.n1608 0.0132571
R9658 VCC.n1919 VCC.n1918 0.0132571
R9659 VCC.n2041 VCC.n2040 0.0132571
R9660 VCC.n2165 VCC.n2164 0.0132571
R9661 VCC.n2477 VCC.n2476 0.0132571
R9662 VCC.n2598 VCC.n2597 0.0132571
R9663 VCC.n2721 VCC.n2717 0.0132571
R9664 VCC.n3028 VCC.n3027 0.0132571
R9665 VCC.n3150 VCC.n3149 0.0132571
R9666 VCC.n3274 VCC.n3273 0.0132571
R9667 VCC.n3586 VCC.n3585 0.0132571
R9668 VCC.n3707 VCC.n3706 0.0132571
R9669 VCC.n3830 VCC.n3826 0.0132571
R9670 VCC.n4137 VCC.n4136 0.0132571
R9671 VCC.n4259 VCC.n4258 0.0132571
R9672 VCC.n4383 VCC.n4382 0.0132571
R9673 VCC.n4695 VCC.n4694 0.0132571
R9674 VCC.n4816 VCC.n4815 0.0132571
R9675 VCC.n4939 VCC.n4935 0.0132571
R9676 VCC.n5246 VCC.n5245 0.0132571
R9677 VCC.n5368 VCC.n5367 0.0132571
R9678 VCC.n5492 VCC.n5491 0.0132571
R9679 VCC.n5803 VCC.n5802 0.0132571
R9680 VCC.n5924 VCC.n5923 0.0132571
R9681 VCC.n6047 VCC.n6043 0.0132571
R9682 VCC.n6353 VCC.n6352 0.0132571
R9683 VCC.n6475 VCC.n6474 0.0132571
R9684 VCC.n6599 VCC.n6598 0.0132571
R9685 VCC.n6910 VCC.n6909 0.0132571
R9686 VCC.n7031 VCC.n7030 0.0132571
R9687 VCC.n7154 VCC.n7150 0.0132571
R9688 VCC.n7460 VCC.n7459 0.0132571
R9689 VCC.n7582 VCC.n7581 0.0132571
R9690 VCC.n7706 VCC.n7705 0.0132571
R9691 VCC.n8017 VCC.n8016 0.0132571
R9692 VCC.n8138 VCC.n8137 0.0132571
R9693 VCC.n8261 VCC.n8257 0.0132571
R9694 VCC.n8502 VCC.n8501 0.0132571
R9695 VCC.n8626 VCC.n8625 0.0132571
R9696 VCC.n202 VCC.n200 0.013
R9697 VCC.n76 VCC.n74 0.013
R9698 VCC.n542 VCC.n9 0.013
R9699 VCC.n550 VCC.n2 0.013
R9700 VCC.n541 VCC.n540 0.013
R9701 VCC.n754 VCC.n752 0.013
R9702 VCC.n628 VCC.n626 0.013
R9703 VCC.n1096 VCC.n563 0.013
R9704 VCC.n1104 VCC.n556 0.013
R9705 VCC.n1095 VCC.n1094 0.013
R9706 VCC.n1642 VCC.n1641 0.013
R9707 VCC.n1658 VCC.n1110 0.013
R9708 VCC.n1643 VCC.n1121 0.013
R9709 VCC.n1185 VCC.n1183 0.013
R9710 VCC.n1312 VCC.n1310 0.013
R9711 VCC.n1863 VCC.n1861 0.013
R9712 VCC.n1737 VCC.n1735 0.013
R9713 VCC.n2205 VCC.n1672 0.013
R9714 VCC.n2213 VCC.n1665 0.013
R9715 VCC.n2204 VCC.n2203 0.013
R9716 VCC.n2751 VCC.n2750 0.013
R9717 VCC.n2767 VCC.n2219 0.013
R9718 VCC.n2752 VCC.n2230 0.013
R9719 VCC.n2294 VCC.n2292 0.013
R9720 VCC.n2421 VCC.n2419 0.013
R9721 VCC.n2972 VCC.n2970 0.013
R9722 VCC.n2846 VCC.n2844 0.013
R9723 VCC.n3314 VCC.n2781 0.013
R9724 VCC.n3322 VCC.n2774 0.013
R9725 VCC.n3313 VCC.n3312 0.013
R9726 VCC.n3860 VCC.n3859 0.013
R9727 VCC.n3876 VCC.n3328 0.013
R9728 VCC.n3861 VCC.n3339 0.013
R9729 VCC.n3403 VCC.n3401 0.013
R9730 VCC.n3530 VCC.n3528 0.013
R9731 VCC.n4081 VCC.n4079 0.013
R9732 VCC.n3955 VCC.n3953 0.013
R9733 VCC.n4423 VCC.n3890 0.013
R9734 VCC.n4431 VCC.n3883 0.013
R9735 VCC.n4422 VCC.n4421 0.013
R9736 VCC.n4969 VCC.n4968 0.013
R9737 VCC.n4985 VCC.n4437 0.013
R9738 VCC.n4970 VCC.n4448 0.013
R9739 VCC.n4512 VCC.n4510 0.013
R9740 VCC.n4639 VCC.n4637 0.013
R9741 VCC.n5190 VCC.n5188 0.013
R9742 VCC.n5064 VCC.n5062 0.013
R9743 VCC.n5532 VCC.n4999 0.013
R9744 VCC.n5540 VCC.n4992 0.013
R9745 VCC.n5531 VCC.n5530 0.013
R9746 VCC.n6077 VCC.n6076 0.013
R9747 VCC.n6093 VCC.n5545 0.013
R9748 VCC.n6078 VCC.n5556 0.013
R9749 VCC.n5620 VCC.n5618 0.013
R9750 VCC.n5747 VCC.n5745 0.013
R9751 VCC.n6297 VCC.n6295 0.013
R9752 VCC.n6171 VCC.n6169 0.013
R9753 VCC.n6639 VCC.n6106 0.013
R9754 VCC.n6647 VCC.n6099 0.013
R9755 VCC.n6638 VCC.n6637 0.013
R9756 VCC.n7184 VCC.n7183 0.013
R9757 VCC.n7200 VCC.n6652 0.013
R9758 VCC.n7185 VCC.n6663 0.013
R9759 VCC.n6727 VCC.n6725 0.013
R9760 VCC.n6854 VCC.n6852 0.013
R9761 VCC.n7404 VCC.n7402 0.013
R9762 VCC.n7278 VCC.n7276 0.013
R9763 VCC.n7746 VCC.n7213 0.013
R9764 VCC.n7754 VCC.n7206 0.013
R9765 VCC.n7745 VCC.n7744 0.013
R9766 VCC.n8291 VCC.n8290 0.013
R9767 VCC.n8307 VCC.n7759 0.013
R9768 VCC.n8292 VCC.n7770 0.013
R9769 VCC.n7834 VCC.n7832 0.013
R9770 VCC.n7961 VCC.n7959 0.013
R9771 VCC.n8385 VCC.n8383 0.013
R9772 VCC.n8666 VCC.n8320 0.013
R9773 VCC.n8674 VCC.n8313 0.013
R9774 VCC.n8665 VCC.n8664 0.013
R9775 VCC.n137 VCC.n135 0.0121071
R9776 VCC.n205 VCC.n204 0.0121071
R9777 VCC.n327 VCC.n324 0.0121071
R9778 VCC.n446 VCC.n445 0.0121071
R9779 VCC.n435 VCC.n75 0.0121071
R9780 VCC.n458 VCC.n451 0.0121071
R9781 VCC.n456 VCC.n453 0.0121071
R9782 VCC.n455 VCC.n454 0.0121071
R9783 VCC.n18 VCC.n15 0.0121071
R9784 VCC.n689 VCC.n687 0.0121071
R9785 VCC.n757 VCC.n756 0.0121071
R9786 VCC.n879 VCC.n876 0.0121071
R9787 VCC.n998 VCC.n997 0.0121071
R9788 VCC.n987 VCC.n627 0.0121071
R9789 VCC.n1010 VCC.n1003 0.0121071
R9790 VCC.n1008 VCC.n1005 0.0121071
R9791 VCC.n1007 VCC.n1006 0.0121071
R9792 VCC.n570 VCC.n567 0.0121071
R9793 VCC.n1569 VCC.n1561 0.0121071
R9794 VCC.n1567 VCC.n1563 0.0121071
R9795 VCC.n1566 VCC.n1565 0.0121071
R9796 VCC.n1645 VCC.n1120 0.0121071
R9797 VCC.n1436 VCC.n1433 0.0121071
R9798 VCC.n1556 VCC.n1555 0.0121071
R9799 VCC.n1545 VCC.n1184 0.0121071
R9800 VCC.n1247 VCC.n1245 0.0121071
R9801 VCC.n1315 VCC.n1314 0.0121071
R9802 VCC.n1798 VCC.n1796 0.0121071
R9803 VCC.n1866 VCC.n1865 0.0121071
R9804 VCC.n1988 VCC.n1985 0.0121071
R9805 VCC.n2107 VCC.n2106 0.0121071
R9806 VCC.n2096 VCC.n1736 0.0121071
R9807 VCC.n2119 VCC.n2112 0.0121071
R9808 VCC.n2117 VCC.n2114 0.0121071
R9809 VCC.n2116 VCC.n2115 0.0121071
R9810 VCC.n1679 VCC.n1676 0.0121071
R9811 VCC.n2678 VCC.n2670 0.0121071
R9812 VCC.n2676 VCC.n2672 0.0121071
R9813 VCC.n2675 VCC.n2674 0.0121071
R9814 VCC.n2754 VCC.n2229 0.0121071
R9815 VCC.n2545 VCC.n2542 0.0121071
R9816 VCC.n2665 VCC.n2664 0.0121071
R9817 VCC.n2654 VCC.n2293 0.0121071
R9818 VCC.n2356 VCC.n2354 0.0121071
R9819 VCC.n2424 VCC.n2423 0.0121071
R9820 VCC.n2907 VCC.n2905 0.0121071
R9821 VCC.n2975 VCC.n2974 0.0121071
R9822 VCC.n3097 VCC.n3094 0.0121071
R9823 VCC.n3216 VCC.n3215 0.0121071
R9824 VCC.n3205 VCC.n2845 0.0121071
R9825 VCC.n3228 VCC.n3221 0.0121071
R9826 VCC.n3226 VCC.n3223 0.0121071
R9827 VCC.n3225 VCC.n3224 0.0121071
R9828 VCC.n2788 VCC.n2785 0.0121071
R9829 VCC.n3787 VCC.n3779 0.0121071
R9830 VCC.n3785 VCC.n3781 0.0121071
R9831 VCC.n3784 VCC.n3783 0.0121071
R9832 VCC.n3863 VCC.n3338 0.0121071
R9833 VCC.n3654 VCC.n3651 0.0121071
R9834 VCC.n3774 VCC.n3773 0.0121071
R9835 VCC.n3763 VCC.n3402 0.0121071
R9836 VCC.n3465 VCC.n3463 0.0121071
R9837 VCC.n3533 VCC.n3532 0.0121071
R9838 VCC.n4016 VCC.n4014 0.0121071
R9839 VCC.n4084 VCC.n4083 0.0121071
R9840 VCC.n4206 VCC.n4203 0.0121071
R9841 VCC.n4325 VCC.n4324 0.0121071
R9842 VCC.n4314 VCC.n3954 0.0121071
R9843 VCC.n4337 VCC.n4330 0.0121071
R9844 VCC.n4335 VCC.n4332 0.0121071
R9845 VCC.n4334 VCC.n4333 0.0121071
R9846 VCC.n3897 VCC.n3894 0.0121071
R9847 VCC.n4896 VCC.n4888 0.0121071
R9848 VCC.n4894 VCC.n4890 0.0121071
R9849 VCC.n4893 VCC.n4892 0.0121071
R9850 VCC.n4972 VCC.n4447 0.0121071
R9851 VCC.n4763 VCC.n4760 0.0121071
R9852 VCC.n4883 VCC.n4882 0.0121071
R9853 VCC.n4872 VCC.n4511 0.0121071
R9854 VCC.n4574 VCC.n4572 0.0121071
R9855 VCC.n4642 VCC.n4641 0.0121071
R9856 VCC.n5125 VCC.n5123 0.0121071
R9857 VCC.n5193 VCC.n5192 0.0121071
R9858 VCC.n5315 VCC.n5312 0.0121071
R9859 VCC.n5434 VCC.n5433 0.0121071
R9860 VCC.n5423 VCC.n5063 0.0121071
R9861 VCC.n5446 VCC.n5439 0.0121071
R9862 VCC.n5444 VCC.n5441 0.0121071
R9863 VCC.n5443 VCC.n5442 0.0121071
R9864 VCC.n5006 VCC.n5003 0.0121071
R9865 VCC.n6004 VCC.n5996 0.0121071
R9866 VCC.n6002 VCC.n5998 0.0121071
R9867 VCC.n6001 VCC.n6000 0.0121071
R9868 VCC.n6080 VCC.n5555 0.0121071
R9869 VCC.n5871 VCC.n5868 0.0121071
R9870 VCC.n5991 VCC.n5990 0.0121071
R9871 VCC.n5980 VCC.n5619 0.0121071
R9872 VCC.n5682 VCC.n5680 0.0121071
R9873 VCC.n5750 VCC.n5749 0.0121071
R9874 VCC.n6232 VCC.n6230 0.0121071
R9875 VCC.n6300 VCC.n6299 0.0121071
R9876 VCC.n6422 VCC.n6419 0.0121071
R9877 VCC.n6541 VCC.n6540 0.0121071
R9878 VCC.n6530 VCC.n6170 0.0121071
R9879 VCC.n6553 VCC.n6546 0.0121071
R9880 VCC.n6551 VCC.n6548 0.0121071
R9881 VCC.n6550 VCC.n6549 0.0121071
R9882 VCC.n6113 VCC.n6110 0.0121071
R9883 VCC.n7111 VCC.n7103 0.0121071
R9884 VCC.n7109 VCC.n7105 0.0121071
R9885 VCC.n7108 VCC.n7107 0.0121071
R9886 VCC.n7187 VCC.n6662 0.0121071
R9887 VCC.n6978 VCC.n6975 0.0121071
R9888 VCC.n7098 VCC.n7097 0.0121071
R9889 VCC.n7087 VCC.n6726 0.0121071
R9890 VCC.n6789 VCC.n6787 0.0121071
R9891 VCC.n6857 VCC.n6856 0.0121071
R9892 VCC.n7339 VCC.n7337 0.0121071
R9893 VCC.n7407 VCC.n7406 0.0121071
R9894 VCC.n7529 VCC.n7526 0.0121071
R9895 VCC.n7648 VCC.n7647 0.0121071
R9896 VCC.n7637 VCC.n7277 0.0121071
R9897 VCC.n7660 VCC.n7653 0.0121071
R9898 VCC.n7658 VCC.n7655 0.0121071
R9899 VCC.n7657 VCC.n7656 0.0121071
R9900 VCC.n7220 VCC.n7217 0.0121071
R9901 VCC.n8218 VCC.n8210 0.0121071
R9902 VCC.n8216 VCC.n8212 0.0121071
R9903 VCC.n8215 VCC.n8214 0.0121071
R9904 VCC.n8294 VCC.n7769 0.0121071
R9905 VCC.n8085 VCC.n8082 0.0121071
R9906 VCC.n8205 VCC.n8204 0.0121071
R9907 VCC.n8194 VCC.n7833 0.0121071
R9908 VCC.n7896 VCC.n7894 0.0121071
R9909 VCC.n7964 VCC.n7963 0.0121071
R9910 VCC.n8449 VCC.n8446 0.0121071
R9911 VCC.n8568 VCC.n8567 0.0121071
R9912 VCC.n8557 VCC.n8384 0.0121071
R9913 VCC.n8580 VCC.n8573 0.0121071
R9914 VCC.n8578 VCC.n8575 0.0121071
R9915 VCC.n8577 VCC.n8576 0.0121071
R9916 VCC.n8327 VCC.n8324 0.0121071
R9917 VCC.n199 VCC.n185 0.0112143
R9918 VCC.n303 VCC.n135 0.0112143
R9919 VCC.n311 VCC.n310 0.0112143
R9920 VCC.n198 VCC.n186 0.0112143
R9921 VCC.n302 VCC.n301 0.0112143
R9922 VCC.n300 VCC.n136 0.0112143
R9923 VCC.n324 VCC.n323 0.0112143
R9924 VCC.n439 VCC.n438 0.0112143
R9925 VCC.n330 VCC.n329 0.0112143
R9926 VCC.n322 VCC.n321 0.0112143
R9927 VCC.n437 VCC.n72 0.0112143
R9928 VCC.n453 VCC.n452 0.0112143
R9929 VCC.n467 VCC.n59 0.0112143
R9930 VCC.n533 VCC.n532 0.0112143
R9931 VCC.n466 VCC.n465 0.0112143
R9932 VCC.n751 VCC.n737 0.0112143
R9933 VCC.n855 VCC.n687 0.0112143
R9934 VCC.n863 VCC.n862 0.0112143
R9935 VCC.n750 VCC.n738 0.0112143
R9936 VCC.n854 VCC.n853 0.0112143
R9937 VCC.n852 VCC.n688 0.0112143
R9938 VCC.n876 VCC.n875 0.0112143
R9939 VCC.n991 VCC.n990 0.0112143
R9940 VCC.n882 VCC.n881 0.0112143
R9941 VCC.n874 VCC.n873 0.0112143
R9942 VCC.n989 VCC.n624 0.0112143
R9943 VCC.n1005 VCC.n1004 0.0112143
R9944 VCC.n1019 VCC.n611 0.0112143
R9945 VCC.n1085 VCC.n1084 0.0112143
R9946 VCC.n1018 VCC.n1017 0.0112143
R9947 VCC.n1563 VCC.n1562 0.0112143
R9948 VCC.n1576 VCC.n1575 0.0112143
R9949 VCC.n1647 VCC.n1118 0.0112143
R9950 VCC.n1574 VCC.n1167 0.0112143
R9951 VCC.n1433 VCC.n1432 0.0112143
R9952 VCC.n1549 VCC.n1548 0.0112143
R9953 VCC.n1439 VCC.n1438 0.0112143
R9954 VCC.n1431 VCC.n1429 0.0112143
R9955 VCC.n1547 VCC.n1181 0.0112143
R9956 VCC.n1309 VCC.n1295 0.0112143
R9957 VCC.n1413 VCC.n1245 0.0112143
R9958 VCC.n1421 VCC.n1420 0.0112143
R9959 VCC.n1308 VCC.n1296 0.0112143
R9960 VCC.n1412 VCC.n1411 0.0112143
R9961 VCC.n1410 VCC.n1246 0.0112143
R9962 VCC.n1860 VCC.n1846 0.0112143
R9963 VCC.n1964 VCC.n1796 0.0112143
R9964 VCC.n1972 VCC.n1971 0.0112143
R9965 VCC.n1859 VCC.n1847 0.0112143
R9966 VCC.n1963 VCC.n1962 0.0112143
R9967 VCC.n1961 VCC.n1797 0.0112143
R9968 VCC.n1985 VCC.n1984 0.0112143
R9969 VCC.n2100 VCC.n2099 0.0112143
R9970 VCC.n1991 VCC.n1990 0.0112143
R9971 VCC.n1983 VCC.n1982 0.0112143
R9972 VCC.n2098 VCC.n1733 0.0112143
R9973 VCC.n2114 VCC.n2113 0.0112143
R9974 VCC.n2128 VCC.n1720 0.0112143
R9975 VCC.n2194 VCC.n2193 0.0112143
R9976 VCC.n2127 VCC.n2126 0.0112143
R9977 VCC.n2672 VCC.n2671 0.0112143
R9978 VCC.n2685 VCC.n2684 0.0112143
R9979 VCC.n2756 VCC.n2227 0.0112143
R9980 VCC.n2683 VCC.n2276 0.0112143
R9981 VCC.n2542 VCC.n2541 0.0112143
R9982 VCC.n2658 VCC.n2657 0.0112143
R9983 VCC.n2548 VCC.n2547 0.0112143
R9984 VCC.n2540 VCC.n2538 0.0112143
R9985 VCC.n2656 VCC.n2290 0.0112143
R9986 VCC.n2418 VCC.n2404 0.0112143
R9987 VCC.n2522 VCC.n2354 0.0112143
R9988 VCC.n2530 VCC.n2529 0.0112143
R9989 VCC.n2417 VCC.n2405 0.0112143
R9990 VCC.n2521 VCC.n2520 0.0112143
R9991 VCC.n2519 VCC.n2355 0.0112143
R9992 VCC.n2969 VCC.n2955 0.0112143
R9993 VCC.n3073 VCC.n2905 0.0112143
R9994 VCC.n3081 VCC.n3080 0.0112143
R9995 VCC.n2968 VCC.n2956 0.0112143
R9996 VCC.n3072 VCC.n3071 0.0112143
R9997 VCC.n3070 VCC.n2906 0.0112143
R9998 VCC.n3094 VCC.n3093 0.0112143
R9999 VCC.n3209 VCC.n3208 0.0112143
R10000 VCC.n3100 VCC.n3099 0.0112143
R10001 VCC.n3092 VCC.n3091 0.0112143
R10002 VCC.n3207 VCC.n2842 0.0112143
R10003 VCC.n3223 VCC.n3222 0.0112143
R10004 VCC.n3237 VCC.n2829 0.0112143
R10005 VCC.n3303 VCC.n3302 0.0112143
R10006 VCC.n3236 VCC.n3235 0.0112143
R10007 VCC.n3781 VCC.n3780 0.0112143
R10008 VCC.n3794 VCC.n3793 0.0112143
R10009 VCC.n3865 VCC.n3336 0.0112143
R10010 VCC.n3792 VCC.n3385 0.0112143
R10011 VCC.n3651 VCC.n3650 0.0112143
R10012 VCC.n3767 VCC.n3766 0.0112143
R10013 VCC.n3657 VCC.n3656 0.0112143
R10014 VCC.n3649 VCC.n3647 0.0112143
R10015 VCC.n3765 VCC.n3399 0.0112143
R10016 VCC.n3527 VCC.n3513 0.0112143
R10017 VCC.n3631 VCC.n3463 0.0112143
R10018 VCC.n3639 VCC.n3638 0.0112143
R10019 VCC.n3526 VCC.n3514 0.0112143
R10020 VCC.n3630 VCC.n3629 0.0112143
R10021 VCC.n3628 VCC.n3464 0.0112143
R10022 VCC.n4078 VCC.n4064 0.0112143
R10023 VCC.n4182 VCC.n4014 0.0112143
R10024 VCC.n4190 VCC.n4189 0.0112143
R10025 VCC.n4077 VCC.n4065 0.0112143
R10026 VCC.n4181 VCC.n4180 0.0112143
R10027 VCC.n4179 VCC.n4015 0.0112143
R10028 VCC.n4203 VCC.n4202 0.0112143
R10029 VCC.n4318 VCC.n4317 0.0112143
R10030 VCC.n4209 VCC.n4208 0.0112143
R10031 VCC.n4201 VCC.n4200 0.0112143
R10032 VCC.n4316 VCC.n3951 0.0112143
R10033 VCC.n4332 VCC.n4331 0.0112143
R10034 VCC.n4346 VCC.n3938 0.0112143
R10035 VCC.n4412 VCC.n4411 0.0112143
R10036 VCC.n4345 VCC.n4344 0.0112143
R10037 VCC.n4890 VCC.n4889 0.0112143
R10038 VCC.n4903 VCC.n4902 0.0112143
R10039 VCC.n4974 VCC.n4445 0.0112143
R10040 VCC.n4901 VCC.n4494 0.0112143
R10041 VCC.n4760 VCC.n4759 0.0112143
R10042 VCC.n4876 VCC.n4875 0.0112143
R10043 VCC.n4766 VCC.n4765 0.0112143
R10044 VCC.n4758 VCC.n4756 0.0112143
R10045 VCC.n4874 VCC.n4508 0.0112143
R10046 VCC.n4636 VCC.n4622 0.0112143
R10047 VCC.n4740 VCC.n4572 0.0112143
R10048 VCC.n4748 VCC.n4747 0.0112143
R10049 VCC.n4635 VCC.n4623 0.0112143
R10050 VCC.n4739 VCC.n4738 0.0112143
R10051 VCC.n4737 VCC.n4573 0.0112143
R10052 VCC.n5187 VCC.n5173 0.0112143
R10053 VCC.n5291 VCC.n5123 0.0112143
R10054 VCC.n5299 VCC.n5298 0.0112143
R10055 VCC.n5186 VCC.n5174 0.0112143
R10056 VCC.n5290 VCC.n5289 0.0112143
R10057 VCC.n5288 VCC.n5124 0.0112143
R10058 VCC.n5312 VCC.n5311 0.0112143
R10059 VCC.n5427 VCC.n5426 0.0112143
R10060 VCC.n5318 VCC.n5317 0.0112143
R10061 VCC.n5310 VCC.n5309 0.0112143
R10062 VCC.n5425 VCC.n5060 0.0112143
R10063 VCC.n5441 VCC.n5440 0.0112143
R10064 VCC.n5455 VCC.n5047 0.0112143
R10065 VCC.n5521 VCC.n5520 0.0112143
R10066 VCC.n5454 VCC.n5453 0.0112143
R10067 VCC.n5998 VCC.n5997 0.0112143
R10068 VCC.n6011 VCC.n6010 0.0112143
R10069 VCC.n6082 VCC.n5553 0.0112143
R10070 VCC.n6009 VCC.n5602 0.0112143
R10071 VCC.n5868 VCC.n5867 0.0112143
R10072 VCC.n5984 VCC.n5983 0.0112143
R10073 VCC.n5874 VCC.n5873 0.0112143
R10074 VCC.n5866 VCC.n5864 0.0112143
R10075 VCC.n5982 VCC.n5616 0.0112143
R10076 VCC.n5744 VCC.n5730 0.0112143
R10077 VCC.n5848 VCC.n5680 0.0112143
R10078 VCC.n5856 VCC.n5855 0.0112143
R10079 VCC.n5743 VCC.n5731 0.0112143
R10080 VCC.n5847 VCC.n5846 0.0112143
R10081 VCC.n5845 VCC.n5681 0.0112143
R10082 VCC.n6294 VCC.n6280 0.0112143
R10083 VCC.n6398 VCC.n6230 0.0112143
R10084 VCC.n6406 VCC.n6405 0.0112143
R10085 VCC.n6293 VCC.n6281 0.0112143
R10086 VCC.n6397 VCC.n6396 0.0112143
R10087 VCC.n6395 VCC.n6231 0.0112143
R10088 VCC.n6419 VCC.n6418 0.0112143
R10089 VCC.n6534 VCC.n6533 0.0112143
R10090 VCC.n6425 VCC.n6424 0.0112143
R10091 VCC.n6417 VCC.n6416 0.0112143
R10092 VCC.n6532 VCC.n6167 0.0112143
R10093 VCC.n6548 VCC.n6547 0.0112143
R10094 VCC.n6562 VCC.n6154 0.0112143
R10095 VCC.n6628 VCC.n6627 0.0112143
R10096 VCC.n6561 VCC.n6560 0.0112143
R10097 VCC.n7105 VCC.n7104 0.0112143
R10098 VCC.n7118 VCC.n7117 0.0112143
R10099 VCC.n7189 VCC.n6660 0.0112143
R10100 VCC.n7116 VCC.n6709 0.0112143
R10101 VCC.n6975 VCC.n6974 0.0112143
R10102 VCC.n7091 VCC.n7090 0.0112143
R10103 VCC.n6981 VCC.n6980 0.0112143
R10104 VCC.n6973 VCC.n6971 0.0112143
R10105 VCC.n7089 VCC.n6723 0.0112143
R10106 VCC.n6851 VCC.n6837 0.0112143
R10107 VCC.n6955 VCC.n6787 0.0112143
R10108 VCC.n6963 VCC.n6962 0.0112143
R10109 VCC.n6850 VCC.n6838 0.0112143
R10110 VCC.n6954 VCC.n6953 0.0112143
R10111 VCC.n6952 VCC.n6788 0.0112143
R10112 VCC.n7401 VCC.n7387 0.0112143
R10113 VCC.n7505 VCC.n7337 0.0112143
R10114 VCC.n7513 VCC.n7512 0.0112143
R10115 VCC.n7400 VCC.n7388 0.0112143
R10116 VCC.n7504 VCC.n7503 0.0112143
R10117 VCC.n7502 VCC.n7338 0.0112143
R10118 VCC.n7526 VCC.n7525 0.0112143
R10119 VCC.n7641 VCC.n7640 0.0112143
R10120 VCC.n7532 VCC.n7531 0.0112143
R10121 VCC.n7524 VCC.n7523 0.0112143
R10122 VCC.n7639 VCC.n7274 0.0112143
R10123 VCC.n7655 VCC.n7654 0.0112143
R10124 VCC.n7669 VCC.n7261 0.0112143
R10125 VCC.n7735 VCC.n7734 0.0112143
R10126 VCC.n7668 VCC.n7667 0.0112143
R10127 VCC.n8212 VCC.n8211 0.0112143
R10128 VCC.n8225 VCC.n8224 0.0112143
R10129 VCC.n8296 VCC.n7767 0.0112143
R10130 VCC.n8223 VCC.n7816 0.0112143
R10131 VCC.n8082 VCC.n8081 0.0112143
R10132 VCC.n8198 VCC.n8197 0.0112143
R10133 VCC.n8088 VCC.n8087 0.0112143
R10134 VCC.n8080 VCC.n8078 0.0112143
R10135 VCC.n8196 VCC.n7830 0.0112143
R10136 VCC.n7958 VCC.n7944 0.0112143
R10137 VCC.n8062 VCC.n7894 0.0112143
R10138 VCC.n8070 VCC.n8069 0.0112143
R10139 VCC.n7957 VCC.n7945 0.0112143
R10140 VCC.n8061 VCC.n8060 0.0112143
R10141 VCC.n8059 VCC.n7895 0.0112143
R10142 VCC.n8446 VCC.n8445 0.0112143
R10143 VCC.n8561 VCC.n8560 0.0112143
R10144 VCC.n8452 VCC.n8451 0.0112143
R10145 VCC.n8444 VCC.n8443 0.0112143
R10146 VCC.n8559 VCC.n8381 0.0112143
R10147 VCC.n8575 VCC.n8574 0.0112143
R10148 VCC.n8589 VCC.n8368 0.0112143
R10149 VCC.n8655 VCC.n8654 0.0112143
R10150 VCC.n8588 VCC.n8587 0.0112143
R10151 VCC.n200 VCC.n199 0.0103214
R10152 VCC.n235 VCC.n170 0.0103214
R10153 VCC.n161 VCC.n158 0.0103214
R10154 VCC.n278 VCC.n277 0.0103214
R10155 VCC.n304 VCC.n303 0.0103214
R10156 VCC.n198 VCC.n197 0.0103214
R10157 VCC.n234 VCC.n171 0.0103214
R10158 VCC.n279 VCC.n149 0.0103214
R10159 VCC.n302 VCC.n133 0.0103214
R10160 VCC.n136 VCC.n130 0.0103214
R10161 VCC.n332 VCC.n331 0.0103214
R10162 VCC.n323 VCC.n116 0.0103214
R10163 VCC.n351 VCC.n350 0.0103214
R10164 VCC.n390 VCC.n389 0.0103214
R10165 VCC.n405 VCC.n404 0.0103214
R10166 VCC.n438 VCC.n74 0.0103214
R10167 VCC.n330 VCC.n319 0.0103214
R10168 VCC.n322 VCC.n115 0.0103214
R10169 VCC.n349 VCC.n103 0.0103214
R10170 VCC.n406 VCC.n89 0.0103214
R10171 VCC.n437 VCC.n436 0.0103214
R10172 VCC.n467 VCC.n58 0.0103214
R10173 VCC.n463 VCC.n462 0.0103214
R10174 VCC.n488 VCC.n45 0.0103214
R10175 VCC.n510 VCC.n26 0.0103214
R10176 VCC.n543 VCC.n542 0.0103214
R10177 VCC.n466 VCC.n60 0.0103214
R10178 VCC.n487 VCC.n486 0.0103214
R10179 VCC.n482 VCC.n36 0.0103214
R10180 VCC.n511 VCC.n28 0.0103214
R10181 VCC.n519 VCC.n518 0.0103214
R10182 VCC.n752 VCC.n751 0.0103214
R10183 VCC.n787 VCC.n722 0.0103214
R10184 VCC.n713 VCC.n710 0.0103214
R10185 VCC.n830 VCC.n829 0.0103214
R10186 VCC.n856 VCC.n855 0.0103214
R10187 VCC.n750 VCC.n749 0.0103214
R10188 VCC.n786 VCC.n723 0.0103214
R10189 VCC.n831 VCC.n701 0.0103214
R10190 VCC.n854 VCC.n685 0.0103214
R10191 VCC.n688 VCC.n682 0.0103214
R10192 VCC.n884 VCC.n883 0.0103214
R10193 VCC.n875 VCC.n668 0.0103214
R10194 VCC.n903 VCC.n902 0.0103214
R10195 VCC.n942 VCC.n941 0.0103214
R10196 VCC.n957 VCC.n956 0.0103214
R10197 VCC.n990 VCC.n626 0.0103214
R10198 VCC.n882 VCC.n871 0.0103214
R10199 VCC.n874 VCC.n667 0.0103214
R10200 VCC.n901 VCC.n655 0.0103214
R10201 VCC.n958 VCC.n641 0.0103214
R10202 VCC.n989 VCC.n988 0.0103214
R10203 VCC.n1019 VCC.n610 0.0103214
R10204 VCC.n1015 VCC.n1014 0.0103214
R10205 VCC.n1040 VCC.n597 0.0103214
R10206 VCC.n1062 VCC.n578 0.0103214
R10207 VCC.n1097 VCC.n1096 0.0103214
R10208 VCC.n1018 VCC.n612 0.0103214
R10209 VCC.n1039 VCC.n1038 0.0103214
R10210 VCC.n1034 VCC.n588 0.0103214
R10211 VCC.n1063 VCC.n580 0.0103214
R10212 VCC.n1071 VCC.n1070 0.0103214
R10213 VCC.n1576 VCC.n1166 0.0103214
R10214 VCC.n1169 VCC.n1168 0.0103214
R10215 VCC.n1589 VCC.n1152 0.0103214
R10216 VCC.n1626 VCC.n1625 0.0103214
R10217 VCC.n1642 VCC.n1125 0.0103214
R10218 VCC.n1564 VCC.n1167 0.0103214
R10219 VCC.n1590 VCC.n1153 0.0103214
R10220 VCC.n1606 VCC.n1151 0.0103214
R10221 VCC.n1627 VCC.n1132 0.0103214
R10222 VCC.n1137 VCC.n1129 0.0103214
R10223 VCC.n1441 VCC.n1235 0.0103214
R10224 VCC.n1432 VCC.n1225 0.0103214
R10225 VCC.n1460 VCC.n1459 0.0103214
R10226 VCC.n1499 VCC.n1498 0.0103214
R10227 VCC.n1514 VCC.n1513 0.0103214
R10228 VCC.n1548 VCC.n1183 0.0103214
R10229 VCC.n1440 VCC.n1439 0.0103214
R10230 VCC.n1431 VCC.n1224 0.0103214
R10231 VCC.n1458 VCC.n1212 0.0103214
R10232 VCC.n1515 VCC.n1198 0.0103214
R10233 VCC.n1547 VCC.n1546 0.0103214
R10234 VCC.n1310 VCC.n1309 0.0103214
R10235 VCC.n1345 VCC.n1280 0.0103214
R10236 VCC.n1271 VCC.n1268 0.0103214
R10237 VCC.n1388 VCC.n1387 0.0103214
R10238 VCC.n1414 VCC.n1413 0.0103214
R10239 VCC.n1308 VCC.n1307 0.0103214
R10240 VCC.n1344 VCC.n1281 0.0103214
R10241 VCC.n1389 VCC.n1259 0.0103214
R10242 VCC.n1412 VCC.n1243 0.0103214
R10243 VCC.n1246 VCC.n1240 0.0103214
R10244 VCC.n1861 VCC.n1860 0.0103214
R10245 VCC.n1896 VCC.n1831 0.0103214
R10246 VCC.n1822 VCC.n1819 0.0103214
R10247 VCC.n1939 VCC.n1938 0.0103214
R10248 VCC.n1965 VCC.n1964 0.0103214
R10249 VCC.n1859 VCC.n1858 0.0103214
R10250 VCC.n1895 VCC.n1832 0.0103214
R10251 VCC.n1940 VCC.n1810 0.0103214
R10252 VCC.n1963 VCC.n1794 0.0103214
R10253 VCC.n1797 VCC.n1791 0.0103214
R10254 VCC.n1993 VCC.n1992 0.0103214
R10255 VCC.n1984 VCC.n1777 0.0103214
R10256 VCC.n2012 VCC.n2011 0.0103214
R10257 VCC.n2051 VCC.n2050 0.0103214
R10258 VCC.n2066 VCC.n2065 0.0103214
R10259 VCC.n2099 VCC.n1735 0.0103214
R10260 VCC.n1991 VCC.n1980 0.0103214
R10261 VCC.n1983 VCC.n1776 0.0103214
R10262 VCC.n2010 VCC.n1764 0.0103214
R10263 VCC.n2067 VCC.n1750 0.0103214
R10264 VCC.n2098 VCC.n2097 0.0103214
R10265 VCC.n2128 VCC.n1719 0.0103214
R10266 VCC.n2124 VCC.n2123 0.0103214
R10267 VCC.n2149 VCC.n1706 0.0103214
R10268 VCC.n2171 VCC.n1687 0.0103214
R10269 VCC.n2206 VCC.n2205 0.0103214
R10270 VCC.n2127 VCC.n1721 0.0103214
R10271 VCC.n2148 VCC.n2147 0.0103214
R10272 VCC.n2143 VCC.n1697 0.0103214
R10273 VCC.n2172 VCC.n1689 0.0103214
R10274 VCC.n2180 VCC.n2179 0.0103214
R10275 VCC.n2685 VCC.n2275 0.0103214
R10276 VCC.n2278 VCC.n2277 0.0103214
R10277 VCC.n2698 VCC.n2261 0.0103214
R10278 VCC.n2735 VCC.n2734 0.0103214
R10279 VCC.n2751 VCC.n2234 0.0103214
R10280 VCC.n2673 VCC.n2276 0.0103214
R10281 VCC.n2699 VCC.n2262 0.0103214
R10282 VCC.n2715 VCC.n2260 0.0103214
R10283 VCC.n2736 VCC.n2241 0.0103214
R10284 VCC.n2246 VCC.n2238 0.0103214
R10285 VCC.n2550 VCC.n2344 0.0103214
R10286 VCC.n2541 VCC.n2334 0.0103214
R10287 VCC.n2569 VCC.n2568 0.0103214
R10288 VCC.n2608 VCC.n2607 0.0103214
R10289 VCC.n2623 VCC.n2622 0.0103214
R10290 VCC.n2657 VCC.n2292 0.0103214
R10291 VCC.n2549 VCC.n2548 0.0103214
R10292 VCC.n2540 VCC.n2333 0.0103214
R10293 VCC.n2567 VCC.n2321 0.0103214
R10294 VCC.n2624 VCC.n2307 0.0103214
R10295 VCC.n2656 VCC.n2655 0.0103214
R10296 VCC.n2419 VCC.n2418 0.0103214
R10297 VCC.n2454 VCC.n2389 0.0103214
R10298 VCC.n2380 VCC.n2377 0.0103214
R10299 VCC.n2497 VCC.n2496 0.0103214
R10300 VCC.n2523 VCC.n2522 0.0103214
R10301 VCC.n2417 VCC.n2416 0.0103214
R10302 VCC.n2453 VCC.n2390 0.0103214
R10303 VCC.n2498 VCC.n2368 0.0103214
R10304 VCC.n2521 VCC.n2352 0.0103214
R10305 VCC.n2355 VCC.n2349 0.0103214
R10306 VCC.n2970 VCC.n2969 0.0103214
R10307 VCC.n3005 VCC.n2940 0.0103214
R10308 VCC.n2931 VCC.n2928 0.0103214
R10309 VCC.n3048 VCC.n3047 0.0103214
R10310 VCC.n3074 VCC.n3073 0.0103214
R10311 VCC.n2968 VCC.n2967 0.0103214
R10312 VCC.n3004 VCC.n2941 0.0103214
R10313 VCC.n3049 VCC.n2919 0.0103214
R10314 VCC.n3072 VCC.n2903 0.0103214
R10315 VCC.n2906 VCC.n2900 0.0103214
R10316 VCC.n3102 VCC.n3101 0.0103214
R10317 VCC.n3093 VCC.n2886 0.0103214
R10318 VCC.n3121 VCC.n3120 0.0103214
R10319 VCC.n3160 VCC.n3159 0.0103214
R10320 VCC.n3175 VCC.n3174 0.0103214
R10321 VCC.n3208 VCC.n2844 0.0103214
R10322 VCC.n3100 VCC.n3089 0.0103214
R10323 VCC.n3092 VCC.n2885 0.0103214
R10324 VCC.n3119 VCC.n2873 0.0103214
R10325 VCC.n3176 VCC.n2859 0.0103214
R10326 VCC.n3207 VCC.n3206 0.0103214
R10327 VCC.n3237 VCC.n2828 0.0103214
R10328 VCC.n3233 VCC.n3232 0.0103214
R10329 VCC.n3258 VCC.n2815 0.0103214
R10330 VCC.n3280 VCC.n2796 0.0103214
R10331 VCC.n3315 VCC.n3314 0.0103214
R10332 VCC.n3236 VCC.n2830 0.0103214
R10333 VCC.n3257 VCC.n3256 0.0103214
R10334 VCC.n3252 VCC.n2806 0.0103214
R10335 VCC.n3281 VCC.n2798 0.0103214
R10336 VCC.n3289 VCC.n3288 0.0103214
R10337 VCC.n3794 VCC.n3384 0.0103214
R10338 VCC.n3387 VCC.n3386 0.0103214
R10339 VCC.n3807 VCC.n3370 0.0103214
R10340 VCC.n3844 VCC.n3843 0.0103214
R10341 VCC.n3860 VCC.n3343 0.0103214
R10342 VCC.n3782 VCC.n3385 0.0103214
R10343 VCC.n3808 VCC.n3371 0.0103214
R10344 VCC.n3824 VCC.n3369 0.0103214
R10345 VCC.n3845 VCC.n3350 0.0103214
R10346 VCC.n3355 VCC.n3347 0.0103214
R10347 VCC.n3659 VCC.n3453 0.0103214
R10348 VCC.n3650 VCC.n3443 0.0103214
R10349 VCC.n3678 VCC.n3677 0.0103214
R10350 VCC.n3717 VCC.n3716 0.0103214
R10351 VCC.n3732 VCC.n3731 0.0103214
R10352 VCC.n3766 VCC.n3401 0.0103214
R10353 VCC.n3658 VCC.n3657 0.0103214
R10354 VCC.n3649 VCC.n3442 0.0103214
R10355 VCC.n3676 VCC.n3430 0.0103214
R10356 VCC.n3733 VCC.n3416 0.0103214
R10357 VCC.n3765 VCC.n3764 0.0103214
R10358 VCC.n3528 VCC.n3527 0.0103214
R10359 VCC.n3563 VCC.n3498 0.0103214
R10360 VCC.n3489 VCC.n3486 0.0103214
R10361 VCC.n3606 VCC.n3605 0.0103214
R10362 VCC.n3632 VCC.n3631 0.0103214
R10363 VCC.n3526 VCC.n3525 0.0103214
R10364 VCC.n3562 VCC.n3499 0.0103214
R10365 VCC.n3607 VCC.n3477 0.0103214
R10366 VCC.n3630 VCC.n3461 0.0103214
R10367 VCC.n3464 VCC.n3458 0.0103214
R10368 VCC.n4079 VCC.n4078 0.0103214
R10369 VCC.n4114 VCC.n4049 0.0103214
R10370 VCC.n4040 VCC.n4037 0.0103214
R10371 VCC.n4157 VCC.n4156 0.0103214
R10372 VCC.n4183 VCC.n4182 0.0103214
R10373 VCC.n4077 VCC.n4076 0.0103214
R10374 VCC.n4113 VCC.n4050 0.0103214
R10375 VCC.n4158 VCC.n4028 0.0103214
R10376 VCC.n4181 VCC.n4012 0.0103214
R10377 VCC.n4015 VCC.n4009 0.0103214
R10378 VCC.n4211 VCC.n4210 0.0103214
R10379 VCC.n4202 VCC.n3995 0.0103214
R10380 VCC.n4230 VCC.n4229 0.0103214
R10381 VCC.n4269 VCC.n4268 0.0103214
R10382 VCC.n4284 VCC.n4283 0.0103214
R10383 VCC.n4317 VCC.n3953 0.0103214
R10384 VCC.n4209 VCC.n4198 0.0103214
R10385 VCC.n4201 VCC.n3994 0.0103214
R10386 VCC.n4228 VCC.n3982 0.0103214
R10387 VCC.n4285 VCC.n3968 0.0103214
R10388 VCC.n4316 VCC.n4315 0.0103214
R10389 VCC.n4346 VCC.n3937 0.0103214
R10390 VCC.n4342 VCC.n4341 0.0103214
R10391 VCC.n4367 VCC.n3924 0.0103214
R10392 VCC.n4389 VCC.n3905 0.0103214
R10393 VCC.n4424 VCC.n4423 0.0103214
R10394 VCC.n4345 VCC.n3939 0.0103214
R10395 VCC.n4366 VCC.n4365 0.0103214
R10396 VCC.n4361 VCC.n3915 0.0103214
R10397 VCC.n4390 VCC.n3907 0.0103214
R10398 VCC.n4398 VCC.n4397 0.0103214
R10399 VCC.n4903 VCC.n4493 0.0103214
R10400 VCC.n4496 VCC.n4495 0.0103214
R10401 VCC.n4916 VCC.n4479 0.0103214
R10402 VCC.n4953 VCC.n4952 0.0103214
R10403 VCC.n4969 VCC.n4452 0.0103214
R10404 VCC.n4891 VCC.n4494 0.0103214
R10405 VCC.n4917 VCC.n4480 0.0103214
R10406 VCC.n4933 VCC.n4478 0.0103214
R10407 VCC.n4954 VCC.n4459 0.0103214
R10408 VCC.n4464 VCC.n4456 0.0103214
R10409 VCC.n4768 VCC.n4562 0.0103214
R10410 VCC.n4759 VCC.n4552 0.0103214
R10411 VCC.n4787 VCC.n4786 0.0103214
R10412 VCC.n4826 VCC.n4825 0.0103214
R10413 VCC.n4841 VCC.n4840 0.0103214
R10414 VCC.n4875 VCC.n4510 0.0103214
R10415 VCC.n4767 VCC.n4766 0.0103214
R10416 VCC.n4758 VCC.n4551 0.0103214
R10417 VCC.n4785 VCC.n4539 0.0103214
R10418 VCC.n4842 VCC.n4525 0.0103214
R10419 VCC.n4874 VCC.n4873 0.0103214
R10420 VCC.n4637 VCC.n4636 0.0103214
R10421 VCC.n4672 VCC.n4607 0.0103214
R10422 VCC.n4598 VCC.n4595 0.0103214
R10423 VCC.n4715 VCC.n4714 0.0103214
R10424 VCC.n4741 VCC.n4740 0.0103214
R10425 VCC.n4635 VCC.n4634 0.0103214
R10426 VCC.n4671 VCC.n4608 0.0103214
R10427 VCC.n4716 VCC.n4586 0.0103214
R10428 VCC.n4739 VCC.n4570 0.0103214
R10429 VCC.n4573 VCC.n4567 0.0103214
R10430 VCC.n5188 VCC.n5187 0.0103214
R10431 VCC.n5223 VCC.n5158 0.0103214
R10432 VCC.n5149 VCC.n5146 0.0103214
R10433 VCC.n5266 VCC.n5265 0.0103214
R10434 VCC.n5292 VCC.n5291 0.0103214
R10435 VCC.n5186 VCC.n5185 0.0103214
R10436 VCC.n5222 VCC.n5159 0.0103214
R10437 VCC.n5267 VCC.n5137 0.0103214
R10438 VCC.n5290 VCC.n5121 0.0103214
R10439 VCC.n5124 VCC.n5118 0.0103214
R10440 VCC.n5320 VCC.n5319 0.0103214
R10441 VCC.n5311 VCC.n5104 0.0103214
R10442 VCC.n5339 VCC.n5338 0.0103214
R10443 VCC.n5378 VCC.n5377 0.0103214
R10444 VCC.n5393 VCC.n5392 0.0103214
R10445 VCC.n5426 VCC.n5062 0.0103214
R10446 VCC.n5318 VCC.n5307 0.0103214
R10447 VCC.n5310 VCC.n5103 0.0103214
R10448 VCC.n5337 VCC.n5091 0.0103214
R10449 VCC.n5394 VCC.n5077 0.0103214
R10450 VCC.n5425 VCC.n5424 0.0103214
R10451 VCC.n5455 VCC.n5046 0.0103214
R10452 VCC.n5451 VCC.n5450 0.0103214
R10453 VCC.n5476 VCC.n5033 0.0103214
R10454 VCC.n5498 VCC.n5014 0.0103214
R10455 VCC.n5533 VCC.n5532 0.0103214
R10456 VCC.n5454 VCC.n5048 0.0103214
R10457 VCC.n5475 VCC.n5474 0.0103214
R10458 VCC.n5470 VCC.n5024 0.0103214
R10459 VCC.n5499 VCC.n5016 0.0103214
R10460 VCC.n5507 VCC.n5506 0.0103214
R10461 VCC.n6011 VCC.n5601 0.0103214
R10462 VCC.n5604 VCC.n5603 0.0103214
R10463 VCC.n6024 VCC.n5587 0.0103214
R10464 VCC.n6061 VCC.n6060 0.0103214
R10465 VCC.n6077 VCC.n5560 0.0103214
R10466 VCC.n5999 VCC.n5602 0.0103214
R10467 VCC.n6025 VCC.n5588 0.0103214
R10468 VCC.n6041 VCC.n5586 0.0103214
R10469 VCC.n6062 VCC.n5567 0.0103214
R10470 VCC.n5572 VCC.n5564 0.0103214
R10471 VCC.n5876 VCC.n5670 0.0103214
R10472 VCC.n5867 VCC.n5660 0.0103214
R10473 VCC.n5895 VCC.n5894 0.0103214
R10474 VCC.n5934 VCC.n5933 0.0103214
R10475 VCC.n5949 VCC.n5948 0.0103214
R10476 VCC.n5983 VCC.n5618 0.0103214
R10477 VCC.n5875 VCC.n5874 0.0103214
R10478 VCC.n5866 VCC.n5659 0.0103214
R10479 VCC.n5893 VCC.n5647 0.0103214
R10480 VCC.n5950 VCC.n5633 0.0103214
R10481 VCC.n5982 VCC.n5981 0.0103214
R10482 VCC.n5745 VCC.n5744 0.0103214
R10483 VCC.n5780 VCC.n5715 0.0103214
R10484 VCC.n5706 VCC.n5703 0.0103214
R10485 VCC.n5823 VCC.n5822 0.0103214
R10486 VCC.n5849 VCC.n5848 0.0103214
R10487 VCC.n5743 VCC.n5742 0.0103214
R10488 VCC.n5779 VCC.n5716 0.0103214
R10489 VCC.n5824 VCC.n5694 0.0103214
R10490 VCC.n5847 VCC.n5678 0.0103214
R10491 VCC.n5681 VCC.n5675 0.0103214
R10492 VCC.n6295 VCC.n6294 0.0103214
R10493 VCC.n6330 VCC.n6265 0.0103214
R10494 VCC.n6256 VCC.n6253 0.0103214
R10495 VCC.n6373 VCC.n6372 0.0103214
R10496 VCC.n6399 VCC.n6398 0.0103214
R10497 VCC.n6293 VCC.n6292 0.0103214
R10498 VCC.n6329 VCC.n6266 0.0103214
R10499 VCC.n6374 VCC.n6244 0.0103214
R10500 VCC.n6397 VCC.n6228 0.0103214
R10501 VCC.n6231 VCC.n6225 0.0103214
R10502 VCC.n6427 VCC.n6426 0.0103214
R10503 VCC.n6418 VCC.n6211 0.0103214
R10504 VCC.n6446 VCC.n6445 0.0103214
R10505 VCC.n6485 VCC.n6484 0.0103214
R10506 VCC.n6500 VCC.n6499 0.0103214
R10507 VCC.n6533 VCC.n6169 0.0103214
R10508 VCC.n6425 VCC.n6414 0.0103214
R10509 VCC.n6417 VCC.n6210 0.0103214
R10510 VCC.n6444 VCC.n6198 0.0103214
R10511 VCC.n6501 VCC.n6184 0.0103214
R10512 VCC.n6532 VCC.n6531 0.0103214
R10513 VCC.n6562 VCC.n6153 0.0103214
R10514 VCC.n6558 VCC.n6557 0.0103214
R10515 VCC.n6583 VCC.n6140 0.0103214
R10516 VCC.n6605 VCC.n6121 0.0103214
R10517 VCC.n6640 VCC.n6639 0.0103214
R10518 VCC.n6561 VCC.n6155 0.0103214
R10519 VCC.n6582 VCC.n6581 0.0103214
R10520 VCC.n6577 VCC.n6131 0.0103214
R10521 VCC.n6606 VCC.n6123 0.0103214
R10522 VCC.n6614 VCC.n6613 0.0103214
R10523 VCC.n7118 VCC.n6708 0.0103214
R10524 VCC.n6711 VCC.n6710 0.0103214
R10525 VCC.n7131 VCC.n6694 0.0103214
R10526 VCC.n7168 VCC.n7167 0.0103214
R10527 VCC.n7184 VCC.n6667 0.0103214
R10528 VCC.n7106 VCC.n6709 0.0103214
R10529 VCC.n7132 VCC.n6695 0.0103214
R10530 VCC.n7148 VCC.n6693 0.0103214
R10531 VCC.n7169 VCC.n6674 0.0103214
R10532 VCC.n6679 VCC.n6671 0.0103214
R10533 VCC.n6983 VCC.n6777 0.0103214
R10534 VCC.n6974 VCC.n6767 0.0103214
R10535 VCC.n7002 VCC.n7001 0.0103214
R10536 VCC.n7041 VCC.n7040 0.0103214
R10537 VCC.n7056 VCC.n7055 0.0103214
R10538 VCC.n7090 VCC.n6725 0.0103214
R10539 VCC.n6982 VCC.n6981 0.0103214
R10540 VCC.n6973 VCC.n6766 0.0103214
R10541 VCC.n7000 VCC.n6754 0.0103214
R10542 VCC.n7057 VCC.n6740 0.0103214
R10543 VCC.n7089 VCC.n7088 0.0103214
R10544 VCC.n6852 VCC.n6851 0.0103214
R10545 VCC.n6887 VCC.n6822 0.0103214
R10546 VCC.n6813 VCC.n6810 0.0103214
R10547 VCC.n6930 VCC.n6929 0.0103214
R10548 VCC.n6956 VCC.n6955 0.0103214
R10549 VCC.n6850 VCC.n6849 0.0103214
R10550 VCC.n6886 VCC.n6823 0.0103214
R10551 VCC.n6931 VCC.n6801 0.0103214
R10552 VCC.n6954 VCC.n6785 0.0103214
R10553 VCC.n6788 VCC.n6782 0.0103214
R10554 VCC.n7402 VCC.n7401 0.0103214
R10555 VCC.n7437 VCC.n7372 0.0103214
R10556 VCC.n7363 VCC.n7360 0.0103214
R10557 VCC.n7480 VCC.n7479 0.0103214
R10558 VCC.n7506 VCC.n7505 0.0103214
R10559 VCC.n7400 VCC.n7399 0.0103214
R10560 VCC.n7436 VCC.n7373 0.0103214
R10561 VCC.n7481 VCC.n7351 0.0103214
R10562 VCC.n7504 VCC.n7335 0.0103214
R10563 VCC.n7338 VCC.n7332 0.0103214
R10564 VCC.n7534 VCC.n7533 0.0103214
R10565 VCC.n7525 VCC.n7318 0.0103214
R10566 VCC.n7553 VCC.n7552 0.0103214
R10567 VCC.n7592 VCC.n7591 0.0103214
R10568 VCC.n7607 VCC.n7606 0.0103214
R10569 VCC.n7640 VCC.n7276 0.0103214
R10570 VCC.n7532 VCC.n7521 0.0103214
R10571 VCC.n7524 VCC.n7317 0.0103214
R10572 VCC.n7551 VCC.n7305 0.0103214
R10573 VCC.n7608 VCC.n7291 0.0103214
R10574 VCC.n7639 VCC.n7638 0.0103214
R10575 VCC.n7669 VCC.n7260 0.0103214
R10576 VCC.n7665 VCC.n7664 0.0103214
R10577 VCC.n7690 VCC.n7247 0.0103214
R10578 VCC.n7712 VCC.n7228 0.0103214
R10579 VCC.n7747 VCC.n7746 0.0103214
R10580 VCC.n7668 VCC.n7262 0.0103214
R10581 VCC.n7689 VCC.n7688 0.0103214
R10582 VCC.n7684 VCC.n7238 0.0103214
R10583 VCC.n7713 VCC.n7230 0.0103214
R10584 VCC.n7721 VCC.n7720 0.0103214
R10585 VCC.n8225 VCC.n7815 0.0103214
R10586 VCC.n7818 VCC.n7817 0.0103214
R10587 VCC.n8238 VCC.n7801 0.0103214
R10588 VCC.n8275 VCC.n8274 0.0103214
R10589 VCC.n8291 VCC.n7774 0.0103214
R10590 VCC.n8213 VCC.n7816 0.0103214
R10591 VCC.n8239 VCC.n7802 0.0103214
R10592 VCC.n8255 VCC.n7800 0.0103214
R10593 VCC.n8276 VCC.n7781 0.0103214
R10594 VCC.n7786 VCC.n7778 0.0103214
R10595 VCC.n8090 VCC.n7884 0.0103214
R10596 VCC.n8081 VCC.n7874 0.0103214
R10597 VCC.n8109 VCC.n8108 0.0103214
R10598 VCC.n8148 VCC.n8147 0.0103214
R10599 VCC.n8163 VCC.n8162 0.0103214
R10600 VCC.n8197 VCC.n7832 0.0103214
R10601 VCC.n8089 VCC.n8088 0.0103214
R10602 VCC.n8080 VCC.n7873 0.0103214
R10603 VCC.n8107 VCC.n7861 0.0103214
R10604 VCC.n8164 VCC.n7847 0.0103214
R10605 VCC.n8196 VCC.n8195 0.0103214
R10606 VCC.n7959 VCC.n7958 0.0103214
R10607 VCC.n7994 VCC.n7929 0.0103214
R10608 VCC.n7920 VCC.n7917 0.0103214
R10609 VCC.n8037 VCC.n8036 0.0103214
R10610 VCC.n8063 VCC.n8062 0.0103214
R10611 VCC.n7957 VCC.n7956 0.0103214
R10612 VCC.n7993 VCC.n7930 0.0103214
R10613 VCC.n8038 VCC.n7908 0.0103214
R10614 VCC.n8061 VCC.n7892 0.0103214
R10615 VCC.n7895 VCC.n7889 0.0103214
R10616 VCC.n8454 VCC.n8453 0.0103214
R10617 VCC.n8445 VCC.n8425 0.0103214
R10618 VCC.n8473 VCC.n8472 0.0103214
R10619 VCC.n8512 VCC.n8511 0.0103214
R10620 VCC.n8527 VCC.n8526 0.0103214
R10621 VCC.n8560 VCC.n8383 0.0103214
R10622 VCC.n8452 VCC.n8441 0.0103214
R10623 VCC.n8444 VCC.n8424 0.0103214
R10624 VCC.n8471 VCC.n8412 0.0103214
R10625 VCC.n8528 VCC.n8398 0.0103214
R10626 VCC.n8559 VCC.n8558 0.0103214
R10627 VCC.n8589 VCC.n8367 0.0103214
R10628 VCC.n8585 VCC.n8584 0.0103214
R10629 VCC.n8610 VCC.n8354 0.0103214
R10630 VCC.n8632 VCC.n8335 0.0103214
R10631 VCC.n8667 VCC.n8666 0.0103214
R10632 VCC.n8588 VCC.n8369 0.0103214
R10633 VCC.n8609 VCC.n8608 0.0103214
R10634 VCC.n8604 VCC.n8345 0.0103214
R10635 VCC.n8633 VCC.n8337 0.0103214
R10636 VCC.n8641 VCC.n8640 0.0103214
R10637 VCC.n206 VCC.n193 0.00942857
R10638 VCC.n246 VCC.n168 0.00942857
R10639 VCC.n262 VCC.n162 0.00942857
R10640 VCC.n294 VCC.n138 0.00942857
R10641 VCC.n205 VCC.n190 0.00942857
R10642 VCC.n261 VCC.n260 0.00942857
R10643 VCC.n367 VCC.n105 0.00942857
R10644 VCC.n383 VCC.n98 0.00942857
R10645 VCC.n77 VCC.n68 0.00942857
R10646 VCC.n382 VCC.n100 0.00942857
R10647 VCC.n75 VCC.n69 0.00942857
R10648 VCC.n457 VCC.n456 0.00942857
R10649 VCC.n534 VCC.n16 0.00942857
R10650 VCC.n19 VCC.n17 0.00942857
R10651 VCC.n455 VCC.n64 0.00942857
R10652 VCC.n479 VCC.n51 0.00942857
R10653 VCC.n507 VCC.n506 0.00942857
R10654 VCC.n18 VCC.n10 0.00942857
R10655 VCC.n758 VCC.n745 0.00942857
R10656 VCC.n798 VCC.n720 0.00942857
R10657 VCC.n814 VCC.n714 0.00942857
R10658 VCC.n846 VCC.n690 0.00942857
R10659 VCC.n757 VCC.n742 0.00942857
R10660 VCC.n813 VCC.n812 0.00942857
R10661 VCC.n919 VCC.n657 0.00942857
R10662 VCC.n935 VCC.n650 0.00942857
R10663 VCC.n629 VCC.n620 0.00942857
R10664 VCC.n934 VCC.n652 0.00942857
R10665 VCC.n627 VCC.n621 0.00942857
R10666 VCC.n1009 VCC.n1008 0.00942857
R10667 VCC.n1086 VCC.n568 0.00942857
R10668 VCC.n571 VCC.n569 0.00942857
R10669 VCC.n1007 VCC.n616 0.00942857
R10670 VCC.n1031 VCC.n603 0.00942857
R10671 VCC.n1059 VCC.n1058 0.00942857
R10672 VCC.n570 VCC.n564 0.00942857
R10673 VCC.n1568 VCC.n1567 0.00942857
R10674 VCC.n1633 VCC.n1632 0.00942857
R10675 VCC.n1646 VCC.n1119 0.00942857
R10676 VCC.n1566 VCC.n1173 0.00942857
R10677 VCC.n1597 VCC.n1156 0.00942857
R10678 VCC.n1610 VCC.n1149 0.00942857
R10679 VCC.n1645 VCC.n1644 0.00942857
R10680 VCC.n1476 VCC.n1214 0.00942857
R10681 VCC.n1492 VCC.n1207 0.00942857
R10682 VCC.n1186 VCC.n1177 0.00942857
R10683 VCC.n1491 VCC.n1209 0.00942857
R10684 VCC.n1184 VCC.n1178 0.00942857
R10685 VCC.n1316 VCC.n1303 0.00942857
R10686 VCC.n1356 VCC.n1278 0.00942857
R10687 VCC.n1372 VCC.n1272 0.00942857
R10688 VCC.n1404 VCC.n1248 0.00942857
R10689 VCC.n1315 VCC.n1300 0.00942857
R10690 VCC.n1371 VCC.n1370 0.00942857
R10691 VCC.n1867 VCC.n1854 0.00942857
R10692 VCC.n1907 VCC.n1829 0.00942857
R10693 VCC.n1923 VCC.n1823 0.00942857
R10694 VCC.n1955 VCC.n1799 0.00942857
R10695 VCC.n1866 VCC.n1851 0.00942857
R10696 VCC.n1922 VCC.n1921 0.00942857
R10697 VCC.n2028 VCC.n1766 0.00942857
R10698 VCC.n2044 VCC.n1759 0.00942857
R10699 VCC.n1738 VCC.n1729 0.00942857
R10700 VCC.n2043 VCC.n1761 0.00942857
R10701 VCC.n1736 VCC.n1730 0.00942857
R10702 VCC.n2118 VCC.n2117 0.00942857
R10703 VCC.n2195 VCC.n1677 0.00942857
R10704 VCC.n1680 VCC.n1678 0.00942857
R10705 VCC.n2116 VCC.n1725 0.00942857
R10706 VCC.n2140 VCC.n1712 0.00942857
R10707 VCC.n2168 VCC.n2167 0.00942857
R10708 VCC.n1679 VCC.n1673 0.00942857
R10709 VCC.n2677 VCC.n2676 0.00942857
R10710 VCC.n2742 VCC.n2741 0.00942857
R10711 VCC.n2755 VCC.n2228 0.00942857
R10712 VCC.n2675 VCC.n2282 0.00942857
R10713 VCC.n2706 VCC.n2265 0.00942857
R10714 VCC.n2719 VCC.n2258 0.00942857
R10715 VCC.n2754 VCC.n2753 0.00942857
R10716 VCC.n2585 VCC.n2323 0.00942857
R10717 VCC.n2601 VCC.n2316 0.00942857
R10718 VCC.n2295 VCC.n2286 0.00942857
R10719 VCC.n2600 VCC.n2318 0.00942857
R10720 VCC.n2293 VCC.n2287 0.00942857
R10721 VCC.n2425 VCC.n2412 0.00942857
R10722 VCC.n2465 VCC.n2387 0.00942857
R10723 VCC.n2481 VCC.n2381 0.00942857
R10724 VCC.n2513 VCC.n2357 0.00942857
R10725 VCC.n2424 VCC.n2409 0.00942857
R10726 VCC.n2480 VCC.n2479 0.00942857
R10727 VCC.n2976 VCC.n2963 0.00942857
R10728 VCC.n3016 VCC.n2938 0.00942857
R10729 VCC.n3032 VCC.n2932 0.00942857
R10730 VCC.n3064 VCC.n2908 0.00942857
R10731 VCC.n2975 VCC.n2960 0.00942857
R10732 VCC.n3031 VCC.n3030 0.00942857
R10733 VCC.n3137 VCC.n2875 0.00942857
R10734 VCC.n3153 VCC.n2868 0.00942857
R10735 VCC.n2847 VCC.n2838 0.00942857
R10736 VCC.n3152 VCC.n2870 0.00942857
R10737 VCC.n2845 VCC.n2839 0.00942857
R10738 VCC.n3227 VCC.n3226 0.00942857
R10739 VCC.n3304 VCC.n2786 0.00942857
R10740 VCC.n2789 VCC.n2787 0.00942857
R10741 VCC.n3225 VCC.n2834 0.00942857
R10742 VCC.n3249 VCC.n2821 0.00942857
R10743 VCC.n3277 VCC.n3276 0.00942857
R10744 VCC.n2788 VCC.n2782 0.00942857
R10745 VCC.n3786 VCC.n3785 0.00942857
R10746 VCC.n3851 VCC.n3850 0.00942857
R10747 VCC.n3864 VCC.n3337 0.00942857
R10748 VCC.n3784 VCC.n3391 0.00942857
R10749 VCC.n3815 VCC.n3374 0.00942857
R10750 VCC.n3828 VCC.n3367 0.00942857
R10751 VCC.n3863 VCC.n3862 0.00942857
R10752 VCC.n3694 VCC.n3432 0.00942857
R10753 VCC.n3710 VCC.n3425 0.00942857
R10754 VCC.n3404 VCC.n3395 0.00942857
R10755 VCC.n3709 VCC.n3427 0.00942857
R10756 VCC.n3402 VCC.n3396 0.00942857
R10757 VCC.n3534 VCC.n3521 0.00942857
R10758 VCC.n3574 VCC.n3496 0.00942857
R10759 VCC.n3590 VCC.n3490 0.00942857
R10760 VCC.n3622 VCC.n3466 0.00942857
R10761 VCC.n3533 VCC.n3518 0.00942857
R10762 VCC.n3589 VCC.n3588 0.00942857
R10763 VCC.n4085 VCC.n4072 0.00942857
R10764 VCC.n4125 VCC.n4047 0.00942857
R10765 VCC.n4141 VCC.n4041 0.00942857
R10766 VCC.n4173 VCC.n4017 0.00942857
R10767 VCC.n4084 VCC.n4069 0.00942857
R10768 VCC.n4140 VCC.n4139 0.00942857
R10769 VCC.n4246 VCC.n3984 0.00942857
R10770 VCC.n4262 VCC.n3977 0.00942857
R10771 VCC.n3956 VCC.n3947 0.00942857
R10772 VCC.n4261 VCC.n3979 0.00942857
R10773 VCC.n3954 VCC.n3948 0.00942857
R10774 VCC.n4336 VCC.n4335 0.00942857
R10775 VCC.n4413 VCC.n3895 0.00942857
R10776 VCC.n3898 VCC.n3896 0.00942857
R10777 VCC.n4334 VCC.n3943 0.00942857
R10778 VCC.n4358 VCC.n3930 0.00942857
R10779 VCC.n4386 VCC.n4385 0.00942857
R10780 VCC.n3897 VCC.n3891 0.00942857
R10781 VCC.n4895 VCC.n4894 0.00942857
R10782 VCC.n4960 VCC.n4959 0.00942857
R10783 VCC.n4973 VCC.n4446 0.00942857
R10784 VCC.n4893 VCC.n4500 0.00942857
R10785 VCC.n4924 VCC.n4483 0.00942857
R10786 VCC.n4937 VCC.n4476 0.00942857
R10787 VCC.n4972 VCC.n4971 0.00942857
R10788 VCC.n4803 VCC.n4541 0.00942857
R10789 VCC.n4819 VCC.n4534 0.00942857
R10790 VCC.n4513 VCC.n4504 0.00942857
R10791 VCC.n4818 VCC.n4536 0.00942857
R10792 VCC.n4511 VCC.n4505 0.00942857
R10793 VCC.n4643 VCC.n4630 0.00942857
R10794 VCC.n4683 VCC.n4605 0.00942857
R10795 VCC.n4699 VCC.n4599 0.00942857
R10796 VCC.n4731 VCC.n4575 0.00942857
R10797 VCC.n4642 VCC.n4627 0.00942857
R10798 VCC.n4698 VCC.n4697 0.00942857
R10799 VCC.n5194 VCC.n5181 0.00942857
R10800 VCC.n5234 VCC.n5156 0.00942857
R10801 VCC.n5250 VCC.n5150 0.00942857
R10802 VCC.n5282 VCC.n5126 0.00942857
R10803 VCC.n5193 VCC.n5178 0.00942857
R10804 VCC.n5249 VCC.n5248 0.00942857
R10805 VCC.n5355 VCC.n5093 0.00942857
R10806 VCC.n5371 VCC.n5086 0.00942857
R10807 VCC.n5065 VCC.n5056 0.00942857
R10808 VCC.n5370 VCC.n5088 0.00942857
R10809 VCC.n5063 VCC.n5057 0.00942857
R10810 VCC.n5445 VCC.n5444 0.00942857
R10811 VCC.n5522 VCC.n5004 0.00942857
R10812 VCC.n5007 VCC.n5005 0.00942857
R10813 VCC.n5443 VCC.n5052 0.00942857
R10814 VCC.n5467 VCC.n5039 0.00942857
R10815 VCC.n5495 VCC.n5494 0.00942857
R10816 VCC.n5006 VCC.n5000 0.00942857
R10817 VCC.n6003 VCC.n6002 0.00942857
R10818 VCC.n6068 VCC.n6067 0.00942857
R10819 VCC.n6081 VCC.n5554 0.00942857
R10820 VCC.n6001 VCC.n5608 0.00942857
R10821 VCC.n6032 VCC.n5591 0.00942857
R10822 VCC.n6045 VCC.n5584 0.00942857
R10823 VCC.n6080 VCC.n6079 0.00942857
R10824 VCC.n5911 VCC.n5649 0.00942857
R10825 VCC.n5927 VCC.n5642 0.00942857
R10826 VCC.n5621 VCC.n5612 0.00942857
R10827 VCC.n5926 VCC.n5644 0.00942857
R10828 VCC.n5619 VCC.n5613 0.00942857
R10829 VCC.n5751 VCC.n5738 0.00942857
R10830 VCC.n5791 VCC.n5713 0.00942857
R10831 VCC.n5807 VCC.n5707 0.00942857
R10832 VCC.n5839 VCC.n5683 0.00942857
R10833 VCC.n5750 VCC.n5735 0.00942857
R10834 VCC.n5806 VCC.n5805 0.00942857
R10835 VCC.n6301 VCC.n6288 0.00942857
R10836 VCC.n6341 VCC.n6263 0.00942857
R10837 VCC.n6357 VCC.n6257 0.00942857
R10838 VCC.n6389 VCC.n6233 0.00942857
R10839 VCC.n6300 VCC.n6285 0.00942857
R10840 VCC.n6356 VCC.n6355 0.00942857
R10841 VCC.n6462 VCC.n6200 0.00942857
R10842 VCC.n6478 VCC.n6193 0.00942857
R10843 VCC.n6172 VCC.n6163 0.00942857
R10844 VCC.n6477 VCC.n6195 0.00942857
R10845 VCC.n6170 VCC.n6164 0.00942857
R10846 VCC.n6552 VCC.n6551 0.00942857
R10847 VCC.n6629 VCC.n6111 0.00942857
R10848 VCC.n6114 VCC.n6112 0.00942857
R10849 VCC.n6550 VCC.n6159 0.00942857
R10850 VCC.n6574 VCC.n6146 0.00942857
R10851 VCC.n6602 VCC.n6601 0.00942857
R10852 VCC.n6113 VCC.n6107 0.00942857
R10853 VCC.n7110 VCC.n7109 0.00942857
R10854 VCC.n7175 VCC.n7174 0.00942857
R10855 VCC.n7188 VCC.n6661 0.00942857
R10856 VCC.n7108 VCC.n6715 0.00942857
R10857 VCC.n7139 VCC.n6698 0.00942857
R10858 VCC.n7152 VCC.n6691 0.00942857
R10859 VCC.n7187 VCC.n7186 0.00942857
R10860 VCC.n7018 VCC.n6756 0.00942857
R10861 VCC.n7034 VCC.n6749 0.00942857
R10862 VCC.n6728 VCC.n6719 0.00942857
R10863 VCC.n7033 VCC.n6751 0.00942857
R10864 VCC.n6726 VCC.n6720 0.00942857
R10865 VCC.n6858 VCC.n6845 0.00942857
R10866 VCC.n6898 VCC.n6820 0.00942857
R10867 VCC.n6914 VCC.n6814 0.00942857
R10868 VCC.n6946 VCC.n6790 0.00942857
R10869 VCC.n6857 VCC.n6842 0.00942857
R10870 VCC.n6913 VCC.n6912 0.00942857
R10871 VCC.n7408 VCC.n7395 0.00942857
R10872 VCC.n7448 VCC.n7370 0.00942857
R10873 VCC.n7464 VCC.n7364 0.00942857
R10874 VCC.n7496 VCC.n7340 0.00942857
R10875 VCC.n7407 VCC.n7392 0.00942857
R10876 VCC.n7463 VCC.n7462 0.00942857
R10877 VCC.n7569 VCC.n7307 0.00942857
R10878 VCC.n7585 VCC.n7300 0.00942857
R10879 VCC.n7279 VCC.n7270 0.00942857
R10880 VCC.n7584 VCC.n7302 0.00942857
R10881 VCC.n7277 VCC.n7271 0.00942857
R10882 VCC.n7659 VCC.n7658 0.00942857
R10883 VCC.n7736 VCC.n7218 0.00942857
R10884 VCC.n7221 VCC.n7219 0.00942857
R10885 VCC.n7657 VCC.n7266 0.00942857
R10886 VCC.n7681 VCC.n7253 0.00942857
R10887 VCC.n7709 VCC.n7708 0.00942857
R10888 VCC.n7220 VCC.n7214 0.00942857
R10889 VCC.n8217 VCC.n8216 0.00942857
R10890 VCC.n8282 VCC.n8281 0.00942857
R10891 VCC.n8295 VCC.n7768 0.00942857
R10892 VCC.n8215 VCC.n7822 0.00942857
R10893 VCC.n8246 VCC.n7805 0.00942857
R10894 VCC.n8259 VCC.n7798 0.00942857
R10895 VCC.n8294 VCC.n8293 0.00942857
R10896 VCC.n8125 VCC.n7863 0.00942857
R10897 VCC.n8141 VCC.n7856 0.00942857
R10898 VCC.n7835 VCC.n7826 0.00942857
R10899 VCC.n8140 VCC.n7858 0.00942857
R10900 VCC.n7833 VCC.n7827 0.00942857
R10901 VCC.n7965 VCC.n7952 0.00942857
R10902 VCC.n8005 VCC.n7927 0.00942857
R10903 VCC.n8021 VCC.n7921 0.00942857
R10904 VCC.n8053 VCC.n7897 0.00942857
R10905 VCC.n7964 VCC.n7949 0.00942857
R10906 VCC.n8020 VCC.n8019 0.00942857
R10907 VCC.n8489 VCC.n8414 0.00942857
R10908 VCC.n8505 VCC.n8407 0.00942857
R10909 VCC.n8386 VCC.n8377 0.00942857
R10910 VCC.n8504 VCC.n8409 0.00942857
R10911 VCC.n8384 VCC.n8378 0.00942857
R10912 VCC.n8579 VCC.n8578 0.00942857
R10913 VCC.n8656 VCC.n8325 0.00942857
R10914 VCC.n8328 VCC.n8326 0.00942857
R10915 VCC.n8577 VCC.n8373 0.00942857
R10916 VCC.n8601 VCC.n8360 0.00942857
R10917 VCC.n8629 VCC.n8628 0.00942857
R10918 VCC.n8327 VCC.n8321 0.00942857
R10919 VCC.n222 VCC.n221 0.00853571
R10920 VCC.n233 VCC.n176 0.00853571
R10921 VCC.n251 VCC.n250 0.00853571
R10922 VCC.n284 VCC.n145 0.00853571
R10923 VCC.n172 VCC.n166 0.00853571
R10924 VCC.n342 VCC.n117 0.00853571
R10925 VCC.n356 VCC.n111 0.00853571
R10926 VCC.n388 VCC.n96 0.00853571
R10927 VCC.n411 VCC.n85 0.00853571
R10928 VCC.n375 VCC.n374 0.00853571
R10929 VCC.n478 VCC.n52 0.00853571
R10930 VCC.n540 VCC.n539 0.00853571
R10931 VCC.n551 VCC.n1 0.00853571
R10932 VCC.n774 VCC.n773 0.00853571
R10933 VCC.n785 VCC.n728 0.00853571
R10934 VCC.n803 VCC.n802 0.00853571
R10935 VCC.n836 VCC.n697 0.00853571
R10936 VCC.n724 VCC.n718 0.00853571
R10937 VCC.n894 VCC.n669 0.00853571
R10938 VCC.n908 VCC.n663 0.00853571
R10939 VCC.n940 VCC.n648 0.00853571
R10940 VCC.n963 VCC.n637 0.00853571
R10941 VCC.n927 VCC.n926 0.00853571
R10942 VCC.n1030 VCC.n604 0.00853571
R10943 VCC.n1094 VCC.n1093 0.00853571
R10944 VCC.n1105 VCC.n555 0.00853571
R10945 VCC.n1596 VCC.n1157 0.00853571
R10946 VCC.n1638 VCC.n1121 0.00853571
R10947 VCC.n1659 VCC.n1109 0.00853571
R10948 VCC.n1451 VCC.n1226 0.00853571
R10949 VCC.n1465 VCC.n1220 0.00853571
R10950 VCC.n1497 VCC.n1205 0.00853571
R10951 VCC.n1520 VCC.n1194 0.00853571
R10952 VCC.n1484 VCC.n1483 0.00853571
R10953 VCC.n1332 VCC.n1331 0.00853571
R10954 VCC.n1343 VCC.n1286 0.00853571
R10955 VCC.n1361 VCC.n1360 0.00853571
R10956 VCC.n1394 VCC.n1255 0.00853571
R10957 VCC.n1282 VCC.n1276 0.00853571
R10958 VCC.n1883 VCC.n1882 0.00853571
R10959 VCC.n1894 VCC.n1837 0.00853571
R10960 VCC.n1912 VCC.n1911 0.00853571
R10961 VCC.n1945 VCC.n1806 0.00853571
R10962 VCC.n1833 VCC.n1827 0.00853571
R10963 VCC.n2003 VCC.n1778 0.00853571
R10964 VCC.n2017 VCC.n1772 0.00853571
R10965 VCC.n2049 VCC.n1757 0.00853571
R10966 VCC.n2072 VCC.n1746 0.00853571
R10967 VCC.n2036 VCC.n2035 0.00853571
R10968 VCC.n2139 VCC.n1713 0.00853571
R10969 VCC.n2203 VCC.n2202 0.00853571
R10970 VCC.n2214 VCC.n1664 0.00853571
R10971 VCC.n2705 VCC.n2266 0.00853571
R10972 VCC.n2747 VCC.n2230 0.00853571
R10973 VCC.n2768 VCC.n2218 0.00853571
R10974 VCC.n2560 VCC.n2335 0.00853571
R10975 VCC.n2574 VCC.n2329 0.00853571
R10976 VCC.n2606 VCC.n2314 0.00853571
R10977 VCC.n2629 VCC.n2303 0.00853571
R10978 VCC.n2593 VCC.n2592 0.00853571
R10979 VCC.n2441 VCC.n2440 0.00853571
R10980 VCC.n2452 VCC.n2395 0.00853571
R10981 VCC.n2470 VCC.n2469 0.00853571
R10982 VCC.n2503 VCC.n2364 0.00853571
R10983 VCC.n2391 VCC.n2385 0.00853571
R10984 VCC.n2992 VCC.n2991 0.00853571
R10985 VCC.n3003 VCC.n2946 0.00853571
R10986 VCC.n3021 VCC.n3020 0.00853571
R10987 VCC.n3054 VCC.n2915 0.00853571
R10988 VCC.n2942 VCC.n2936 0.00853571
R10989 VCC.n3112 VCC.n2887 0.00853571
R10990 VCC.n3126 VCC.n2881 0.00853571
R10991 VCC.n3158 VCC.n2866 0.00853571
R10992 VCC.n3181 VCC.n2855 0.00853571
R10993 VCC.n3145 VCC.n3144 0.00853571
R10994 VCC.n3248 VCC.n2822 0.00853571
R10995 VCC.n3312 VCC.n3311 0.00853571
R10996 VCC.n3323 VCC.n2773 0.00853571
R10997 VCC.n3814 VCC.n3375 0.00853571
R10998 VCC.n3856 VCC.n3339 0.00853571
R10999 VCC.n3877 VCC.n3327 0.00853571
R11000 VCC.n3669 VCC.n3444 0.00853571
R11001 VCC.n3683 VCC.n3438 0.00853571
R11002 VCC.n3715 VCC.n3423 0.00853571
R11003 VCC.n3738 VCC.n3412 0.00853571
R11004 VCC.n3702 VCC.n3701 0.00853571
R11005 VCC.n3550 VCC.n3549 0.00853571
R11006 VCC.n3561 VCC.n3504 0.00853571
R11007 VCC.n3579 VCC.n3578 0.00853571
R11008 VCC.n3612 VCC.n3473 0.00853571
R11009 VCC.n3500 VCC.n3494 0.00853571
R11010 VCC.n4101 VCC.n4100 0.00853571
R11011 VCC.n4112 VCC.n4055 0.00853571
R11012 VCC.n4130 VCC.n4129 0.00853571
R11013 VCC.n4163 VCC.n4024 0.00853571
R11014 VCC.n4051 VCC.n4045 0.00853571
R11015 VCC.n4221 VCC.n3996 0.00853571
R11016 VCC.n4235 VCC.n3990 0.00853571
R11017 VCC.n4267 VCC.n3975 0.00853571
R11018 VCC.n4290 VCC.n3964 0.00853571
R11019 VCC.n4254 VCC.n4253 0.00853571
R11020 VCC.n4357 VCC.n3931 0.00853571
R11021 VCC.n4421 VCC.n4420 0.00853571
R11022 VCC.n4432 VCC.n3882 0.00853571
R11023 VCC.n4923 VCC.n4484 0.00853571
R11024 VCC.n4965 VCC.n4448 0.00853571
R11025 VCC.n4986 VCC.n4436 0.00853571
R11026 VCC.n4778 VCC.n4553 0.00853571
R11027 VCC.n4792 VCC.n4547 0.00853571
R11028 VCC.n4824 VCC.n4532 0.00853571
R11029 VCC.n4847 VCC.n4521 0.00853571
R11030 VCC.n4811 VCC.n4810 0.00853571
R11031 VCC.n4659 VCC.n4658 0.00853571
R11032 VCC.n4670 VCC.n4613 0.00853571
R11033 VCC.n4688 VCC.n4687 0.00853571
R11034 VCC.n4721 VCC.n4582 0.00853571
R11035 VCC.n4609 VCC.n4603 0.00853571
R11036 VCC.n5210 VCC.n5209 0.00853571
R11037 VCC.n5221 VCC.n5164 0.00853571
R11038 VCC.n5239 VCC.n5238 0.00853571
R11039 VCC.n5272 VCC.n5133 0.00853571
R11040 VCC.n5160 VCC.n5154 0.00853571
R11041 VCC.n5330 VCC.n5105 0.00853571
R11042 VCC.n5344 VCC.n5099 0.00853571
R11043 VCC.n5376 VCC.n5084 0.00853571
R11044 VCC.n5399 VCC.n5073 0.00853571
R11045 VCC.n5363 VCC.n5362 0.00853571
R11046 VCC.n5466 VCC.n5040 0.00853571
R11047 VCC.n5530 VCC.n5529 0.00853571
R11048 VCC.n5541 VCC.n4991 0.00853571
R11049 VCC.n6031 VCC.n5592 0.00853571
R11050 VCC.n6073 VCC.n5556 0.00853571
R11051 VCC.n6094 VCC.n5544 0.00853571
R11052 VCC.n5886 VCC.n5661 0.00853571
R11053 VCC.n5900 VCC.n5655 0.00853571
R11054 VCC.n5932 VCC.n5640 0.00853571
R11055 VCC.n5955 VCC.n5629 0.00853571
R11056 VCC.n5919 VCC.n5918 0.00853571
R11057 VCC.n5767 VCC.n5766 0.00853571
R11058 VCC.n5778 VCC.n5721 0.00853571
R11059 VCC.n5796 VCC.n5795 0.00853571
R11060 VCC.n5829 VCC.n5690 0.00853571
R11061 VCC.n5717 VCC.n5711 0.00853571
R11062 VCC.n6317 VCC.n6316 0.00853571
R11063 VCC.n6328 VCC.n6271 0.00853571
R11064 VCC.n6346 VCC.n6345 0.00853571
R11065 VCC.n6379 VCC.n6240 0.00853571
R11066 VCC.n6267 VCC.n6261 0.00853571
R11067 VCC.n6437 VCC.n6212 0.00853571
R11068 VCC.n6451 VCC.n6206 0.00853571
R11069 VCC.n6483 VCC.n6191 0.00853571
R11070 VCC.n6506 VCC.n6180 0.00853571
R11071 VCC.n6470 VCC.n6469 0.00853571
R11072 VCC.n6573 VCC.n6147 0.00853571
R11073 VCC.n6637 VCC.n6636 0.00853571
R11074 VCC.n6648 VCC.n6098 0.00853571
R11075 VCC.n7138 VCC.n6699 0.00853571
R11076 VCC.n7180 VCC.n6663 0.00853571
R11077 VCC.n7201 VCC.n6651 0.00853571
R11078 VCC.n6993 VCC.n6768 0.00853571
R11079 VCC.n7007 VCC.n6762 0.00853571
R11080 VCC.n7039 VCC.n6747 0.00853571
R11081 VCC.n7062 VCC.n6736 0.00853571
R11082 VCC.n7026 VCC.n7025 0.00853571
R11083 VCC.n6874 VCC.n6873 0.00853571
R11084 VCC.n6885 VCC.n6828 0.00853571
R11085 VCC.n6903 VCC.n6902 0.00853571
R11086 VCC.n6936 VCC.n6797 0.00853571
R11087 VCC.n6824 VCC.n6818 0.00853571
R11088 VCC.n7424 VCC.n7423 0.00853571
R11089 VCC.n7435 VCC.n7378 0.00853571
R11090 VCC.n7453 VCC.n7452 0.00853571
R11091 VCC.n7486 VCC.n7347 0.00853571
R11092 VCC.n7374 VCC.n7368 0.00853571
R11093 VCC.n7544 VCC.n7319 0.00853571
R11094 VCC.n7558 VCC.n7313 0.00853571
R11095 VCC.n7590 VCC.n7298 0.00853571
R11096 VCC.n7613 VCC.n7287 0.00853571
R11097 VCC.n7577 VCC.n7576 0.00853571
R11098 VCC.n7680 VCC.n7254 0.00853571
R11099 VCC.n7744 VCC.n7743 0.00853571
R11100 VCC.n7755 VCC.n7205 0.00853571
R11101 VCC.n8245 VCC.n7806 0.00853571
R11102 VCC.n8287 VCC.n7770 0.00853571
R11103 VCC.n8308 VCC.n7758 0.00853571
R11104 VCC.n8100 VCC.n7875 0.00853571
R11105 VCC.n8114 VCC.n7869 0.00853571
R11106 VCC.n8146 VCC.n7854 0.00853571
R11107 VCC.n8169 VCC.n7843 0.00853571
R11108 VCC.n8133 VCC.n8132 0.00853571
R11109 VCC.n7981 VCC.n7980 0.00853571
R11110 VCC.n7992 VCC.n7935 0.00853571
R11111 VCC.n8010 VCC.n8009 0.00853571
R11112 VCC.n8043 VCC.n7904 0.00853571
R11113 VCC.n7931 VCC.n7925 0.00853571
R11114 VCC.n8464 VCC.n8426 0.00853571
R11115 VCC.n8478 VCC.n8420 0.00853571
R11116 VCC.n8510 VCC.n8405 0.00853571
R11117 VCC.n8533 VCC.n8394 0.00853571
R11118 VCC.n8497 VCC.n8496 0.00853571
R11119 VCC.n8600 VCC.n8361 0.00853571
R11120 VCC.n8664 VCC.n8663 0.00853571
R11121 VCC.n8675 VCC.n8312 0.00853571
R11122 VCC.n191 VCC.n188 0.00822143
R11123 VCC.n241 VCC.n173 0.00822143
R11124 VCC.n281 VCC.n131 0.00822143
R11125 VCC.n313 VCC.n127 0.00822143
R11126 VCC.n316 VCC.n315 0.00822143
R11127 VCC.n347 VCC.n346 0.00822143
R11128 VCC.n408 VCC.n70 0.00822143
R11129 VCC.n448 VCC.n66 0.00822143
R11130 VCC.n449 VCC.n62 0.00822143
R11131 VCC.n481 VCC.n49 0.00822143
R11132 VCC.n513 VCC.n13 0.00822143
R11133 VCC.n552 VCC.n0 0.00822143
R11134 VCC.n743 VCC.n740 0.00822143
R11135 VCC.n793 VCC.n725 0.00822143
R11136 VCC.n833 VCC.n683 0.00822143
R11137 VCC.n865 VCC.n679 0.00822143
R11138 VCC.n868 VCC.n867 0.00822143
R11139 VCC.n899 VCC.n898 0.00822143
R11140 VCC.n960 VCC.n622 0.00822143
R11141 VCC.n1000 VCC.n618 0.00822143
R11142 VCC.n1001 VCC.n614 0.00822143
R11143 VCC.n1033 VCC.n601 0.00822143
R11144 VCC.n1065 VCC.n565 0.00822143
R11145 VCC.n1106 VCC.n554 0.00822143
R11146 VCC.n1301 VCC.n1298 0.00822143
R11147 VCC.n1351 VCC.n1283 0.00822143
R11148 VCC.n1391 VCC.n1241 0.00822143
R11149 VCC.n1423 VCC.n1237 0.00822143
R11150 VCC.n1426 VCC.n1425 0.00822143
R11151 VCC.n1456 VCC.n1455 0.00822143
R11152 VCC.n1517 VCC.n1179 0.00822143
R11153 VCC.n1558 VCC.n1175 0.00822143
R11154 VCC.n1559 VCC.n1171 0.00822143
R11155 VCC.n1599 VCC.n1154 0.00822143
R11156 VCC.n1629 VCC.n1126 0.00822143
R11157 VCC.n1660 VCC.n1108 0.00822143
R11158 VCC.n1852 VCC.n1849 0.00822143
R11159 VCC.n1902 VCC.n1834 0.00822143
R11160 VCC.n1942 VCC.n1792 0.00822143
R11161 VCC.n1974 VCC.n1788 0.00822143
R11162 VCC.n1977 VCC.n1976 0.00822143
R11163 VCC.n2008 VCC.n2007 0.00822143
R11164 VCC.n2069 VCC.n1731 0.00822143
R11165 VCC.n2109 VCC.n1727 0.00822143
R11166 VCC.n2110 VCC.n1723 0.00822143
R11167 VCC.n2142 VCC.n1710 0.00822143
R11168 VCC.n2174 VCC.n1674 0.00822143
R11169 VCC.n2215 VCC.n1663 0.00822143
R11170 VCC.n2410 VCC.n2407 0.00822143
R11171 VCC.n2460 VCC.n2392 0.00822143
R11172 VCC.n2500 VCC.n2350 0.00822143
R11173 VCC.n2532 VCC.n2346 0.00822143
R11174 VCC.n2535 VCC.n2534 0.00822143
R11175 VCC.n2565 VCC.n2564 0.00822143
R11176 VCC.n2626 VCC.n2288 0.00822143
R11177 VCC.n2667 VCC.n2284 0.00822143
R11178 VCC.n2668 VCC.n2280 0.00822143
R11179 VCC.n2708 VCC.n2263 0.00822143
R11180 VCC.n2738 VCC.n2235 0.00822143
R11181 VCC.n2769 VCC.n2217 0.00822143
R11182 VCC.n2961 VCC.n2958 0.00822143
R11183 VCC.n3011 VCC.n2943 0.00822143
R11184 VCC.n3051 VCC.n2901 0.00822143
R11185 VCC.n3083 VCC.n2897 0.00822143
R11186 VCC.n3086 VCC.n3085 0.00822143
R11187 VCC.n3117 VCC.n3116 0.00822143
R11188 VCC.n3178 VCC.n2840 0.00822143
R11189 VCC.n3218 VCC.n2836 0.00822143
R11190 VCC.n3219 VCC.n2832 0.00822143
R11191 VCC.n3251 VCC.n2819 0.00822143
R11192 VCC.n3283 VCC.n2783 0.00822143
R11193 VCC.n3324 VCC.n2772 0.00822143
R11194 VCC.n3519 VCC.n3516 0.00822143
R11195 VCC.n3569 VCC.n3501 0.00822143
R11196 VCC.n3609 VCC.n3459 0.00822143
R11197 VCC.n3641 VCC.n3455 0.00822143
R11198 VCC.n3644 VCC.n3643 0.00822143
R11199 VCC.n3674 VCC.n3673 0.00822143
R11200 VCC.n3735 VCC.n3397 0.00822143
R11201 VCC.n3776 VCC.n3393 0.00822143
R11202 VCC.n3777 VCC.n3389 0.00822143
R11203 VCC.n3817 VCC.n3372 0.00822143
R11204 VCC.n3847 VCC.n3344 0.00822143
R11205 VCC.n3878 VCC.n3326 0.00822143
R11206 VCC.n4070 VCC.n4067 0.00822143
R11207 VCC.n4120 VCC.n4052 0.00822143
R11208 VCC.n4160 VCC.n4010 0.00822143
R11209 VCC.n4192 VCC.n4006 0.00822143
R11210 VCC.n4195 VCC.n4194 0.00822143
R11211 VCC.n4226 VCC.n4225 0.00822143
R11212 VCC.n4287 VCC.n3949 0.00822143
R11213 VCC.n4327 VCC.n3945 0.00822143
R11214 VCC.n4328 VCC.n3941 0.00822143
R11215 VCC.n4360 VCC.n3928 0.00822143
R11216 VCC.n4392 VCC.n3892 0.00822143
R11217 VCC.n4433 VCC.n3881 0.00822143
R11218 VCC.n4628 VCC.n4625 0.00822143
R11219 VCC.n4678 VCC.n4610 0.00822143
R11220 VCC.n4718 VCC.n4568 0.00822143
R11221 VCC.n4750 VCC.n4564 0.00822143
R11222 VCC.n4753 VCC.n4752 0.00822143
R11223 VCC.n4783 VCC.n4782 0.00822143
R11224 VCC.n4844 VCC.n4506 0.00822143
R11225 VCC.n4885 VCC.n4502 0.00822143
R11226 VCC.n4886 VCC.n4498 0.00822143
R11227 VCC.n4926 VCC.n4481 0.00822143
R11228 VCC.n4956 VCC.n4453 0.00822143
R11229 VCC.n4987 VCC.n4435 0.00822143
R11230 VCC.n5179 VCC.n5176 0.00822143
R11231 VCC.n5229 VCC.n5161 0.00822143
R11232 VCC.n5269 VCC.n5119 0.00822143
R11233 VCC.n5301 VCC.n5115 0.00822143
R11234 VCC.n5304 VCC.n5303 0.00822143
R11235 VCC.n5335 VCC.n5334 0.00822143
R11236 VCC.n5396 VCC.n5058 0.00822143
R11237 VCC.n5436 VCC.n5054 0.00822143
R11238 VCC.n5437 VCC.n5050 0.00822143
R11239 VCC.n5469 VCC.n5037 0.00822143
R11240 VCC.n5501 VCC.n5001 0.00822143
R11241 VCC.n5542 VCC.n4990 0.00822143
R11242 VCC.n5736 VCC.n5733 0.00822143
R11243 VCC.n5786 VCC.n5718 0.00822143
R11244 VCC.n5826 VCC.n5676 0.00822143
R11245 VCC.n5858 VCC.n5672 0.00822143
R11246 VCC.n5861 VCC.n5860 0.00822143
R11247 VCC.n5891 VCC.n5890 0.00822143
R11248 VCC.n5952 VCC.n5614 0.00822143
R11249 VCC.n5993 VCC.n5610 0.00822143
R11250 VCC.n5994 VCC.n5606 0.00822143
R11251 VCC.n6034 VCC.n5589 0.00822143
R11252 VCC.n6064 VCC.n5561 0.00822143
R11253 VCC.n6095 VCC.n5543 0.00822143
R11254 VCC.n6286 VCC.n6283 0.00822143
R11255 VCC.n6336 VCC.n6268 0.00822143
R11256 VCC.n6376 VCC.n6226 0.00822143
R11257 VCC.n6408 VCC.n6222 0.00822143
R11258 VCC.n6411 VCC.n6410 0.00822143
R11259 VCC.n6442 VCC.n6441 0.00822143
R11260 VCC.n6503 VCC.n6165 0.00822143
R11261 VCC.n6543 VCC.n6161 0.00822143
R11262 VCC.n6544 VCC.n6157 0.00822143
R11263 VCC.n6576 VCC.n6144 0.00822143
R11264 VCC.n6608 VCC.n6108 0.00822143
R11265 VCC.n6649 VCC.n6097 0.00822143
R11266 VCC.n6843 VCC.n6840 0.00822143
R11267 VCC.n6893 VCC.n6825 0.00822143
R11268 VCC.n6933 VCC.n6783 0.00822143
R11269 VCC.n6965 VCC.n6779 0.00822143
R11270 VCC.n6968 VCC.n6967 0.00822143
R11271 VCC.n6998 VCC.n6997 0.00822143
R11272 VCC.n7059 VCC.n6721 0.00822143
R11273 VCC.n7100 VCC.n6717 0.00822143
R11274 VCC.n7101 VCC.n6713 0.00822143
R11275 VCC.n7141 VCC.n6696 0.00822143
R11276 VCC.n7171 VCC.n6668 0.00822143
R11277 VCC.n7202 VCC.n6650 0.00822143
R11278 VCC.n7393 VCC.n7390 0.00822143
R11279 VCC.n7443 VCC.n7375 0.00822143
R11280 VCC.n7483 VCC.n7333 0.00822143
R11281 VCC.n7515 VCC.n7329 0.00822143
R11282 VCC.n7518 VCC.n7517 0.00822143
R11283 VCC.n7549 VCC.n7548 0.00822143
R11284 VCC.n7610 VCC.n7272 0.00822143
R11285 VCC.n7650 VCC.n7268 0.00822143
R11286 VCC.n7651 VCC.n7264 0.00822143
R11287 VCC.n7683 VCC.n7251 0.00822143
R11288 VCC.n7715 VCC.n7215 0.00822143
R11289 VCC.n7756 VCC.n7204 0.00822143
R11290 VCC.n7950 VCC.n7947 0.00822143
R11291 VCC.n8000 VCC.n7932 0.00822143
R11292 VCC.n8040 VCC.n7890 0.00822143
R11293 VCC.n8072 VCC.n7886 0.00822143
R11294 VCC.n8075 VCC.n8074 0.00822143
R11295 VCC.n8105 VCC.n8104 0.00822143
R11296 VCC.n8166 VCC.n7828 0.00822143
R11297 VCC.n8207 VCC.n7824 0.00822143
R11298 VCC.n8208 VCC.n7820 0.00822143
R11299 VCC.n8248 VCC.n7803 0.00822143
R11300 VCC.n8278 VCC.n7775 0.00822143
R11301 VCC.n8309 VCC.n7757 0.00822143
R11302 VCC.n8438 VCC.n8437 0.00822143
R11303 VCC.n8469 VCC.n8468 0.00822143
R11304 VCC.n8530 VCC.n8379 0.00822143
R11305 VCC.n8570 VCC.n8375 0.00822143
R11306 VCC.n8571 VCC.n8371 0.00822143
R11307 VCC.n8603 VCC.n8358 0.00822143
R11308 VCC.n8635 VCC.n8322 0.00822143
R11309 VCC.n8676 VCC.n8311 0.00822143
R11310 VCC.n221 VCC.n176 0.00764286
R11311 VCC.n236 VCC.n235 0.00764286
R11312 VCC.n276 VCC.n274 0.00764286
R11313 VCC.n273 VCC.n145 0.00764286
R11314 VCC.n284 VCC.n134 0.00764286
R11315 VCC.n192 VCC.n189 0.00764286
R11316 VCC.n234 VCC.n175 0.00764286
R11317 VCC.n244 VCC.n172 0.00764286
R11318 VCC.n260 VCC.n164 0.00764286
R11319 VCC.n279 VCC.n148 0.00764286
R11320 VCC.n275 VCC.n146 0.00764286
R11321 VCC.n117 VCC.n111 0.00764286
R11322 VCC.n404 VCC.n403 0.00764286
R11323 VCC.n400 VCC.n85 0.00764286
R11324 VCC.n411 VCC.n73 0.00764286
R11325 VCC.n354 VCC.n353 0.00764286
R11326 VCC.n368 VCC.n103 0.00764286
R11327 VCC.n369 VCC.n100 0.00764286
R11328 VCC.n374 VCC.n373 0.00764286
R11329 VCC.n402 VCC.n89 0.00764286
R11330 VCC.n447 VCC.n67 0.00764286
R11331 VCC.n477 VCC.n53 0.00764286
R11332 VCC.n516 VCC.n27 0.00764286
R11333 VCC.n450 VCC.n63 0.00764286
R11334 VCC.n480 VCC.n479 0.00764286
R11335 VCC.n487 VCC.n46 0.00764286
R11336 VCC.n483 VCC.n482 0.00764286
R11337 VCC.n506 VCC.n34 0.00764286
R11338 VCC.n520 VCC.n28 0.00764286
R11339 VCC.n773 VCC.n728 0.00764286
R11340 VCC.n788 VCC.n787 0.00764286
R11341 VCC.n828 VCC.n826 0.00764286
R11342 VCC.n825 VCC.n697 0.00764286
R11343 VCC.n836 VCC.n686 0.00764286
R11344 VCC.n744 VCC.n741 0.00764286
R11345 VCC.n786 VCC.n727 0.00764286
R11346 VCC.n796 VCC.n724 0.00764286
R11347 VCC.n812 VCC.n716 0.00764286
R11348 VCC.n831 VCC.n700 0.00764286
R11349 VCC.n827 VCC.n698 0.00764286
R11350 VCC.n669 VCC.n663 0.00764286
R11351 VCC.n956 VCC.n955 0.00764286
R11352 VCC.n952 VCC.n637 0.00764286
R11353 VCC.n963 VCC.n625 0.00764286
R11354 VCC.n906 VCC.n905 0.00764286
R11355 VCC.n920 VCC.n655 0.00764286
R11356 VCC.n921 VCC.n652 0.00764286
R11357 VCC.n926 VCC.n925 0.00764286
R11358 VCC.n954 VCC.n641 0.00764286
R11359 VCC.n999 VCC.n619 0.00764286
R11360 VCC.n1029 VCC.n605 0.00764286
R11361 VCC.n1068 VCC.n579 0.00764286
R11362 VCC.n1002 VCC.n615 0.00764286
R11363 VCC.n1032 VCC.n1031 0.00764286
R11364 VCC.n1039 VCC.n598 0.00764286
R11365 VCC.n1035 VCC.n1034 0.00764286
R11366 VCC.n1058 VCC.n586 0.00764286
R11367 VCC.n1072 VCC.n580 0.00764286
R11368 VCC.n1595 VCC.n1158 0.00764286
R11369 VCC.n1139 VCC.n1138 0.00764286
R11370 VCC.n1560 VCC.n1172 0.00764286
R11371 VCC.n1598 VCC.n1597 0.00764286
R11372 VCC.n1591 VCC.n1590 0.00764286
R11373 VCC.n1602 VCC.n1151 0.00764286
R11374 VCC.n1610 VCC.n1609 0.00764286
R11375 VCC.n1136 VCC.n1132 0.00764286
R11376 VCC.n1226 VCC.n1220 0.00764286
R11377 VCC.n1513 VCC.n1512 0.00764286
R11378 VCC.n1509 VCC.n1194 0.00764286
R11379 VCC.n1520 VCC.n1182 0.00764286
R11380 VCC.n1463 VCC.n1462 0.00764286
R11381 VCC.n1477 VCC.n1212 0.00764286
R11382 VCC.n1478 VCC.n1209 0.00764286
R11383 VCC.n1483 VCC.n1482 0.00764286
R11384 VCC.n1511 VCC.n1198 0.00764286
R11385 VCC.n1557 VCC.n1176 0.00764286
R11386 VCC.n1331 VCC.n1286 0.00764286
R11387 VCC.n1346 VCC.n1345 0.00764286
R11388 VCC.n1386 VCC.n1384 0.00764286
R11389 VCC.n1383 VCC.n1255 0.00764286
R11390 VCC.n1394 VCC.n1244 0.00764286
R11391 VCC.n1302 VCC.n1299 0.00764286
R11392 VCC.n1344 VCC.n1285 0.00764286
R11393 VCC.n1354 VCC.n1282 0.00764286
R11394 VCC.n1370 VCC.n1274 0.00764286
R11395 VCC.n1389 VCC.n1258 0.00764286
R11396 VCC.n1385 VCC.n1256 0.00764286
R11397 VCC.n1882 VCC.n1837 0.00764286
R11398 VCC.n1897 VCC.n1896 0.00764286
R11399 VCC.n1937 VCC.n1935 0.00764286
R11400 VCC.n1934 VCC.n1806 0.00764286
R11401 VCC.n1945 VCC.n1795 0.00764286
R11402 VCC.n1853 VCC.n1850 0.00764286
R11403 VCC.n1895 VCC.n1836 0.00764286
R11404 VCC.n1905 VCC.n1833 0.00764286
R11405 VCC.n1921 VCC.n1825 0.00764286
R11406 VCC.n1940 VCC.n1809 0.00764286
R11407 VCC.n1936 VCC.n1807 0.00764286
R11408 VCC.n1778 VCC.n1772 0.00764286
R11409 VCC.n2065 VCC.n2064 0.00764286
R11410 VCC.n2061 VCC.n1746 0.00764286
R11411 VCC.n2072 VCC.n1734 0.00764286
R11412 VCC.n2015 VCC.n2014 0.00764286
R11413 VCC.n2029 VCC.n1764 0.00764286
R11414 VCC.n2030 VCC.n1761 0.00764286
R11415 VCC.n2035 VCC.n2034 0.00764286
R11416 VCC.n2063 VCC.n1750 0.00764286
R11417 VCC.n2108 VCC.n1728 0.00764286
R11418 VCC.n2138 VCC.n1714 0.00764286
R11419 VCC.n2177 VCC.n1688 0.00764286
R11420 VCC.n2111 VCC.n1724 0.00764286
R11421 VCC.n2141 VCC.n2140 0.00764286
R11422 VCC.n2148 VCC.n1707 0.00764286
R11423 VCC.n2144 VCC.n2143 0.00764286
R11424 VCC.n2167 VCC.n1695 0.00764286
R11425 VCC.n2181 VCC.n1689 0.00764286
R11426 VCC.n2704 VCC.n2267 0.00764286
R11427 VCC.n2248 VCC.n2247 0.00764286
R11428 VCC.n2669 VCC.n2281 0.00764286
R11429 VCC.n2707 VCC.n2706 0.00764286
R11430 VCC.n2700 VCC.n2699 0.00764286
R11431 VCC.n2711 VCC.n2260 0.00764286
R11432 VCC.n2719 VCC.n2718 0.00764286
R11433 VCC.n2245 VCC.n2241 0.00764286
R11434 VCC.n2335 VCC.n2329 0.00764286
R11435 VCC.n2622 VCC.n2621 0.00764286
R11436 VCC.n2618 VCC.n2303 0.00764286
R11437 VCC.n2629 VCC.n2291 0.00764286
R11438 VCC.n2572 VCC.n2571 0.00764286
R11439 VCC.n2586 VCC.n2321 0.00764286
R11440 VCC.n2587 VCC.n2318 0.00764286
R11441 VCC.n2592 VCC.n2591 0.00764286
R11442 VCC.n2620 VCC.n2307 0.00764286
R11443 VCC.n2666 VCC.n2285 0.00764286
R11444 VCC.n2440 VCC.n2395 0.00764286
R11445 VCC.n2455 VCC.n2454 0.00764286
R11446 VCC.n2495 VCC.n2493 0.00764286
R11447 VCC.n2492 VCC.n2364 0.00764286
R11448 VCC.n2503 VCC.n2353 0.00764286
R11449 VCC.n2411 VCC.n2408 0.00764286
R11450 VCC.n2453 VCC.n2394 0.00764286
R11451 VCC.n2463 VCC.n2391 0.00764286
R11452 VCC.n2479 VCC.n2383 0.00764286
R11453 VCC.n2498 VCC.n2367 0.00764286
R11454 VCC.n2494 VCC.n2365 0.00764286
R11455 VCC.n2991 VCC.n2946 0.00764286
R11456 VCC.n3006 VCC.n3005 0.00764286
R11457 VCC.n3046 VCC.n3044 0.00764286
R11458 VCC.n3043 VCC.n2915 0.00764286
R11459 VCC.n3054 VCC.n2904 0.00764286
R11460 VCC.n2962 VCC.n2959 0.00764286
R11461 VCC.n3004 VCC.n2945 0.00764286
R11462 VCC.n3014 VCC.n2942 0.00764286
R11463 VCC.n3030 VCC.n2934 0.00764286
R11464 VCC.n3049 VCC.n2918 0.00764286
R11465 VCC.n3045 VCC.n2916 0.00764286
R11466 VCC.n2887 VCC.n2881 0.00764286
R11467 VCC.n3174 VCC.n3173 0.00764286
R11468 VCC.n3170 VCC.n2855 0.00764286
R11469 VCC.n3181 VCC.n2843 0.00764286
R11470 VCC.n3124 VCC.n3123 0.00764286
R11471 VCC.n3138 VCC.n2873 0.00764286
R11472 VCC.n3139 VCC.n2870 0.00764286
R11473 VCC.n3144 VCC.n3143 0.00764286
R11474 VCC.n3172 VCC.n2859 0.00764286
R11475 VCC.n3217 VCC.n2837 0.00764286
R11476 VCC.n3247 VCC.n2823 0.00764286
R11477 VCC.n3286 VCC.n2797 0.00764286
R11478 VCC.n3220 VCC.n2833 0.00764286
R11479 VCC.n3250 VCC.n3249 0.00764286
R11480 VCC.n3257 VCC.n2816 0.00764286
R11481 VCC.n3253 VCC.n3252 0.00764286
R11482 VCC.n3276 VCC.n2804 0.00764286
R11483 VCC.n3290 VCC.n2798 0.00764286
R11484 VCC.n3813 VCC.n3376 0.00764286
R11485 VCC.n3357 VCC.n3356 0.00764286
R11486 VCC.n3778 VCC.n3390 0.00764286
R11487 VCC.n3816 VCC.n3815 0.00764286
R11488 VCC.n3809 VCC.n3808 0.00764286
R11489 VCC.n3820 VCC.n3369 0.00764286
R11490 VCC.n3828 VCC.n3827 0.00764286
R11491 VCC.n3354 VCC.n3350 0.00764286
R11492 VCC.n3444 VCC.n3438 0.00764286
R11493 VCC.n3731 VCC.n3730 0.00764286
R11494 VCC.n3727 VCC.n3412 0.00764286
R11495 VCC.n3738 VCC.n3400 0.00764286
R11496 VCC.n3681 VCC.n3680 0.00764286
R11497 VCC.n3695 VCC.n3430 0.00764286
R11498 VCC.n3696 VCC.n3427 0.00764286
R11499 VCC.n3701 VCC.n3700 0.00764286
R11500 VCC.n3729 VCC.n3416 0.00764286
R11501 VCC.n3775 VCC.n3394 0.00764286
R11502 VCC.n3549 VCC.n3504 0.00764286
R11503 VCC.n3564 VCC.n3563 0.00764286
R11504 VCC.n3604 VCC.n3602 0.00764286
R11505 VCC.n3601 VCC.n3473 0.00764286
R11506 VCC.n3612 VCC.n3462 0.00764286
R11507 VCC.n3520 VCC.n3517 0.00764286
R11508 VCC.n3562 VCC.n3503 0.00764286
R11509 VCC.n3572 VCC.n3500 0.00764286
R11510 VCC.n3588 VCC.n3492 0.00764286
R11511 VCC.n3607 VCC.n3476 0.00764286
R11512 VCC.n3603 VCC.n3474 0.00764286
R11513 VCC.n4100 VCC.n4055 0.00764286
R11514 VCC.n4115 VCC.n4114 0.00764286
R11515 VCC.n4155 VCC.n4153 0.00764286
R11516 VCC.n4152 VCC.n4024 0.00764286
R11517 VCC.n4163 VCC.n4013 0.00764286
R11518 VCC.n4071 VCC.n4068 0.00764286
R11519 VCC.n4113 VCC.n4054 0.00764286
R11520 VCC.n4123 VCC.n4051 0.00764286
R11521 VCC.n4139 VCC.n4043 0.00764286
R11522 VCC.n4158 VCC.n4027 0.00764286
R11523 VCC.n4154 VCC.n4025 0.00764286
R11524 VCC.n3996 VCC.n3990 0.00764286
R11525 VCC.n4283 VCC.n4282 0.00764286
R11526 VCC.n4279 VCC.n3964 0.00764286
R11527 VCC.n4290 VCC.n3952 0.00764286
R11528 VCC.n4233 VCC.n4232 0.00764286
R11529 VCC.n4247 VCC.n3982 0.00764286
R11530 VCC.n4248 VCC.n3979 0.00764286
R11531 VCC.n4253 VCC.n4252 0.00764286
R11532 VCC.n4281 VCC.n3968 0.00764286
R11533 VCC.n4326 VCC.n3946 0.00764286
R11534 VCC.n4356 VCC.n3932 0.00764286
R11535 VCC.n4395 VCC.n3906 0.00764286
R11536 VCC.n4329 VCC.n3942 0.00764286
R11537 VCC.n4359 VCC.n4358 0.00764286
R11538 VCC.n4366 VCC.n3925 0.00764286
R11539 VCC.n4362 VCC.n4361 0.00764286
R11540 VCC.n4385 VCC.n3913 0.00764286
R11541 VCC.n4399 VCC.n3907 0.00764286
R11542 VCC.n4922 VCC.n4485 0.00764286
R11543 VCC.n4466 VCC.n4465 0.00764286
R11544 VCC.n4887 VCC.n4499 0.00764286
R11545 VCC.n4925 VCC.n4924 0.00764286
R11546 VCC.n4918 VCC.n4917 0.00764286
R11547 VCC.n4929 VCC.n4478 0.00764286
R11548 VCC.n4937 VCC.n4936 0.00764286
R11549 VCC.n4463 VCC.n4459 0.00764286
R11550 VCC.n4553 VCC.n4547 0.00764286
R11551 VCC.n4840 VCC.n4839 0.00764286
R11552 VCC.n4836 VCC.n4521 0.00764286
R11553 VCC.n4847 VCC.n4509 0.00764286
R11554 VCC.n4790 VCC.n4789 0.00764286
R11555 VCC.n4804 VCC.n4539 0.00764286
R11556 VCC.n4805 VCC.n4536 0.00764286
R11557 VCC.n4810 VCC.n4809 0.00764286
R11558 VCC.n4838 VCC.n4525 0.00764286
R11559 VCC.n4884 VCC.n4503 0.00764286
R11560 VCC.n4658 VCC.n4613 0.00764286
R11561 VCC.n4673 VCC.n4672 0.00764286
R11562 VCC.n4713 VCC.n4711 0.00764286
R11563 VCC.n4710 VCC.n4582 0.00764286
R11564 VCC.n4721 VCC.n4571 0.00764286
R11565 VCC.n4629 VCC.n4626 0.00764286
R11566 VCC.n4671 VCC.n4612 0.00764286
R11567 VCC.n4681 VCC.n4609 0.00764286
R11568 VCC.n4697 VCC.n4601 0.00764286
R11569 VCC.n4716 VCC.n4585 0.00764286
R11570 VCC.n4712 VCC.n4583 0.00764286
R11571 VCC.n5209 VCC.n5164 0.00764286
R11572 VCC.n5224 VCC.n5223 0.00764286
R11573 VCC.n5264 VCC.n5262 0.00764286
R11574 VCC.n5261 VCC.n5133 0.00764286
R11575 VCC.n5272 VCC.n5122 0.00764286
R11576 VCC.n5180 VCC.n5177 0.00764286
R11577 VCC.n5222 VCC.n5163 0.00764286
R11578 VCC.n5232 VCC.n5160 0.00764286
R11579 VCC.n5248 VCC.n5152 0.00764286
R11580 VCC.n5267 VCC.n5136 0.00764286
R11581 VCC.n5263 VCC.n5134 0.00764286
R11582 VCC.n5105 VCC.n5099 0.00764286
R11583 VCC.n5392 VCC.n5391 0.00764286
R11584 VCC.n5388 VCC.n5073 0.00764286
R11585 VCC.n5399 VCC.n5061 0.00764286
R11586 VCC.n5342 VCC.n5341 0.00764286
R11587 VCC.n5356 VCC.n5091 0.00764286
R11588 VCC.n5357 VCC.n5088 0.00764286
R11589 VCC.n5362 VCC.n5361 0.00764286
R11590 VCC.n5390 VCC.n5077 0.00764286
R11591 VCC.n5435 VCC.n5055 0.00764286
R11592 VCC.n5465 VCC.n5041 0.00764286
R11593 VCC.n5504 VCC.n5015 0.00764286
R11594 VCC.n5438 VCC.n5051 0.00764286
R11595 VCC.n5468 VCC.n5467 0.00764286
R11596 VCC.n5475 VCC.n5034 0.00764286
R11597 VCC.n5471 VCC.n5470 0.00764286
R11598 VCC.n5494 VCC.n5022 0.00764286
R11599 VCC.n5508 VCC.n5016 0.00764286
R11600 VCC.n6030 VCC.n5593 0.00764286
R11601 VCC.n5574 VCC.n5573 0.00764286
R11602 VCC.n5995 VCC.n5607 0.00764286
R11603 VCC.n6033 VCC.n6032 0.00764286
R11604 VCC.n6026 VCC.n6025 0.00764286
R11605 VCC.n6037 VCC.n5586 0.00764286
R11606 VCC.n6045 VCC.n6044 0.00764286
R11607 VCC.n5571 VCC.n5567 0.00764286
R11608 VCC.n5661 VCC.n5655 0.00764286
R11609 VCC.n5948 VCC.n5947 0.00764286
R11610 VCC.n5944 VCC.n5629 0.00764286
R11611 VCC.n5955 VCC.n5617 0.00764286
R11612 VCC.n5898 VCC.n5897 0.00764286
R11613 VCC.n5912 VCC.n5647 0.00764286
R11614 VCC.n5913 VCC.n5644 0.00764286
R11615 VCC.n5918 VCC.n5917 0.00764286
R11616 VCC.n5946 VCC.n5633 0.00764286
R11617 VCC.n5992 VCC.n5611 0.00764286
R11618 VCC.n5766 VCC.n5721 0.00764286
R11619 VCC.n5781 VCC.n5780 0.00764286
R11620 VCC.n5821 VCC.n5819 0.00764286
R11621 VCC.n5818 VCC.n5690 0.00764286
R11622 VCC.n5829 VCC.n5679 0.00764286
R11623 VCC.n5737 VCC.n5734 0.00764286
R11624 VCC.n5779 VCC.n5720 0.00764286
R11625 VCC.n5789 VCC.n5717 0.00764286
R11626 VCC.n5805 VCC.n5709 0.00764286
R11627 VCC.n5824 VCC.n5693 0.00764286
R11628 VCC.n5820 VCC.n5691 0.00764286
R11629 VCC.n6316 VCC.n6271 0.00764286
R11630 VCC.n6331 VCC.n6330 0.00764286
R11631 VCC.n6371 VCC.n6369 0.00764286
R11632 VCC.n6368 VCC.n6240 0.00764286
R11633 VCC.n6379 VCC.n6229 0.00764286
R11634 VCC.n6287 VCC.n6284 0.00764286
R11635 VCC.n6329 VCC.n6270 0.00764286
R11636 VCC.n6339 VCC.n6267 0.00764286
R11637 VCC.n6355 VCC.n6259 0.00764286
R11638 VCC.n6374 VCC.n6243 0.00764286
R11639 VCC.n6370 VCC.n6241 0.00764286
R11640 VCC.n6212 VCC.n6206 0.00764286
R11641 VCC.n6499 VCC.n6498 0.00764286
R11642 VCC.n6495 VCC.n6180 0.00764286
R11643 VCC.n6506 VCC.n6168 0.00764286
R11644 VCC.n6449 VCC.n6448 0.00764286
R11645 VCC.n6463 VCC.n6198 0.00764286
R11646 VCC.n6464 VCC.n6195 0.00764286
R11647 VCC.n6469 VCC.n6468 0.00764286
R11648 VCC.n6497 VCC.n6184 0.00764286
R11649 VCC.n6542 VCC.n6162 0.00764286
R11650 VCC.n6572 VCC.n6148 0.00764286
R11651 VCC.n6611 VCC.n6122 0.00764286
R11652 VCC.n6545 VCC.n6158 0.00764286
R11653 VCC.n6575 VCC.n6574 0.00764286
R11654 VCC.n6582 VCC.n6141 0.00764286
R11655 VCC.n6578 VCC.n6577 0.00764286
R11656 VCC.n6601 VCC.n6129 0.00764286
R11657 VCC.n6615 VCC.n6123 0.00764286
R11658 VCC.n7137 VCC.n6700 0.00764286
R11659 VCC.n6681 VCC.n6680 0.00764286
R11660 VCC.n7102 VCC.n6714 0.00764286
R11661 VCC.n7140 VCC.n7139 0.00764286
R11662 VCC.n7133 VCC.n7132 0.00764286
R11663 VCC.n7144 VCC.n6693 0.00764286
R11664 VCC.n7152 VCC.n7151 0.00764286
R11665 VCC.n6678 VCC.n6674 0.00764286
R11666 VCC.n6768 VCC.n6762 0.00764286
R11667 VCC.n7055 VCC.n7054 0.00764286
R11668 VCC.n7051 VCC.n6736 0.00764286
R11669 VCC.n7062 VCC.n6724 0.00764286
R11670 VCC.n7005 VCC.n7004 0.00764286
R11671 VCC.n7019 VCC.n6754 0.00764286
R11672 VCC.n7020 VCC.n6751 0.00764286
R11673 VCC.n7025 VCC.n7024 0.00764286
R11674 VCC.n7053 VCC.n6740 0.00764286
R11675 VCC.n7099 VCC.n6718 0.00764286
R11676 VCC.n6873 VCC.n6828 0.00764286
R11677 VCC.n6888 VCC.n6887 0.00764286
R11678 VCC.n6928 VCC.n6926 0.00764286
R11679 VCC.n6925 VCC.n6797 0.00764286
R11680 VCC.n6936 VCC.n6786 0.00764286
R11681 VCC.n6844 VCC.n6841 0.00764286
R11682 VCC.n6886 VCC.n6827 0.00764286
R11683 VCC.n6896 VCC.n6824 0.00764286
R11684 VCC.n6912 VCC.n6816 0.00764286
R11685 VCC.n6931 VCC.n6800 0.00764286
R11686 VCC.n6927 VCC.n6798 0.00764286
R11687 VCC.n7423 VCC.n7378 0.00764286
R11688 VCC.n7438 VCC.n7437 0.00764286
R11689 VCC.n7478 VCC.n7476 0.00764286
R11690 VCC.n7475 VCC.n7347 0.00764286
R11691 VCC.n7486 VCC.n7336 0.00764286
R11692 VCC.n7394 VCC.n7391 0.00764286
R11693 VCC.n7436 VCC.n7377 0.00764286
R11694 VCC.n7446 VCC.n7374 0.00764286
R11695 VCC.n7462 VCC.n7366 0.00764286
R11696 VCC.n7481 VCC.n7350 0.00764286
R11697 VCC.n7477 VCC.n7348 0.00764286
R11698 VCC.n7319 VCC.n7313 0.00764286
R11699 VCC.n7606 VCC.n7605 0.00764286
R11700 VCC.n7602 VCC.n7287 0.00764286
R11701 VCC.n7613 VCC.n7275 0.00764286
R11702 VCC.n7556 VCC.n7555 0.00764286
R11703 VCC.n7570 VCC.n7305 0.00764286
R11704 VCC.n7571 VCC.n7302 0.00764286
R11705 VCC.n7576 VCC.n7575 0.00764286
R11706 VCC.n7604 VCC.n7291 0.00764286
R11707 VCC.n7649 VCC.n7269 0.00764286
R11708 VCC.n7679 VCC.n7255 0.00764286
R11709 VCC.n7718 VCC.n7229 0.00764286
R11710 VCC.n7652 VCC.n7265 0.00764286
R11711 VCC.n7682 VCC.n7681 0.00764286
R11712 VCC.n7689 VCC.n7248 0.00764286
R11713 VCC.n7685 VCC.n7684 0.00764286
R11714 VCC.n7708 VCC.n7236 0.00764286
R11715 VCC.n7722 VCC.n7230 0.00764286
R11716 VCC.n8244 VCC.n7807 0.00764286
R11717 VCC.n7788 VCC.n7787 0.00764286
R11718 VCC.n8209 VCC.n7821 0.00764286
R11719 VCC.n8247 VCC.n8246 0.00764286
R11720 VCC.n8240 VCC.n8239 0.00764286
R11721 VCC.n8251 VCC.n7800 0.00764286
R11722 VCC.n8259 VCC.n8258 0.00764286
R11723 VCC.n7785 VCC.n7781 0.00764286
R11724 VCC.n7875 VCC.n7869 0.00764286
R11725 VCC.n8162 VCC.n8161 0.00764286
R11726 VCC.n8158 VCC.n7843 0.00764286
R11727 VCC.n8169 VCC.n7831 0.00764286
R11728 VCC.n8112 VCC.n8111 0.00764286
R11729 VCC.n8126 VCC.n7861 0.00764286
R11730 VCC.n8127 VCC.n7858 0.00764286
R11731 VCC.n8132 VCC.n8131 0.00764286
R11732 VCC.n8160 VCC.n7847 0.00764286
R11733 VCC.n8206 VCC.n7825 0.00764286
R11734 VCC.n7980 VCC.n7935 0.00764286
R11735 VCC.n7995 VCC.n7994 0.00764286
R11736 VCC.n8035 VCC.n8033 0.00764286
R11737 VCC.n8032 VCC.n7904 0.00764286
R11738 VCC.n8043 VCC.n7893 0.00764286
R11739 VCC.n7951 VCC.n7948 0.00764286
R11740 VCC.n7993 VCC.n7934 0.00764286
R11741 VCC.n8003 VCC.n7931 0.00764286
R11742 VCC.n8019 VCC.n7923 0.00764286
R11743 VCC.n8038 VCC.n7907 0.00764286
R11744 VCC.n8034 VCC.n7905 0.00764286
R11745 VCC.n8426 VCC.n8420 0.00764286
R11746 VCC.n8526 VCC.n8525 0.00764286
R11747 VCC.n8522 VCC.n8394 0.00764286
R11748 VCC.n8533 VCC.n8382 0.00764286
R11749 VCC.n8476 VCC.n8475 0.00764286
R11750 VCC.n8490 VCC.n8412 0.00764286
R11751 VCC.n8491 VCC.n8409 0.00764286
R11752 VCC.n8496 VCC.n8495 0.00764286
R11753 VCC.n8524 VCC.n8398 0.00764286
R11754 VCC.n8569 VCC.n8376 0.00764286
R11755 VCC.n8599 VCC.n8362 0.00764286
R11756 VCC.n8638 VCC.n8336 0.00764286
R11757 VCC.n8572 VCC.n8372 0.00764286
R11758 VCC.n8602 VCC.n8601 0.00764286
R11759 VCC.n8609 VCC.n8355 0.00764286
R11760 VCC.n8605 VCC.n8604 0.00764286
R11761 VCC.n8628 VCC.n8343 0.00764286
R11762 VCC.n8642 VCC.n8337 0.00764286
R11763 VCC.n203 VCC.n196 0.00675
R11764 VCC.n246 VCC.n170 0.00675
R11765 VCC.n277 VCC.n276 0.00675
R11766 VCC.n298 VCC.n138 0.00675
R11767 VCC.n239 VCC.n175 0.00675
R11768 VCC.n245 VCC.n171 0.00675
R11769 VCC.n275 VCC.n149 0.00675
R11770 VCC.n283 VCC.n132 0.00675
R11771 VCC.n312 VCC.n128 0.00675
R11772 VCC.n352 VCC.n351 0.00675
R11773 VCC.n367 VCC.n104 0.00675
R11774 VCC.n403 VCC.n401 0.00675
R11775 VCC.n433 VCC.n77 0.00675
R11776 VCC.n314 VCC.n126 0.00675
R11777 VCC.n345 VCC.n113 0.00675
R11778 VCC.n353 VCC.n349 0.00675
R11779 VCC.n406 VCC.n88 0.00675
R11780 VCC.n402 VCC.n86 0.00675
R11781 VCC.n53 VCC.n44 0.00675
R11782 VCC.n47 VCC.n45 0.00675
R11783 VCC.n521 VCC.n27 0.00675
R11784 VCC.n51 VCC.n46 0.00675
R11785 VCC.n486 VCC.n48 0.00675
R11786 VCC.n34 VCC.n31 0.00675
R11787 VCC.n520 VCC.n519 0.00675
R11788 VCC.n518 VCC.n514 0.00675
R11789 VCC.n755 VCC.n748 0.00675
R11790 VCC.n798 VCC.n722 0.00675
R11791 VCC.n829 VCC.n828 0.00675
R11792 VCC.n850 VCC.n690 0.00675
R11793 VCC.n791 VCC.n727 0.00675
R11794 VCC.n797 VCC.n723 0.00675
R11795 VCC.n827 VCC.n701 0.00675
R11796 VCC.n835 VCC.n684 0.00675
R11797 VCC.n864 VCC.n680 0.00675
R11798 VCC.n904 VCC.n903 0.00675
R11799 VCC.n919 VCC.n656 0.00675
R11800 VCC.n955 VCC.n953 0.00675
R11801 VCC.n985 VCC.n629 0.00675
R11802 VCC.n866 VCC.n678 0.00675
R11803 VCC.n897 VCC.n665 0.00675
R11804 VCC.n905 VCC.n901 0.00675
R11805 VCC.n958 VCC.n640 0.00675
R11806 VCC.n954 VCC.n638 0.00675
R11807 VCC.n605 VCC.n596 0.00675
R11808 VCC.n599 VCC.n597 0.00675
R11809 VCC.n1073 VCC.n579 0.00675
R11810 VCC.n603 VCC.n598 0.00675
R11811 VCC.n1038 VCC.n600 0.00675
R11812 VCC.n586 VCC.n583 0.00675
R11813 VCC.n1072 VCC.n1071 0.00675
R11814 VCC.n1070 VCC.n1066 0.00675
R11815 VCC.n1592 VCC.n1158 0.00675
R11816 VCC.n1604 VCC.n1152 0.00675
R11817 VCC.n1138 VCC.n1134 0.00675
R11818 VCC.n1591 VCC.n1156 0.00675
R11819 VCC.n1603 VCC.n1153 0.00675
R11820 VCC.n1609 VCC.n1131 0.00675
R11821 VCC.n1137 VCC.n1136 0.00675
R11822 VCC.n1630 VCC.n1129 0.00675
R11823 VCC.n1461 VCC.n1460 0.00675
R11824 VCC.n1476 VCC.n1213 0.00675
R11825 VCC.n1512 VCC.n1510 0.00675
R11826 VCC.n1543 VCC.n1186 0.00675
R11827 VCC.n1424 VCC.n1236 0.00675
R11828 VCC.n1454 VCC.n1222 0.00675
R11829 VCC.n1462 VCC.n1458 0.00675
R11830 VCC.n1515 VCC.n1197 0.00675
R11831 VCC.n1511 VCC.n1195 0.00675
R11832 VCC.n1313 VCC.n1306 0.00675
R11833 VCC.n1356 VCC.n1280 0.00675
R11834 VCC.n1387 VCC.n1386 0.00675
R11835 VCC.n1408 VCC.n1248 0.00675
R11836 VCC.n1349 VCC.n1285 0.00675
R11837 VCC.n1355 VCC.n1281 0.00675
R11838 VCC.n1385 VCC.n1259 0.00675
R11839 VCC.n1393 VCC.n1242 0.00675
R11840 VCC.n1422 VCC.n1238 0.00675
R11841 VCC.n1864 VCC.n1857 0.00675
R11842 VCC.n1907 VCC.n1831 0.00675
R11843 VCC.n1938 VCC.n1937 0.00675
R11844 VCC.n1959 VCC.n1799 0.00675
R11845 VCC.n1900 VCC.n1836 0.00675
R11846 VCC.n1906 VCC.n1832 0.00675
R11847 VCC.n1936 VCC.n1810 0.00675
R11848 VCC.n1944 VCC.n1793 0.00675
R11849 VCC.n1973 VCC.n1789 0.00675
R11850 VCC.n2013 VCC.n2012 0.00675
R11851 VCC.n2028 VCC.n1765 0.00675
R11852 VCC.n2064 VCC.n2062 0.00675
R11853 VCC.n2094 VCC.n1738 0.00675
R11854 VCC.n1975 VCC.n1787 0.00675
R11855 VCC.n2006 VCC.n1774 0.00675
R11856 VCC.n2014 VCC.n2010 0.00675
R11857 VCC.n2067 VCC.n1749 0.00675
R11858 VCC.n2063 VCC.n1747 0.00675
R11859 VCC.n1714 VCC.n1705 0.00675
R11860 VCC.n1708 VCC.n1706 0.00675
R11861 VCC.n2182 VCC.n1688 0.00675
R11862 VCC.n1712 VCC.n1707 0.00675
R11863 VCC.n2147 VCC.n1709 0.00675
R11864 VCC.n1695 VCC.n1692 0.00675
R11865 VCC.n2181 VCC.n2180 0.00675
R11866 VCC.n2179 VCC.n2175 0.00675
R11867 VCC.n2701 VCC.n2267 0.00675
R11868 VCC.n2713 VCC.n2261 0.00675
R11869 VCC.n2247 VCC.n2243 0.00675
R11870 VCC.n2700 VCC.n2265 0.00675
R11871 VCC.n2712 VCC.n2262 0.00675
R11872 VCC.n2718 VCC.n2240 0.00675
R11873 VCC.n2246 VCC.n2245 0.00675
R11874 VCC.n2739 VCC.n2238 0.00675
R11875 VCC.n2570 VCC.n2569 0.00675
R11876 VCC.n2585 VCC.n2322 0.00675
R11877 VCC.n2621 VCC.n2619 0.00675
R11878 VCC.n2652 VCC.n2295 0.00675
R11879 VCC.n2533 VCC.n2345 0.00675
R11880 VCC.n2563 VCC.n2331 0.00675
R11881 VCC.n2571 VCC.n2567 0.00675
R11882 VCC.n2624 VCC.n2306 0.00675
R11883 VCC.n2620 VCC.n2304 0.00675
R11884 VCC.n2422 VCC.n2415 0.00675
R11885 VCC.n2465 VCC.n2389 0.00675
R11886 VCC.n2496 VCC.n2495 0.00675
R11887 VCC.n2517 VCC.n2357 0.00675
R11888 VCC.n2458 VCC.n2394 0.00675
R11889 VCC.n2464 VCC.n2390 0.00675
R11890 VCC.n2494 VCC.n2368 0.00675
R11891 VCC.n2502 VCC.n2351 0.00675
R11892 VCC.n2531 VCC.n2347 0.00675
R11893 VCC.n2973 VCC.n2966 0.00675
R11894 VCC.n3016 VCC.n2940 0.00675
R11895 VCC.n3047 VCC.n3046 0.00675
R11896 VCC.n3068 VCC.n2908 0.00675
R11897 VCC.n3009 VCC.n2945 0.00675
R11898 VCC.n3015 VCC.n2941 0.00675
R11899 VCC.n3045 VCC.n2919 0.00675
R11900 VCC.n3053 VCC.n2902 0.00675
R11901 VCC.n3082 VCC.n2898 0.00675
R11902 VCC.n3122 VCC.n3121 0.00675
R11903 VCC.n3137 VCC.n2874 0.00675
R11904 VCC.n3173 VCC.n3171 0.00675
R11905 VCC.n3203 VCC.n2847 0.00675
R11906 VCC.n3084 VCC.n2896 0.00675
R11907 VCC.n3115 VCC.n2883 0.00675
R11908 VCC.n3123 VCC.n3119 0.00675
R11909 VCC.n3176 VCC.n2858 0.00675
R11910 VCC.n3172 VCC.n2856 0.00675
R11911 VCC.n2823 VCC.n2814 0.00675
R11912 VCC.n2817 VCC.n2815 0.00675
R11913 VCC.n3291 VCC.n2797 0.00675
R11914 VCC.n2821 VCC.n2816 0.00675
R11915 VCC.n3256 VCC.n2818 0.00675
R11916 VCC.n2804 VCC.n2801 0.00675
R11917 VCC.n3290 VCC.n3289 0.00675
R11918 VCC.n3288 VCC.n3284 0.00675
R11919 VCC.n3810 VCC.n3376 0.00675
R11920 VCC.n3822 VCC.n3370 0.00675
R11921 VCC.n3356 VCC.n3352 0.00675
R11922 VCC.n3809 VCC.n3374 0.00675
R11923 VCC.n3821 VCC.n3371 0.00675
R11924 VCC.n3827 VCC.n3349 0.00675
R11925 VCC.n3355 VCC.n3354 0.00675
R11926 VCC.n3848 VCC.n3347 0.00675
R11927 VCC.n3679 VCC.n3678 0.00675
R11928 VCC.n3694 VCC.n3431 0.00675
R11929 VCC.n3730 VCC.n3728 0.00675
R11930 VCC.n3761 VCC.n3404 0.00675
R11931 VCC.n3642 VCC.n3454 0.00675
R11932 VCC.n3672 VCC.n3440 0.00675
R11933 VCC.n3680 VCC.n3676 0.00675
R11934 VCC.n3733 VCC.n3415 0.00675
R11935 VCC.n3729 VCC.n3413 0.00675
R11936 VCC.n3531 VCC.n3524 0.00675
R11937 VCC.n3574 VCC.n3498 0.00675
R11938 VCC.n3605 VCC.n3604 0.00675
R11939 VCC.n3626 VCC.n3466 0.00675
R11940 VCC.n3567 VCC.n3503 0.00675
R11941 VCC.n3573 VCC.n3499 0.00675
R11942 VCC.n3603 VCC.n3477 0.00675
R11943 VCC.n3611 VCC.n3460 0.00675
R11944 VCC.n3640 VCC.n3456 0.00675
R11945 VCC.n4082 VCC.n4075 0.00675
R11946 VCC.n4125 VCC.n4049 0.00675
R11947 VCC.n4156 VCC.n4155 0.00675
R11948 VCC.n4177 VCC.n4017 0.00675
R11949 VCC.n4118 VCC.n4054 0.00675
R11950 VCC.n4124 VCC.n4050 0.00675
R11951 VCC.n4154 VCC.n4028 0.00675
R11952 VCC.n4162 VCC.n4011 0.00675
R11953 VCC.n4191 VCC.n4007 0.00675
R11954 VCC.n4231 VCC.n4230 0.00675
R11955 VCC.n4246 VCC.n3983 0.00675
R11956 VCC.n4282 VCC.n4280 0.00675
R11957 VCC.n4312 VCC.n3956 0.00675
R11958 VCC.n4193 VCC.n4005 0.00675
R11959 VCC.n4224 VCC.n3992 0.00675
R11960 VCC.n4232 VCC.n4228 0.00675
R11961 VCC.n4285 VCC.n3967 0.00675
R11962 VCC.n4281 VCC.n3965 0.00675
R11963 VCC.n3932 VCC.n3923 0.00675
R11964 VCC.n3926 VCC.n3924 0.00675
R11965 VCC.n4400 VCC.n3906 0.00675
R11966 VCC.n3930 VCC.n3925 0.00675
R11967 VCC.n4365 VCC.n3927 0.00675
R11968 VCC.n3913 VCC.n3910 0.00675
R11969 VCC.n4399 VCC.n4398 0.00675
R11970 VCC.n4397 VCC.n4393 0.00675
R11971 VCC.n4919 VCC.n4485 0.00675
R11972 VCC.n4931 VCC.n4479 0.00675
R11973 VCC.n4465 VCC.n4461 0.00675
R11974 VCC.n4918 VCC.n4483 0.00675
R11975 VCC.n4930 VCC.n4480 0.00675
R11976 VCC.n4936 VCC.n4458 0.00675
R11977 VCC.n4464 VCC.n4463 0.00675
R11978 VCC.n4957 VCC.n4456 0.00675
R11979 VCC.n4788 VCC.n4787 0.00675
R11980 VCC.n4803 VCC.n4540 0.00675
R11981 VCC.n4839 VCC.n4837 0.00675
R11982 VCC.n4870 VCC.n4513 0.00675
R11983 VCC.n4751 VCC.n4563 0.00675
R11984 VCC.n4781 VCC.n4549 0.00675
R11985 VCC.n4789 VCC.n4785 0.00675
R11986 VCC.n4842 VCC.n4524 0.00675
R11987 VCC.n4838 VCC.n4522 0.00675
R11988 VCC.n4640 VCC.n4633 0.00675
R11989 VCC.n4683 VCC.n4607 0.00675
R11990 VCC.n4714 VCC.n4713 0.00675
R11991 VCC.n4735 VCC.n4575 0.00675
R11992 VCC.n4676 VCC.n4612 0.00675
R11993 VCC.n4682 VCC.n4608 0.00675
R11994 VCC.n4712 VCC.n4586 0.00675
R11995 VCC.n4720 VCC.n4569 0.00675
R11996 VCC.n4749 VCC.n4565 0.00675
R11997 VCC.n5191 VCC.n5184 0.00675
R11998 VCC.n5234 VCC.n5158 0.00675
R11999 VCC.n5265 VCC.n5264 0.00675
R12000 VCC.n5286 VCC.n5126 0.00675
R12001 VCC.n5227 VCC.n5163 0.00675
R12002 VCC.n5233 VCC.n5159 0.00675
R12003 VCC.n5263 VCC.n5137 0.00675
R12004 VCC.n5271 VCC.n5120 0.00675
R12005 VCC.n5300 VCC.n5116 0.00675
R12006 VCC.n5340 VCC.n5339 0.00675
R12007 VCC.n5355 VCC.n5092 0.00675
R12008 VCC.n5391 VCC.n5389 0.00675
R12009 VCC.n5421 VCC.n5065 0.00675
R12010 VCC.n5302 VCC.n5114 0.00675
R12011 VCC.n5333 VCC.n5101 0.00675
R12012 VCC.n5341 VCC.n5337 0.00675
R12013 VCC.n5394 VCC.n5076 0.00675
R12014 VCC.n5390 VCC.n5074 0.00675
R12015 VCC.n5041 VCC.n5032 0.00675
R12016 VCC.n5035 VCC.n5033 0.00675
R12017 VCC.n5509 VCC.n5015 0.00675
R12018 VCC.n5039 VCC.n5034 0.00675
R12019 VCC.n5474 VCC.n5036 0.00675
R12020 VCC.n5022 VCC.n5019 0.00675
R12021 VCC.n5508 VCC.n5507 0.00675
R12022 VCC.n5506 VCC.n5502 0.00675
R12023 VCC.n6027 VCC.n5593 0.00675
R12024 VCC.n6039 VCC.n5587 0.00675
R12025 VCC.n5573 VCC.n5569 0.00675
R12026 VCC.n6026 VCC.n5591 0.00675
R12027 VCC.n6038 VCC.n5588 0.00675
R12028 VCC.n6044 VCC.n5566 0.00675
R12029 VCC.n5572 VCC.n5571 0.00675
R12030 VCC.n6065 VCC.n5564 0.00675
R12031 VCC.n5896 VCC.n5895 0.00675
R12032 VCC.n5911 VCC.n5648 0.00675
R12033 VCC.n5947 VCC.n5945 0.00675
R12034 VCC.n5978 VCC.n5621 0.00675
R12035 VCC.n5859 VCC.n5671 0.00675
R12036 VCC.n5889 VCC.n5657 0.00675
R12037 VCC.n5897 VCC.n5893 0.00675
R12038 VCC.n5950 VCC.n5632 0.00675
R12039 VCC.n5946 VCC.n5630 0.00675
R12040 VCC.n5748 VCC.n5741 0.00675
R12041 VCC.n5791 VCC.n5715 0.00675
R12042 VCC.n5822 VCC.n5821 0.00675
R12043 VCC.n5843 VCC.n5683 0.00675
R12044 VCC.n5784 VCC.n5720 0.00675
R12045 VCC.n5790 VCC.n5716 0.00675
R12046 VCC.n5820 VCC.n5694 0.00675
R12047 VCC.n5828 VCC.n5677 0.00675
R12048 VCC.n5857 VCC.n5673 0.00675
R12049 VCC.n6298 VCC.n6291 0.00675
R12050 VCC.n6341 VCC.n6265 0.00675
R12051 VCC.n6372 VCC.n6371 0.00675
R12052 VCC.n6393 VCC.n6233 0.00675
R12053 VCC.n6334 VCC.n6270 0.00675
R12054 VCC.n6340 VCC.n6266 0.00675
R12055 VCC.n6370 VCC.n6244 0.00675
R12056 VCC.n6378 VCC.n6227 0.00675
R12057 VCC.n6407 VCC.n6223 0.00675
R12058 VCC.n6447 VCC.n6446 0.00675
R12059 VCC.n6462 VCC.n6199 0.00675
R12060 VCC.n6498 VCC.n6496 0.00675
R12061 VCC.n6528 VCC.n6172 0.00675
R12062 VCC.n6409 VCC.n6221 0.00675
R12063 VCC.n6440 VCC.n6208 0.00675
R12064 VCC.n6448 VCC.n6444 0.00675
R12065 VCC.n6501 VCC.n6183 0.00675
R12066 VCC.n6497 VCC.n6181 0.00675
R12067 VCC.n6148 VCC.n6139 0.00675
R12068 VCC.n6142 VCC.n6140 0.00675
R12069 VCC.n6616 VCC.n6122 0.00675
R12070 VCC.n6146 VCC.n6141 0.00675
R12071 VCC.n6581 VCC.n6143 0.00675
R12072 VCC.n6129 VCC.n6126 0.00675
R12073 VCC.n6615 VCC.n6614 0.00675
R12074 VCC.n6613 VCC.n6609 0.00675
R12075 VCC.n7134 VCC.n6700 0.00675
R12076 VCC.n7146 VCC.n6694 0.00675
R12077 VCC.n6680 VCC.n6676 0.00675
R12078 VCC.n7133 VCC.n6698 0.00675
R12079 VCC.n7145 VCC.n6695 0.00675
R12080 VCC.n7151 VCC.n6673 0.00675
R12081 VCC.n6679 VCC.n6678 0.00675
R12082 VCC.n7172 VCC.n6671 0.00675
R12083 VCC.n7003 VCC.n7002 0.00675
R12084 VCC.n7018 VCC.n6755 0.00675
R12085 VCC.n7054 VCC.n7052 0.00675
R12086 VCC.n7085 VCC.n6728 0.00675
R12087 VCC.n6966 VCC.n6778 0.00675
R12088 VCC.n6996 VCC.n6764 0.00675
R12089 VCC.n7004 VCC.n7000 0.00675
R12090 VCC.n7057 VCC.n6739 0.00675
R12091 VCC.n7053 VCC.n6737 0.00675
R12092 VCC.n6855 VCC.n6848 0.00675
R12093 VCC.n6898 VCC.n6822 0.00675
R12094 VCC.n6929 VCC.n6928 0.00675
R12095 VCC.n6950 VCC.n6790 0.00675
R12096 VCC.n6891 VCC.n6827 0.00675
R12097 VCC.n6897 VCC.n6823 0.00675
R12098 VCC.n6927 VCC.n6801 0.00675
R12099 VCC.n6935 VCC.n6784 0.00675
R12100 VCC.n6964 VCC.n6780 0.00675
R12101 VCC.n7405 VCC.n7398 0.00675
R12102 VCC.n7448 VCC.n7372 0.00675
R12103 VCC.n7479 VCC.n7478 0.00675
R12104 VCC.n7500 VCC.n7340 0.00675
R12105 VCC.n7441 VCC.n7377 0.00675
R12106 VCC.n7447 VCC.n7373 0.00675
R12107 VCC.n7477 VCC.n7351 0.00675
R12108 VCC.n7485 VCC.n7334 0.00675
R12109 VCC.n7514 VCC.n7330 0.00675
R12110 VCC.n7554 VCC.n7553 0.00675
R12111 VCC.n7569 VCC.n7306 0.00675
R12112 VCC.n7605 VCC.n7603 0.00675
R12113 VCC.n7635 VCC.n7279 0.00675
R12114 VCC.n7516 VCC.n7328 0.00675
R12115 VCC.n7547 VCC.n7315 0.00675
R12116 VCC.n7555 VCC.n7551 0.00675
R12117 VCC.n7608 VCC.n7290 0.00675
R12118 VCC.n7604 VCC.n7288 0.00675
R12119 VCC.n7255 VCC.n7246 0.00675
R12120 VCC.n7249 VCC.n7247 0.00675
R12121 VCC.n7723 VCC.n7229 0.00675
R12122 VCC.n7253 VCC.n7248 0.00675
R12123 VCC.n7688 VCC.n7250 0.00675
R12124 VCC.n7236 VCC.n7233 0.00675
R12125 VCC.n7722 VCC.n7721 0.00675
R12126 VCC.n7720 VCC.n7716 0.00675
R12127 VCC.n8241 VCC.n7807 0.00675
R12128 VCC.n8253 VCC.n7801 0.00675
R12129 VCC.n7787 VCC.n7783 0.00675
R12130 VCC.n8240 VCC.n7805 0.00675
R12131 VCC.n8252 VCC.n7802 0.00675
R12132 VCC.n8258 VCC.n7780 0.00675
R12133 VCC.n7786 VCC.n7785 0.00675
R12134 VCC.n8279 VCC.n7778 0.00675
R12135 VCC.n8110 VCC.n8109 0.00675
R12136 VCC.n8125 VCC.n7862 0.00675
R12137 VCC.n8161 VCC.n8159 0.00675
R12138 VCC.n8192 VCC.n7835 0.00675
R12139 VCC.n8073 VCC.n7885 0.00675
R12140 VCC.n8103 VCC.n7871 0.00675
R12141 VCC.n8111 VCC.n8107 0.00675
R12142 VCC.n8164 VCC.n7846 0.00675
R12143 VCC.n8160 VCC.n7844 0.00675
R12144 VCC.n7962 VCC.n7955 0.00675
R12145 VCC.n8005 VCC.n7929 0.00675
R12146 VCC.n8036 VCC.n8035 0.00675
R12147 VCC.n8057 VCC.n7897 0.00675
R12148 VCC.n7998 VCC.n7934 0.00675
R12149 VCC.n8004 VCC.n7930 0.00675
R12150 VCC.n8034 VCC.n7908 0.00675
R12151 VCC.n8042 VCC.n7891 0.00675
R12152 VCC.n8071 VCC.n7887 0.00675
R12153 VCC.n8474 VCC.n8473 0.00675
R12154 VCC.n8489 VCC.n8413 0.00675
R12155 VCC.n8525 VCC.n8523 0.00675
R12156 VCC.n8555 VCC.n8386 0.00675
R12157 VCC.n8436 VCC.n8435 0.00675
R12158 VCC.n8467 VCC.n8422 0.00675
R12159 VCC.n8475 VCC.n8471 0.00675
R12160 VCC.n8528 VCC.n8397 0.00675
R12161 VCC.n8524 VCC.n8395 0.00675
R12162 VCC.n8362 VCC.n8353 0.00675
R12163 VCC.n8356 VCC.n8354 0.00675
R12164 VCC.n8643 VCC.n8336 0.00675
R12165 VCC.n8360 VCC.n8355 0.00675
R12166 VCC.n8608 VCC.n8357 0.00675
R12167 VCC.n8343 VCC.n8340 0.00675
R12168 VCC.n8642 VCC.n8641 0.00675
R12169 VCC.n8640 VCC.n8636 0.00675
R12170 VCC.n206 VCC.n196 0.00585714
R12171 VCC.n238 VCC.n237 0.00585714
R12172 VCC.n158 VCC.n150 0.00585714
R12173 VCC.n187 VCC.n174 0.00585714
R12174 VCC.n245 VCC.n244 0.00585714
R12175 VCC.n331 VCC.n320 0.00585714
R12176 VCC.n328 VCC.n320 0.00585714
R12177 VCC.n355 VCC.n112 0.00585714
R12178 VCC.n390 VCC.n90 0.00585714
R12179 VCC.n434 VCC.n433 0.00585714
R12180 VCC.n373 VCC.n88 0.00585714
R12181 VCC.n410 VCC.n71 0.00585714
R12182 VCC.n452 VCC.n58 0.00585714
R12183 VCC.n489 VCC.n488 0.00585714
R12184 VCC.n510 VCC.n509 0.00585714
R12185 VCC.n522 VCC.n26 0.00585714
R12186 VCC.n17 VCC.n8 0.00585714
R12187 VCC.n11 VCC.n9 0.00585714
R12188 VCC.n61 VCC.n50 0.00585714
R12189 VCC.n483 VCC.n48 0.00585714
R12190 VCC.n511 VCC.n31 0.00585714
R12191 VCC.n758 VCC.n748 0.00585714
R12192 VCC.n790 VCC.n789 0.00585714
R12193 VCC.n710 VCC.n702 0.00585714
R12194 VCC.n739 VCC.n726 0.00585714
R12195 VCC.n797 VCC.n796 0.00585714
R12196 VCC.n883 VCC.n872 0.00585714
R12197 VCC.n880 VCC.n872 0.00585714
R12198 VCC.n907 VCC.n664 0.00585714
R12199 VCC.n942 VCC.n642 0.00585714
R12200 VCC.n986 VCC.n985 0.00585714
R12201 VCC.n925 VCC.n640 0.00585714
R12202 VCC.n962 VCC.n623 0.00585714
R12203 VCC.n1004 VCC.n610 0.00585714
R12204 VCC.n1041 VCC.n1040 0.00585714
R12205 VCC.n1062 VCC.n1061 0.00585714
R12206 VCC.n1074 VCC.n578 0.00585714
R12207 VCC.n569 VCC.n562 0.00585714
R12208 VCC.n1091 VCC.n563 0.00585714
R12209 VCC.n613 VCC.n602 0.00585714
R12210 VCC.n1035 VCC.n600 0.00585714
R12211 VCC.n1063 VCC.n583 0.00585714
R12212 VCC.n1562 VCC.n1166 0.00585714
R12213 VCC.n1589 VCC.n1588 0.00585714
R12214 VCC.n1626 VCC.n1133 0.00585714
R12215 VCC.n1625 VCC.n1624 0.00585714
R12216 VCC.n1122 VCC.n1119 0.00585714
R12217 VCC.n1641 VCC.n1640 0.00585714
R12218 VCC.n1170 VCC.n1155 0.00585714
R12219 VCC.n1603 VCC.n1602 0.00585714
R12220 VCC.n1627 VCC.n1131 0.00585714
R12221 VCC.n1430 VCC.n1235 0.00585714
R12222 VCC.n1437 VCC.n1430 0.00585714
R12223 VCC.n1464 VCC.n1221 0.00585714
R12224 VCC.n1499 VCC.n1199 0.00585714
R12225 VCC.n1544 VCC.n1543 0.00585714
R12226 VCC.n1482 VCC.n1197 0.00585714
R12227 VCC.n1519 VCC.n1180 0.00585714
R12228 VCC.n1316 VCC.n1306 0.00585714
R12229 VCC.n1348 VCC.n1347 0.00585714
R12230 VCC.n1268 VCC.n1260 0.00585714
R12231 VCC.n1297 VCC.n1284 0.00585714
R12232 VCC.n1355 VCC.n1354 0.00585714
R12233 VCC.n1867 VCC.n1857 0.00585714
R12234 VCC.n1899 VCC.n1898 0.00585714
R12235 VCC.n1819 VCC.n1811 0.00585714
R12236 VCC.n1848 VCC.n1835 0.00585714
R12237 VCC.n1906 VCC.n1905 0.00585714
R12238 VCC.n1992 VCC.n1981 0.00585714
R12239 VCC.n1989 VCC.n1981 0.00585714
R12240 VCC.n2016 VCC.n1773 0.00585714
R12241 VCC.n2051 VCC.n1751 0.00585714
R12242 VCC.n2095 VCC.n2094 0.00585714
R12243 VCC.n2034 VCC.n1749 0.00585714
R12244 VCC.n2071 VCC.n1732 0.00585714
R12245 VCC.n2113 VCC.n1719 0.00585714
R12246 VCC.n2150 VCC.n2149 0.00585714
R12247 VCC.n2171 VCC.n2170 0.00585714
R12248 VCC.n2183 VCC.n1687 0.00585714
R12249 VCC.n1678 VCC.n1671 0.00585714
R12250 VCC.n2200 VCC.n1672 0.00585714
R12251 VCC.n1722 VCC.n1711 0.00585714
R12252 VCC.n2144 VCC.n1709 0.00585714
R12253 VCC.n2172 VCC.n1692 0.00585714
R12254 VCC.n2671 VCC.n2275 0.00585714
R12255 VCC.n2698 VCC.n2697 0.00585714
R12256 VCC.n2735 VCC.n2242 0.00585714
R12257 VCC.n2734 VCC.n2733 0.00585714
R12258 VCC.n2231 VCC.n2228 0.00585714
R12259 VCC.n2750 VCC.n2749 0.00585714
R12260 VCC.n2279 VCC.n2264 0.00585714
R12261 VCC.n2712 VCC.n2711 0.00585714
R12262 VCC.n2736 VCC.n2240 0.00585714
R12263 VCC.n2539 VCC.n2344 0.00585714
R12264 VCC.n2546 VCC.n2539 0.00585714
R12265 VCC.n2573 VCC.n2330 0.00585714
R12266 VCC.n2608 VCC.n2308 0.00585714
R12267 VCC.n2653 VCC.n2652 0.00585714
R12268 VCC.n2591 VCC.n2306 0.00585714
R12269 VCC.n2628 VCC.n2289 0.00585714
R12270 VCC.n2425 VCC.n2415 0.00585714
R12271 VCC.n2457 VCC.n2456 0.00585714
R12272 VCC.n2377 VCC.n2369 0.00585714
R12273 VCC.n2406 VCC.n2393 0.00585714
R12274 VCC.n2464 VCC.n2463 0.00585714
R12275 VCC.n2976 VCC.n2966 0.00585714
R12276 VCC.n3008 VCC.n3007 0.00585714
R12277 VCC.n2928 VCC.n2920 0.00585714
R12278 VCC.n2957 VCC.n2944 0.00585714
R12279 VCC.n3015 VCC.n3014 0.00585714
R12280 VCC.n3101 VCC.n3090 0.00585714
R12281 VCC.n3098 VCC.n3090 0.00585714
R12282 VCC.n3125 VCC.n2882 0.00585714
R12283 VCC.n3160 VCC.n2860 0.00585714
R12284 VCC.n3204 VCC.n3203 0.00585714
R12285 VCC.n3143 VCC.n2858 0.00585714
R12286 VCC.n3180 VCC.n2841 0.00585714
R12287 VCC.n3222 VCC.n2828 0.00585714
R12288 VCC.n3259 VCC.n3258 0.00585714
R12289 VCC.n3280 VCC.n3279 0.00585714
R12290 VCC.n3292 VCC.n2796 0.00585714
R12291 VCC.n2787 VCC.n2780 0.00585714
R12292 VCC.n3309 VCC.n2781 0.00585714
R12293 VCC.n2831 VCC.n2820 0.00585714
R12294 VCC.n3253 VCC.n2818 0.00585714
R12295 VCC.n3281 VCC.n2801 0.00585714
R12296 VCC.n3780 VCC.n3384 0.00585714
R12297 VCC.n3807 VCC.n3806 0.00585714
R12298 VCC.n3844 VCC.n3351 0.00585714
R12299 VCC.n3843 VCC.n3842 0.00585714
R12300 VCC.n3340 VCC.n3337 0.00585714
R12301 VCC.n3859 VCC.n3858 0.00585714
R12302 VCC.n3388 VCC.n3373 0.00585714
R12303 VCC.n3821 VCC.n3820 0.00585714
R12304 VCC.n3845 VCC.n3349 0.00585714
R12305 VCC.n3648 VCC.n3453 0.00585714
R12306 VCC.n3655 VCC.n3648 0.00585714
R12307 VCC.n3682 VCC.n3439 0.00585714
R12308 VCC.n3717 VCC.n3417 0.00585714
R12309 VCC.n3762 VCC.n3761 0.00585714
R12310 VCC.n3700 VCC.n3415 0.00585714
R12311 VCC.n3737 VCC.n3398 0.00585714
R12312 VCC.n3534 VCC.n3524 0.00585714
R12313 VCC.n3566 VCC.n3565 0.00585714
R12314 VCC.n3486 VCC.n3478 0.00585714
R12315 VCC.n3515 VCC.n3502 0.00585714
R12316 VCC.n3573 VCC.n3572 0.00585714
R12317 VCC.n4085 VCC.n4075 0.00585714
R12318 VCC.n4117 VCC.n4116 0.00585714
R12319 VCC.n4037 VCC.n4029 0.00585714
R12320 VCC.n4066 VCC.n4053 0.00585714
R12321 VCC.n4124 VCC.n4123 0.00585714
R12322 VCC.n4210 VCC.n4199 0.00585714
R12323 VCC.n4207 VCC.n4199 0.00585714
R12324 VCC.n4234 VCC.n3991 0.00585714
R12325 VCC.n4269 VCC.n3969 0.00585714
R12326 VCC.n4313 VCC.n4312 0.00585714
R12327 VCC.n4252 VCC.n3967 0.00585714
R12328 VCC.n4289 VCC.n3950 0.00585714
R12329 VCC.n4331 VCC.n3937 0.00585714
R12330 VCC.n4368 VCC.n4367 0.00585714
R12331 VCC.n4389 VCC.n4388 0.00585714
R12332 VCC.n4401 VCC.n3905 0.00585714
R12333 VCC.n3896 VCC.n3889 0.00585714
R12334 VCC.n4418 VCC.n3890 0.00585714
R12335 VCC.n3940 VCC.n3929 0.00585714
R12336 VCC.n4362 VCC.n3927 0.00585714
R12337 VCC.n4390 VCC.n3910 0.00585714
R12338 VCC.n4889 VCC.n4493 0.00585714
R12339 VCC.n4916 VCC.n4915 0.00585714
R12340 VCC.n4953 VCC.n4460 0.00585714
R12341 VCC.n4952 VCC.n4951 0.00585714
R12342 VCC.n4449 VCC.n4446 0.00585714
R12343 VCC.n4968 VCC.n4967 0.00585714
R12344 VCC.n4497 VCC.n4482 0.00585714
R12345 VCC.n4930 VCC.n4929 0.00585714
R12346 VCC.n4954 VCC.n4458 0.00585714
R12347 VCC.n4757 VCC.n4562 0.00585714
R12348 VCC.n4764 VCC.n4757 0.00585714
R12349 VCC.n4791 VCC.n4548 0.00585714
R12350 VCC.n4826 VCC.n4526 0.00585714
R12351 VCC.n4871 VCC.n4870 0.00585714
R12352 VCC.n4809 VCC.n4524 0.00585714
R12353 VCC.n4846 VCC.n4507 0.00585714
R12354 VCC.n4643 VCC.n4633 0.00585714
R12355 VCC.n4675 VCC.n4674 0.00585714
R12356 VCC.n4595 VCC.n4587 0.00585714
R12357 VCC.n4624 VCC.n4611 0.00585714
R12358 VCC.n4682 VCC.n4681 0.00585714
R12359 VCC.n5194 VCC.n5184 0.00585714
R12360 VCC.n5226 VCC.n5225 0.00585714
R12361 VCC.n5146 VCC.n5138 0.00585714
R12362 VCC.n5175 VCC.n5162 0.00585714
R12363 VCC.n5233 VCC.n5232 0.00585714
R12364 VCC.n5319 VCC.n5308 0.00585714
R12365 VCC.n5316 VCC.n5308 0.00585714
R12366 VCC.n5343 VCC.n5100 0.00585714
R12367 VCC.n5378 VCC.n5078 0.00585714
R12368 VCC.n5422 VCC.n5421 0.00585714
R12369 VCC.n5361 VCC.n5076 0.00585714
R12370 VCC.n5398 VCC.n5059 0.00585714
R12371 VCC.n5440 VCC.n5046 0.00585714
R12372 VCC.n5477 VCC.n5476 0.00585714
R12373 VCC.n5498 VCC.n5497 0.00585714
R12374 VCC.n5510 VCC.n5014 0.00585714
R12375 VCC.n5005 VCC.n4998 0.00585714
R12376 VCC.n5527 VCC.n4999 0.00585714
R12377 VCC.n5049 VCC.n5038 0.00585714
R12378 VCC.n5471 VCC.n5036 0.00585714
R12379 VCC.n5499 VCC.n5019 0.00585714
R12380 VCC.n5997 VCC.n5601 0.00585714
R12381 VCC.n6024 VCC.n6023 0.00585714
R12382 VCC.n6061 VCC.n5568 0.00585714
R12383 VCC.n6060 VCC.n6059 0.00585714
R12384 VCC.n5557 VCC.n5554 0.00585714
R12385 VCC.n6076 VCC.n6075 0.00585714
R12386 VCC.n5605 VCC.n5590 0.00585714
R12387 VCC.n6038 VCC.n6037 0.00585714
R12388 VCC.n6062 VCC.n5566 0.00585714
R12389 VCC.n5865 VCC.n5670 0.00585714
R12390 VCC.n5872 VCC.n5865 0.00585714
R12391 VCC.n5899 VCC.n5656 0.00585714
R12392 VCC.n5934 VCC.n5634 0.00585714
R12393 VCC.n5979 VCC.n5978 0.00585714
R12394 VCC.n5917 VCC.n5632 0.00585714
R12395 VCC.n5954 VCC.n5615 0.00585714
R12396 VCC.n5751 VCC.n5741 0.00585714
R12397 VCC.n5783 VCC.n5782 0.00585714
R12398 VCC.n5703 VCC.n5695 0.00585714
R12399 VCC.n5732 VCC.n5719 0.00585714
R12400 VCC.n5790 VCC.n5789 0.00585714
R12401 VCC.n6301 VCC.n6291 0.00585714
R12402 VCC.n6333 VCC.n6332 0.00585714
R12403 VCC.n6253 VCC.n6245 0.00585714
R12404 VCC.n6282 VCC.n6269 0.00585714
R12405 VCC.n6340 VCC.n6339 0.00585714
R12406 VCC.n6426 VCC.n6415 0.00585714
R12407 VCC.n6423 VCC.n6415 0.00585714
R12408 VCC.n6450 VCC.n6207 0.00585714
R12409 VCC.n6485 VCC.n6185 0.00585714
R12410 VCC.n6529 VCC.n6528 0.00585714
R12411 VCC.n6468 VCC.n6183 0.00585714
R12412 VCC.n6505 VCC.n6166 0.00585714
R12413 VCC.n6547 VCC.n6153 0.00585714
R12414 VCC.n6584 VCC.n6583 0.00585714
R12415 VCC.n6605 VCC.n6604 0.00585714
R12416 VCC.n6617 VCC.n6121 0.00585714
R12417 VCC.n6112 VCC.n6105 0.00585714
R12418 VCC.n6634 VCC.n6106 0.00585714
R12419 VCC.n6156 VCC.n6145 0.00585714
R12420 VCC.n6578 VCC.n6143 0.00585714
R12421 VCC.n6606 VCC.n6126 0.00585714
R12422 VCC.n7104 VCC.n6708 0.00585714
R12423 VCC.n7131 VCC.n7130 0.00585714
R12424 VCC.n7168 VCC.n6675 0.00585714
R12425 VCC.n7167 VCC.n7166 0.00585714
R12426 VCC.n6664 VCC.n6661 0.00585714
R12427 VCC.n7183 VCC.n7182 0.00585714
R12428 VCC.n6712 VCC.n6697 0.00585714
R12429 VCC.n7145 VCC.n7144 0.00585714
R12430 VCC.n7169 VCC.n6673 0.00585714
R12431 VCC.n6972 VCC.n6777 0.00585714
R12432 VCC.n6979 VCC.n6972 0.00585714
R12433 VCC.n7006 VCC.n6763 0.00585714
R12434 VCC.n7041 VCC.n6741 0.00585714
R12435 VCC.n7086 VCC.n7085 0.00585714
R12436 VCC.n7024 VCC.n6739 0.00585714
R12437 VCC.n7061 VCC.n6722 0.00585714
R12438 VCC.n6858 VCC.n6848 0.00585714
R12439 VCC.n6890 VCC.n6889 0.00585714
R12440 VCC.n6810 VCC.n6802 0.00585714
R12441 VCC.n6839 VCC.n6826 0.00585714
R12442 VCC.n6897 VCC.n6896 0.00585714
R12443 VCC.n7408 VCC.n7398 0.00585714
R12444 VCC.n7440 VCC.n7439 0.00585714
R12445 VCC.n7360 VCC.n7352 0.00585714
R12446 VCC.n7389 VCC.n7376 0.00585714
R12447 VCC.n7447 VCC.n7446 0.00585714
R12448 VCC.n7533 VCC.n7522 0.00585714
R12449 VCC.n7530 VCC.n7522 0.00585714
R12450 VCC.n7557 VCC.n7314 0.00585714
R12451 VCC.n7592 VCC.n7292 0.00585714
R12452 VCC.n7636 VCC.n7635 0.00585714
R12453 VCC.n7575 VCC.n7290 0.00585714
R12454 VCC.n7612 VCC.n7273 0.00585714
R12455 VCC.n7654 VCC.n7260 0.00585714
R12456 VCC.n7691 VCC.n7690 0.00585714
R12457 VCC.n7712 VCC.n7711 0.00585714
R12458 VCC.n7724 VCC.n7228 0.00585714
R12459 VCC.n7219 VCC.n7212 0.00585714
R12460 VCC.n7741 VCC.n7213 0.00585714
R12461 VCC.n7263 VCC.n7252 0.00585714
R12462 VCC.n7685 VCC.n7250 0.00585714
R12463 VCC.n7713 VCC.n7233 0.00585714
R12464 VCC.n8211 VCC.n7815 0.00585714
R12465 VCC.n8238 VCC.n8237 0.00585714
R12466 VCC.n8275 VCC.n7782 0.00585714
R12467 VCC.n8274 VCC.n8273 0.00585714
R12468 VCC.n7771 VCC.n7768 0.00585714
R12469 VCC.n8290 VCC.n8289 0.00585714
R12470 VCC.n7819 VCC.n7804 0.00585714
R12471 VCC.n8252 VCC.n8251 0.00585714
R12472 VCC.n8276 VCC.n7780 0.00585714
R12473 VCC.n8079 VCC.n7884 0.00585714
R12474 VCC.n8086 VCC.n8079 0.00585714
R12475 VCC.n8113 VCC.n7870 0.00585714
R12476 VCC.n8148 VCC.n7848 0.00585714
R12477 VCC.n8193 VCC.n8192 0.00585714
R12478 VCC.n8131 VCC.n7846 0.00585714
R12479 VCC.n8168 VCC.n7829 0.00585714
R12480 VCC.n7965 VCC.n7955 0.00585714
R12481 VCC.n7997 VCC.n7996 0.00585714
R12482 VCC.n7917 VCC.n7909 0.00585714
R12483 VCC.n7946 VCC.n7933 0.00585714
R12484 VCC.n8004 VCC.n8003 0.00585714
R12485 VCC.n8453 VCC.n8442 0.00585714
R12486 VCC.n8450 VCC.n8442 0.00585714
R12487 VCC.n8477 VCC.n8421 0.00585714
R12488 VCC.n8512 VCC.n8399 0.00585714
R12489 VCC.n8556 VCC.n8555 0.00585714
R12490 VCC.n8495 VCC.n8397 0.00585714
R12491 VCC.n8532 VCC.n8380 0.00585714
R12492 VCC.n8574 VCC.n8367 0.00585714
R12493 VCC.n8611 VCC.n8610 0.00585714
R12494 VCC.n8632 VCC.n8631 0.00585714
R12495 VCC.n8644 VCC.n8335 0.00585714
R12496 VCC.n8326 VCC.n8319 0.00585714
R12497 VCC.n8661 VCC.n8320 0.00585714
R12498 VCC.n8370 VCC.n8359 0.00585714
R12499 VCC.n8605 VCC.n8357 0.00585714
R12500 VCC.n8633 VCC.n8340 0.00585714
R12501 VCC.n299 VCC.n137 0.00496429
R12502 VCC.n299 VCC.n298 0.00496429
R12503 VCC.n216 VCC.n189 0.00496429
R12504 VCC.n219 VCC.n187 0.00496429
R12505 VCC.n164 VCC.n148 0.00496429
R12506 VCC.n306 VCC.n132 0.00496429
R12507 VCC.n309 VCC.n128 0.00496429
R12508 VCC.n328 VCC.n327 0.00496429
R12509 VCC.n318 VCC.n126 0.00496429
R12510 VCC.n345 VCC.n344 0.00496429
R12511 VCC.n369 VCC.n368 0.00496429
R12512 VCC.n441 VCC.n71 0.00496429
R12513 VCC.n444 VCC.n67 0.00496429
R12514 VCC.n459 VCC.n63 0.00496429
R12515 VCC.n464 VCC.n61 0.00496429
R12516 VCC.n29 VCC.n14 0.00496429
R12517 VCC.n535 VCC.n14 0.00496429
R12518 VCC.n538 VCC.n1 0.00496429
R12519 VCC.n851 VCC.n689 0.00496429
R12520 VCC.n851 VCC.n850 0.00496429
R12521 VCC.n768 VCC.n741 0.00496429
R12522 VCC.n771 VCC.n739 0.00496429
R12523 VCC.n716 VCC.n700 0.00496429
R12524 VCC.n858 VCC.n684 0.00496429
R12525 VCC.n861 VCC.n680 0.00496429
R12526 VCC.n880 VCC.n879 0.00496429
R12527 VCC.n870 VCC.n678 0.00496429
R12528 VCC.n897 VCC.n896 0.00496429
R12529 VCC.n921 VCC.n920 0.00496429
R12530 VCC.n993 VCC.n623 0.00496429
R12531 VCC.n996 VCC.n619 0.00496429
R12532 VCC.n1011 VCC.n615 0.00496429
R12533 VCC.n1016 VCC.n613 0.00496429
R12534 VCC.n581 VCC.n566 0.00496429
R12535 VCC.n1087 VCC.n566 0.00496429
R12536 VCC.n1090 VCC.n555 0.00496429
R12537 VCC.n1570 VCC.n1172 0.00496429
R12538 VCC.n1573 VCC.n1170 0.00496429
R12539 VCC.n1631 VCC.n1127 0.00496429
R12540 VCC.n1634 VCC.n1127 0.00496429
R12541 VCC.n1637 VCC.n1109 0.00496429
R12542 VCC.n1437 VCC.n1436 0.00496429
R12543 VCC.n1428 VCC.n1236 0.00496429
R12544 VCC.n1454 VCC.n1453 0.00496429
R12545 VCC.n1478 VCC.n1477 0.00496429
R12546 VCC.n1551 VCC.n1180 0.00496429
R12547 VCC.n1554 VCC.n1176 0.00496429
R12548 VCC.n1409 VCC.n1247 0.00496429
R12549 VCC.n1409 VCC.n1408 0.00496429
R12550 VCC.n1326 VCC.n1299 0.00496429
R12551 VCC.n1329 VCC.n1297 0.00496429
R12552 VCC.n1274 VCC.n1258 0.00496429
R12553 VCC.n1416 VCC.n1242 0.00496429
R12554 VCC.n1419 VCC.n1238 0.00496429
R12555 VCC.n1960 VCC.n1798 0.00496429
R12556 VCC.n1960 VCC.n1959 0.00496429
R12557 VCC.n1877 VCC.n1850 0.00496429
R12558 VCC.n1880 VCC.n1848 0.00496429
R12559 VCC.n1825 VCC.n1809 0.00496429
R12560 VCC.n1967 VCC.n1793 0.00496429
R12561 VCC.n1970 VCC.n1789 0.00496429
R12562 VCC.n1989 VCC.n1988 0.00496429
R12563 VCC.n1979 VCC.n1787 0.00496429
R12564 VCC.n2006 VCC.n2005 0.00496429
R12565 VCC.n2030 VCC.n2029 0.00496429
R12566 VCC.n2102 VCC.n1732 0.00496429
R12567 VCC.n2105 VCC.n1728 0.00496429
R12568 VCC.n2120 VCC.n1724 0.00496429
R12569 VCC.n2125 VCC.n1722 0.00496429
R12570 VCC.n1690 VCC.n1675 0.00496429
R12571 VCC.n2196 VCC.n1675 0.00496429
R12572 VCC.n2199 VCC.n1664 0.00496429
R12573 VCC.n2679 VCC.n2281 0.00496429
R12574 VCC.n2682 VCC.n2279 0.00496429
R12575 VCC.n2740 VCC.n2236 0.00496429
R12576 VCC.n2743 VCC.n2236 0.00496429
R12577 VCC.n2746 VCC.n2218 0.00496429
R12578 VCC.n2546 VCC.n2545 0.00496429
R12579 VCC.n2537 VCC.n2345 0.00496429
R12580 VCC.n2563 VCC.n2562 0.00496429
R12581 VCC.n2587 VCC.n2586 0.00496429
R12582 VCC.n2660 VCC.n2289 0.00496429
R12583 VCC.n2663 VCC.n2285 0.00496429
R12584 VCC.n2518 VCC.n2356 0.00496429
R12585 VCC.n2518 VCC.n2517 0.00496429
R12586 VCC.n2435 VCC.n2408 0.00496429
R12587 VCC.n2438 VCC.n2406 0.00496429
R12588 VCC.n2383 VCC.n2367 0.00496429
R12589 VCC.n2525 VCC.n2351 0.00496429
R12590 VCC.n2528 VCC.n2347 0.00496429
R12591 VCC.n3069 VCC.n2907 0.00496429
R12592 VCC.n3069 VCC.n3068 0.00496429
R12593 VCC.n2986 VCC.n2959 0.00496429
R12594 VCC.n2989 VCC.n2957 0.00496429
R12595 VCC.n2934 VCC.n2918 0.00496429
R12596 VCC.n3076 VCC.n2902 0.00496429
R12597 VCC.n3079 VCC.n2898 0.00496429
R12598 VCC.n3098 VCC.n3097 0.00496429
R12599 VCC.n3088 VCC.n2896 0.00496429
R12600 VCC.n3115 VCC.n3114 0.00496429
R12601 VCC.n3139 VCC.n3138 0.00496429
R12602 VCC.n3211 VCC.n2841 0.00496429
R12603 VCC.n3214 VCC.n2837 0.00496429
R12604 VCC.n3229 VCC.n2833 0.00496429
R12605 VCC.n3234 VCC.n2831 0.00496429
R12606 VCC.n2799 VCC.n2784 0.00496429
R12607 VCC.n3305 VCC.n2784 0.00496429
R12608 VCC.n3308 VCC.n2773 0.00496429
R12609 VCC.n3788 VCC.n3390 0.00496429
R12610 VCC.n3791 VCC.n3388 0.00496429
R12611 VCC.n3849 VCC.n3345 0.00496429
R12612 VCC.n3852 VCC.n3345 0.00496429
R12613 VCC.n3855 VCC.n3327 0.00496429
R12614 VCC.n3655 VCC.n3654 0.00496429
R12615 VCC.n3646 VCC.n3454 0.00496429
R12616 VCC.n3672 VCC.n3671 0.00496429
R12617 VCC.n3696 VCC.n3695 0.00496429
R12618 VCC.n3769 VCC.n3398 0.00496429
R12619 VCC.n3772 VCC.n3394 0.00496429
R12620 VCC.n3627 VCC.n3465 0.00496429
R12621 VCC.n3627 VCC.n3626 0.00496429
R12622 VCC.n3544 VCC.n3517 0.00496429
R12623 VCC.n3547 VCC.n3515 0.00496429
R12624 VCC.n3492 VCC.n3476 0.00496429
R12625 VCC.n3634 VCC.n3460 0.00496429
R12626 VCC.n3637 VCC.n3456 0.00496429
R12627 VCC.n4178 VCC.n4016 0.00496429
R12628 VCC.n4178 VCC.n4177 0.00496429
R12629 VCC.n4095 VCC.n4068 0.00496429
R12630 VCC.n4098 VCC.n4066 0.00496429
R12631 VCC.n4043 VCC.n4027 0.00496429
R12632 VCC.n4185 VCC.n4011 0.00496429
R12633 VCC.n4188 VCC.n4007 0.00496429
R12634 VCC.n4207 VCC.n4206 0.00496429
R12635 VCC.n4197 VCC.n4005 0.00496429
R12636 VCC.n4224 VCC.n4223 0.00496429
R12637 VCC.n4248 VCC.n4247 0.00496429
R12638 VCC.n4320 VCC.n3950 0.00496429
R12639 VCC.n4323 VCC.n3946 0.00496429
R12640 VCC.n4338 VCC.n3942 0.00496429
R12641 VCC.n4343 VCC.n3940 0.00496429
R12642 VCC.n3908 VCC.n3893 0.00496429
R12643 VCC.n4414 VCC.n3893 0.00496429
R12644 VCC.n4417 VCC.n3882 0.00496429
R12645 VCC.n4897 VCC.n4499 0.00496429
R12646 VCC.n4900 VCC.n4497 0.00496429
R12647 VCC.n4958 VCC.n4454 0.00496429
R12648 VCC.n4961 VCC.n4454 0.00496429
R12649 VCC.n4964 VCC.n4436 0.00496429
R12650 VCC.n4764 VCC.n4763 0.00496429
R12651 VCC.n4755 VCC.n4563 0.00496429
R12652 VCC.n4781 VCC.n4780 0.00496429
R12653 VCC.n4805 VCC.n4804 0.00496429
R12654 VCC.n4878 VCC.n4507 0.00496429
R12655 VCC.n4881 VCC.n4503 0.00496429
R12656 VCC.n4736 VCC.n4574 0.00496429
R12657 VCC.n4736 VCC.n4735 0.00496429
R12658 VCC.n4653 VCC.n4626 0.00496429
R12659 VCC.n4656 VCC.n4624 0.00496429
R12660 VCC.n4601 VCC.n4585 0.00496429
R12661 VCC.n4743 VCC.n4569 0.00496429
R12662 VCC.n4746 VCC.n4565 0.00496429
R12663 VCC.n5287 VCC.n5125 0.00496429
R12664 VCC.n5287 VCC.n5286 0.00496429
R12665 VCC.n5204 VCC.n5177 0.00496429
R12666 VCC.n5207 VCC.n5175 0.00496429
R12667 VCC.n5152 VCC.n5136 0.00496429
R12668 VCC.n5294 VCC.n5120 0.00496429
R12669 VCC.n5297 VCC.n5116 0.00496429
R12670 VCC.n5316 VCC.n5315 0.00496429
R12671 VCC.n5306 VCC.n5114 0.00496429
R12672 VCC.n5333 VCC.n5332 0.00496429
R12673 VCC.n5357 VCC.n5356 0.00496429
R12674 VCC.n5429 VCC.n5059 0.00496429
R12675 VCC.n5432 VCC.n5055 0.00496429
R12676 VCC.n5447 VCC.n5051 0.00496429
R12677 VCC.n5452 VCC.n5049 0.00496429
R12678 VCC.n5017 VCC.n5002 0.00496429
R12679 VCC.n5523 VCC.n5002 0.00496429
R12680 VCC.n5526 VCC.n4991 0.00496429
R12681 VCC.n6005 VCC.n5607 0.00496429
R12682 VCC.n6008 VCC.n5605 0.00496429
R12683 VCC.n6066 VCC.n5562 0.00496429
R12684 VCC.n6069 VCC.n5562 0.00496429
R12685 VCC.n6072 VCC.n5544 0.00496429
R12686 VCC.n5872 VCC.n5871 0.00496429
R12687 VCC.n5863 VCC.n5671 0.00496429
R12688 VCC.n5889 VCC.n5888 0.00496429
R12689 VCC.n5913 VCC.n5912 0.00496429
R12690 VCC.n5986 VCC.n5615 0.00496429
R12691 VCC.n5989 VCC.n5611 0.00496429
R12692 VCC.n5844 VCC.n5682 0.00496429
R12693 VCC.n5844 VCC.n5843 0.00496429
R12694 VCC.n5761 VCC.n5734 0.00496429
R12695 VCC.n5764 VCC.n5732 0.00496429
R12696 VCC.n5709 VCC.n5693 0.00496429
R12697 VCC.n5851 VCC.n5677 0.00496429
R12698 VCC.n5854 VCC.n5673 0.00496429
R12699 VCC.n6394 VCC.n6232 0.00496429
R12700 VCC.n6394 VCC.n6393 0.00496429
R12701 VCC.n6311 VCC.n6284 0.00496429
R12702 VCC.n6314 VCC.n6282 0.00496429
R12703 VCC.n6259 VCC.n6243 0.00496429
R12704 VCC.n6401 VCC.n6227 0.00496429
R12705 VCC.n6404 VCC.n6223 0.00496429
R12706 VCC.n6423 VCC.n6422 0.00496429
R12707 VCC.n6413 VCC.n6221 0.00496429
R12708 VCC.n6440 VCC.n6439 0.00496429
R12709 VCC.n6464 VCC.n6463 0.00496429
R12710 VCC.n6536 VCC.n6166 0.00496429
R12711 VCC.n6539 VCC.n6162 0.00496429
R12712 VCC.n6554 VCC.n6158 0.00496429
R12713 VCC.n6559 VCC.n6156 0.00496429
R12714 VCC.n6124 VCC.n6109 0.00496429
R12715 VCC.n6630 VCC.n6109 0.00496429
R12716 VCC.n6633 VCC.n6098 0.00496429
R12717 VCC.n7112 VCC.n6714 0.00496429
R12718 VCC.n7115 VCC.n6712 0.00496429
R12719 VCC.n7173 VCC.n6669 0.00496429
R12720 VCC.n7176 VCC.n6669 0.00496429
R12721 VCC.n7179 VCC.n6651 0.00496429
R12722 VCC.n6979 VCC.n6978 0.00496429
R12723 VCC.n6970 VCC.n6778 0.00496429
R12724 VCC.n6996 VCC.n6995 0.00496429
R12725 VCC.n7020 VCC.n7019 0.00496429
R12726 VCC.n7093 VCC.n6722 0.00496429
R12727 VCC.n7096 VCC.n6718 0.00496429
R12728 VCC.n6951 VCC.n6789 0.00496429
R12729 VCC.n6951 VCC.n6950 0.00496429
R12730 VCC.n6868 VCC.n6841 0.00496429
R12731 VCC.n6871 VCC.n6839 0.00496429
R12732 VCC.n6816 VCC.n6800 0.00496429
R12733 VCC.n6958 VCC.n6784 0.00496429
R12734 VCC.n6961 VCC.n6780 0.00496429
R12735 VCC.n7501 VCC.n7339 0.00496429
R12736 VCC.n7501 VCC.n7500 0.00496429
R12737 VCC.n7418 VCC.n7391 0.00496429
R12738 VCC.n7421 VCC.n7389 0.00496429
R12739 VCC.n7366 VCC.n7350 0.00496429
R12740 VCC.n7508 VCC.n7334 0.00496429
R12741 VCC.n7511 VCC.n7330 0.00496429
R12742 VCC.n7530 VCC.n7529 0.00496429
R12743 VCC.n7520 VCC.n7328 0.00496429
R12744 VCC.n7547 VCC.n7546 0.00496429
R12745 VCC.n7571 VCC.n7570 0.00496429
R12746 VCC.n7643 VCC.n7273 0.00496429
R12747 VCC.n7646 VCC.n7269 0.00496429
R12748 VCC.n7661 VCC.n7265 0.00496429
R12749 VCC.n7666 VCC.n7263 0.00496429
R12750 VCC.n7231 VCC.n7216 0.00496429
R12751 VCC.n7737 VCC.n7216 0.00496429
R12752 VCC.n7740 VCC.n7205 0.00496429
R12753 VCC.n8219 VCC.n7821 0.00496429
R12754 VCC.n8222 VCC.n7819 0.00496429
R12755 VCC.n8280 VCC.n7776 0.00496429
R12756 VCC.n8283 VCC.n7776 0.00496429
R12757 VCC.n8286 VCC.n7758 0.00496429
R12758 VCC.n8086 VCC.n8085 0.00496429
R12759 VCC.n8077 VCC.n7885 0.00496429
R12760 VCC.n8103 VCC.n8102 0.00496429
R12761 VCC.n8127 VCC.n8126 0.00496429
R12762 VCC.n8200 VCC.n7829 0.00496429
R12763 VCC.n8203 VCC.n7825 0.00496429
R12764 VCC.n8058 VCC.n7896 0.00496429
R12765 VCC.n8058 VCC.n8057 0.00496429
R12766 VCC.n7975 VCC.n7948 0.00496429
R12767 VCC.n7978 VCC.n7946 0.00496429
R12768 VCC.n7923 VCC.n7907 0.00496429
R12769 VCC.n8065 VCC.n7891 0.00496429
R12770 VCC.n8068 VCC.n7887 0.00496429
R12771 VCC.n8450 VCC.n8449 0.00496429
R12772 VCC.n8440 VCC.n8435 0.00496429
R12773 VCC.n8467 VCC.n8466 0.00496429
R12774 VCC.n8491 VCC.n8490 0.00496429
R12775 VCC.n8563 VCC.n8380 0.00496429
R12776 VCC.n8566 VCC.n8376 0.00496429
R12777 VCC.n8581 VCC.n8372 0.00496429
R12778 VCC.n8586 VCC.n8370 0.00496429
R12779 VCC.n8338 VCC.n8323 0.00496429
R12780 VCC.n8657 VCC.n8323 0.00496429
R12781 VCC.n8660 VCC.n8312 0.00496429
R12782 VCC.n243 VCC.n242 0.00486429
R12783 VCC.n257 VCC.n165 0.00486429
R12784 VCC.n259 VCC.n258 0.00486429
R12785 VCC.n280 VCC.n147 0.00486429
R12786 VCC.n370 VCC.n102 0.00486429
R12787 VCC.n380 VCC.n371 0.00486429
R12788 VCC.n379 VCC.n372 0.00486429
R12789 VCC.n407 VCC.n87 0.00486429
R12790 VCC.n485 VCC.n484 0.00486429
R12791 VCC.n503 VCC.n35 0.00486429
R12792 VCC.n505 VCC.n504 0.00486429
R12793 VCC.n512 VCC.n30 0.00486429
R12794 VCC.n795 VCC.n794 0.00486429
R12795 VCC.n809 VCC.n717 0.00486429
R12796 VCC.n811 VCC.n810 0.00486429
R12797 VCC.n832 VCC.n699 0.00486429
R12798 VCC.n922 VCC.n654 0.00486429
R12799 VCC.n932 VCC.n923 0.00486429
R12800 VCC.n931 VCC.n924 0.00486429
R12801 VCC.n959 VCC.n639 0.00486429
R12802 VCC.n1037 VCC.n1036 0.00486429
R12803 VCC.n1055 VCC.n587 0.00486429
R12804 VCC.n1057 VCC.n1056 0.00486429
R12805 VCC.n1064 VCC.n582 0.00486429
R12806 VCC.n1353 VCC.n1352 0.00486429
R12807 VCC.n1367 VCC.n1275 0.00486429
R12808 VCC.n1369 VCC.n1368 0.00486429
R12809 VCC.n1390 VCC.n1257 0.00486429
R12810 VCC.n1479 VCC.n1211 0.00486429
R12811 VCC.n1489 VCC.n1480 0.00486429
R12812 VCC.n1488 VCC.n1481 0.00486429
R12813 VCC.n1516 VCC.n1196 0.00486429
R12814 VCC.n1601 VCC.n1600 0.00486429
R12815 VCC.n1608 VCC.n1150 0.00486429
R12816 VCC.n1612 VCC.n1611 0.00486429
R12817 VCC.n1628 VCC.n1130 0.00486429
R12818 VCC.n1904 VCC.n1903 0.00486429
R12819 VCC.n1918 VCC.n1826 0.00486429
R12820 VCC.n1920 VCC.n1919 0.00486429
R12821 VCC.n1941 VCC.n1808 0.00486429
R12822 VCC.n2031 VCC.n1763 0.00486429
R12823 VCC.n2041 VCC.n2032 0.00486429
R12824 VCC.n2040 VCC.n2033 0.00486429
R12825 VCC.n2068 VCC.n1748 0.00486429
R12826 VCC.n2146 VCC.n2145 0.00486429
R12827 VCC.n2164 VCC.n1696 0.00486429
R12828 VCC.n2166 VCC.n2165 0.00486429
R12829 VCC.n2173 VCC.n1691 0.00486429
R12830 VCC.n2462 VCC.n2461 0.00486429
R12831 VCC.n2476 VCC.n2384 0.00486429
R12832 VCC.n2478 VCC.n2477 0.00486429
R12833 VCC.n2499 VCC.n2366 0.00486429
R12834 VCC.n2588 VCC.n2320 0.00486429
R12835 VCC.n2598 VCC.n2589 0.00486429
R12836 VCC.n2597 VCC.n2590 0.00486429
R12837 VCC.n2625 VCC.n2305 0.00486429
R12838 VCC.n2710 VCC.n2709 0.00486429
R12839 VCC.n2717 VCC.n2259 0.00486429
R12840 VCC.n2721 VCC.n2720 0.00486429
R12841 VCC.n2737 VCC.n2239 0.00486429
R12842 VCC.n3013 VCC.n3012 0.00486429
R12843 VCC.n3027 VCC.n2935 0.00486429
R12844 VCC.n3029 VCC.n3028 0.00486429
R12845 VCC.n3050 VCC.n2917 0.00486429
R12846 VCC.n3140 VCC.n2872 0.00486429
R12847 VCC.n3150 VCC.n3141 0.00486429
R12848 VCC.n3149 VCC.n3142 0.00486429
R12849 VCC.n3177 VCC.n2857 0.00486429
R12850 VCC.n3255 VCC.n3254 0.00486429
R12851 VCC.n3273 VCC.n2805 0.00486429
R12852 VCC.n3275 VCC.n3274 0.00486429
R12853 VCC.n3282 VCC.n2800 0.00486429
R12854 VCC.n3571 VCC.n3570 0.00486429
R12855 VCC.n3585 VCC.n3493 0.00486429
R12856 VCC.n3587 VCC.n3586 0.00486429
R12857 VCC.n3608 VCC.n3475 0.00486429
R12858 VCC.n3697 VCC.n3429 0.00486429
R12859 VCC.n3707 VCC.n3698 0.00486429
R12860 VCC.n3706 VCC.n3699 0.00486429
R12861 VCC.n3734 VCC.n3414 0.00486429
R12862 VCC.n3819 VCC.n3818 0.00486429
R12863 VCC.n3826 VCC.n3368 0.00486429
R12864 VCC.n3830 VCC.n3829 0.00486429
R12865 VCC.n3846 VCC.n3348 0.00486429
R12866 VCC.n4122 VCC.n4121 0.00486429
R12867 VCC.n4136 VCC.n4044 0.00486429
R12868 VCC.n4138 VCC.n4137 0.00486429
R12869 VCC.n4159 VCC.n4026 0.00486429
R12870 VCC.n4249 VCC.n3981 0.00486429
R12871 VCC.n4259 VCC.n4250 0.00486429
R12872 VCC.n4258 VCC.n4251 0.00486429
R12873 VCC.n4286 VCC.n3966 0.00486429
R12874 VCC.n4364 VCC.n4363 0.00486429
R12875 VCC.n4382 VCC.n3914 0.00486429
R12876 VCC.n4384 VCC.n4383 0.00486429
R12877 VCC.n4391 VCC.n3909 0.00486429
R12878 VCC.n4680 VCC.n4679 0.00486429
R12879 VCC.n4694 VCC.n4602 0.00486429
R12880 VCC.n4696 VCC.n4695 0.00486429
R12881 VCC.n4717 VCC.n4584 0.00486429
R12882 VCC.n4806 VCC.n4538 0.00486429
R12883 VCC.n4816 VCC.n4807 0.00486429
R12884 VCC.n4815 VCC.n4808 0.00486429
R12885 VCC.n4843 VCC.n4523 0.00486429
R12886 VCC.n4928 VCC.n4927 0.00486429
R12887 VCC.n4935 VCC.n4477 0.00486429
R12888 VCC.n4939 VCC.n4938 0.00486429
R12889 VCC.n4955 VCC.n4457 0.00486429
R12890 VCC.n5231 VCC.n5230 0.00486429
R12891 VCC.n5245 VCC.n5153 0.00486429
R12892 VCC.n5247 VCC.n5246 0.00486429
R12893 VCC.n5268 VCC.n5135 0.00486429
R12894 VCC.n5358 VCC.n5090 0.00486429
R12895 VCC.n5368 VCC.n5359 0.00486429
R12896 VCC.n5367 VCC.n5360 0.00486429
R12897 VCC.n5395 VCC.n5075 0.00486429
R12898 VCC.n5473 VCC.n5472 0.00486429
R12899 VCC.n5491 VCC.n5023 0.00486429
R12900 VCC.n5493 VCC.n5492 0.00486429
R12901 VCC.n5500 VCC.n5018 0.00486429
R12902 VCC.n5788 VCC.n5787 0.00486429
R12903 VCC.n5802 VCC.n5710 0.00486429
R12904 VCC.n5804 VCC.n5803 0.00486429
R12905 VCC.n5825 VCC.n5692 0.00486429
R12906 VCC.n5914 VCC.n5646 0.00486429
R12907 VCC.n5924 VCC.n5915 0.00486429
R12908 VCC.n5923 VCC.n5916 0.00486429
R12909 VCC.n5951 VCC.n5631 0.00486429
R12910 VCC.n6036 VCC.n6035 0.00486429
R12911 VCC.n6043 VCC.n5585 0.00486429
R12912 VCC.n6047 VCC.n6046 0.00486429
R12913 VCC.n6063 VCC.n5565 0.00486429
R12914 VCC.n6338 VCC.n6337 0.00486429
R12915 VCC.n6352 VCC.n6260 0.00486429
R12916 VCC.n6354 VCC.n6353 0.00486429
R12917 VCC.n6375 VCC.n6242 0.00486429
R12918 VCC.n6465 VCC.n6197 0.00486429
R12919 VCC.n6475 VCC.n6466 0.00486429
R12920 VCC.n6474 VCC.n6467 0.00486429
R12921 VCC.n6502 VCC.n6182 0.00486429
R12922 VCC.n6580 VCC.n6579 0.00486429
R12923 VCC.n6598 VCC.n6130 0.00486429
R12924 VCC.n6600 VCC.n6599 0.00486429
R12925 VCC.n6607 VCC.n6125 0.00486429
R12926 VCC.n6895 VCC.n6894 0.00486429
R12927 VCC.n6909 VCC.n6817 0.00486429
R12928 VCC.n6911 VCC.n6910 0.00486429
R12929 VCC.n6932 VCC.n6799 0.00486429
R12930 VCC.n7021 VCC.n6753 0.00486429
R12931 VCC.n7031 VCC.n7022 0.00486429
R12932 VCC.n7030 VCC.n7023 0.00486429
R12933 VCC.n7058 VCC.n6738 0.00486429
R12934 VCC.n7143 VCC.n7142 0.00486429
R12935 VCC.n7150 VCC.n6692 0.00486429
R12936 VCC.n7154 VCC.n7153 0.00486429
R12937 VCC.n7170 VCC.n6672 0.00486429
R12938 VCC.n7445 VCC.n7444 0.00486429
R12939 VCC.n7459 VCC.n7367 0.00486429
R12940 VCC.n7461 VCC.n7460 0.00486429
R12941 VCC.n7482 VCC.n7349 0.00486429
R12942 VCC.n7572 VCC.n7304 0.00486429
R12943 VCC.n7582 VCC.n7573 0.00486429
R12944 VCC.n7581 VCC.n7574 0.00486429
R12945 VCC.n7609 VCC.n7289 0.00486429
R12946 VCC.n7687 VCC.n7686 0.00486429
R12947 VCC.n7705 VCC.n7237 0.00486429
R12948 VCC.n7707 VCC.n7706 0.00486429
R12949 VCC.n7714 VCC.n7232 0.00486429
R12950 VCC.n8002 VCC.n8001 0.00486429
R12951 VCC.n8016 VCC.n7924 0.00486429
R12952 VCC.n8018 VCC.n8017 0.00486429
R12953 VCC.n8039 VCC.n7906 0.00486429
R12954 VCC.n8128 VCC.n7860 0.00486429
R12955 VCC.n8138 VCC.n8129 0.00486429
R12956 VCC.n8137 VCC.n8130 0.00486429
R12957 VCC.n8165 VCC.n7845 0.00486429
R12958 VCC.n8250 VCC.n8249 0.00486429
R12959 VCC.n8257 VCC.n7799 0.00486429
R12960 VCC.n8261 VCC.n8260 0.00486429
R12961 VCC.n8277 VCC.n7779 0.00486429
R12962 VCC.n8492 VCC.n8411 0.00486429
R12963 VCC.n8502 VCC.n8493 0.00486429
R12964 VCC.n8501 VCC.n8494 0.00486429
R12965 VCC.n8529 VCC.n8396 0.00486429
R12966 VCC.n8607 VCC.n8606 0.00486429
R12967 VCC.n8625 VCC.n8344 0.00486429
R12968 VCC.n8627 VCC.n8626 0.00486429
R12969 VCC.n8634 VCC.n8339 0.00486429
R12970 VCC.n203 VCC.n202 0.00407143
R12971 VCC.n250 VCC.n168 0.00407143
R12972 VCC.n255 VCC.n251 0.00407143
R12973 VCC.n305 VCC.n134 0.00407143
R12974 VCC.n256 VCC.n166 0.00407143
R12975 VCC.n377 VCC.n96 0.00407143
R12976 VCC.n434 VCC.n76 0.00407143
R12977 VCC.n378 VCC.n375 0.00407143
R12978 VCC.n755 VCC.n754 0.00407143
R12979 VCC.n802 VCC.n720 0.00407143
R12980 VCC.n807 VCC.n803 0.00407143
R12981 VCC.n857 VCC.n686 0.00407143
R12982 VCC.n808 VCC.n718 0.00407143
R12983 VCC.n929 VCC.n648 0.00407143
R12984 VCC.n986 VCC.n628 0.00407143
R12985 VCC.n930 VCC.n927 0.00407143
R12986 VCC.n1486 VCC.n1205 0.00407143
R12987 VCC.n1544 VCC.n1185 0.00407143
R12988 VCC.n1487 VCC.n1484 0.00407143
R12989 VCC.n1313 VCC.n1312 0.00407143
R12990 VCC.n1360 VCC.n1278 0.00407143
R12991 VCC.n1365 VCC.n1361 0.00407143
R12992 VCC.n1415 VCC.n1244 0.00407143
R12993 VCC.n1366 VCC.n1276 0.00407143
R12994 VCC.n1864 VCC.n1863 0.00407143
R12995 VCC.n1911 VCC.n1829 0.00407143
R12996 VCC.n1916 VCC.n1912 0.00407143
R12997 VCC.n1966 VCC.n1795 0.00407143
R12998 VCC.n1917 VCC.n1827 0.00407143
R12999 VCC.n2038 VCC.n1757 0.00407143
R13000 VCC.n2095 VCC.n1737 0.00407143
R13001 VCC.n2039 VCC.n2036 0.00407143
R13002 VCC.n2595 VCC.n2314 0.00407143
R13003 VCC.n2653 VCC.n2294 0.00407143
R13004 VCC.n2596 VCC.n2593 0.00407143
R13005 VCC.n2422 VCC.n2421 0.00407143
R13006 VCC.n2469 VCC.n2387 0.00407143
R13007 VCC.n2474 VCC.n2470 0.00407143
R13008 VCC.n2524 VCC.n2353 0.00407143
R13009 VCC.n2475 VCC.n2385 0.00407143
R13010 VCC.n2973 VCC.n2972 0.00407143
R13011 VCC.n3020 VCC.n2938 0.00407143
R13012 VCC.n3025 VCC.n3021 0.00407143
R13013 VCC.n3075 VCC.n2904 0.00407143
R13014 VCC.n3026 VCC.n2936 0.00407143
R13015 VCC.n3147 VCC.n2866 0.00407143
R13016 VCC.n3204 VCC.n2846 0.00407143
R13017 VCC.n3148 VCC.n3145 0.00407143
R13018 VCC.n3704 VCC.n3423 0.00407143
R13019 VCC.n3762 VCC.n3403 0.00407143
R13020 VCC.n3705 VCC.n3702 0.00407143
R13021 VCC.n3531 VCC.n3530 0.00407143
R13022 VCC.n3578 VCC.n3496 0.00407143
R13023 VCC.n3583 VCC.n3579 0.00407143
R13024 VCC.n3633 VCC.n3462 0.00407143
R13025 VCC.n3584 VCC.n3494 0.00407143
R13026 VCC.n4082 VCC.n4081 0.00407143
R13027 VCC.n4129 VCC.n4047 0.00407143
R13028 VCC.n4134 VCC.n4130 0.00407143
R13029 VCC.n4184 VCC.n4013 0.00407143
R13030 VCC.n4135 VCC.n4045 0.00407143
R13031 VCC.n4256 VCC.n3975 0.00407143
R13032 VCC.n4313 VCC.n3955 0.00407143
R13033 VCC.n4257 VCC.n4254 0.00407143
R13034 VCC.n4813 VCC.n4532 0.00407143
R13035 VCC.n4871 VCC.n4512 0.00407143
R13036 VCC.n4814 VCC.n4811 0.00407143
R13037 VCC.n4640 VCC.n4639 0.00407143
R13038 VCC.n4687 VCC.n4605 0.00407143
R13039 VCC.n4692 VCC.n4688 0.00407143
R13040 VCC.n4742 VCC.n4571 0.00407143
R13041 VCC.n4693 VCC.n4603 0.00407143
R13042 VCC.n5191 VCC.n5190 0.00407143
R13043 VCC.n5238 VCC.n5156 0.00407143
R13044 VCC.n5243 VCC.n5239 0.00407143
R13045 VCC.n5293 VCC.n5122 0.00407143
R13046 VCC.n5244 VCC.n5154 0.00407143
R13047 VCC.n5365 VCC.n5084 0.00407143
R13048 VCC.n5422 VCC.n5064 0.00407143
R13049 VCC.n5366 VCC.n5363 0.00407143
R13050 VCC.n5921 VCC.n5640 0.00407143
R13051 VCC.n5979 VCC.n5620 0.00407143
R13052 VCC.n5922 VCC.n5919 0.00407143
R13053 VCC.n5748 VCC.n5747 0.00407143
R13054 VCC.n5795 VCC.n5713 0.00407143
R13055 VCC.n5800 VCC.n5796 0.00407143
R13056 VCC.n5850 VCC.n5679 0.00407143
R13057 VCC.n5801 VCC.n5711 0.00407143
R13058 VCC.n6298 VCC.n6297 0.00407143
R13059 VCC.n6345 VCC.n6263 0.00407143
R13060 VCC.n6350 VCC.n6346 0.00407143
R13061 VCC.n6400 VCC.n6229 0.00407143
R13062 VCC.n6351 VCC.n6261 0.00407143
R13063 VCC.n6472 VCC.n6191 0.00407143
R13064 VCC.n6529 VCC.n6171 0.00407143
R13065 VCC.n6473 VCC.n6470 0.00407143
R13066 VCC.n7028 VCC.n6747 0.00407143
R13067 VCC.n7086 VCC.n6727 0.00407143
R13068 VCC.n7029 VCC.n7026 0.00407143
R13069 VCC.n6855 VCC.n6854 0.00407143
R13070 VCC.n6902 VCC.n6820 0.00407143
R13071 VCC.n6907 VCC.n6903 0.00407143
R13072 VCC.n6957 VCC.n6786 0.00407143
R13073 VCC.n6908 VCC.n6818 0.00407143
R13074 VCC.n7405 VCC.n7404 0.00407143
R13075 VCC.n7452 VCC.n7370 0.00407143
R13076 VCC.n7457 VCC.n7453 0.00407143
R13077 VCC.n7507 VCC.n7336 0.00407143
R13078 VCC.n7458 VCC.n7368 0.00407143
R13079 VCC.n7579 VCC.n7298 0.00407143
R13080 VCC.n7636 VCC.n7278 0.00407143
R13081 VCC.n7580 VCC.n7577 0.00407143
R13082 VCC.n8135 VCC.n7854 0.00407143
R13083 VCC.n8193 VCC.n7834 0.00407143
R13084 VCC.n8136 VCC.n8133 0.00407143
R13085 VCC.n7962 VCC.n7961 0.00407143
R13086 VCC.n8009 VCC.n7927 0.00407143
R13087 VCC.n8014 VCC.n8010 0.00407143
R13088 VCC.n8064 VCC.n7893 0.00407143
R13089 VCC.n8015 VCC.n7925 0.00407143
R13090 VCC.n8499 VCC.n8405 0.00407143
R13091 VCC.n8556 VCC.n8385 0.00407143
R13092 VCC.n8500 VCC.n8497 0.00407143
R13093 VCC.n243 VCC.n165 0.00318571
R13094 VCC.n259 VCC.n147 0.00318571
R13095 VCC.n371 VCC.n370 0.00318571
R13096 VCC.n372 VCC.n87 0.00318571
R13097 VCC.n484 VCC.n35 0.00318571
R13098 VCC.n505 VCC.n30 0.00318571
R13099 VCC.n795 VCC.n717 0.00318571
R13100 VCC.n811 VCC.n699 0.00318571
R13101 VCC.n923 VCC.n922 0.00318571
R13102 VCC.n924 VCC.n639 0.00318571
R13103 VCC.n1036 VCC.n587 0.00318571
R13104 VCC.n1057 VCC.n582 0.00318571
R13105 VCC.n1353 VCC.n1275 0.00318571
R13106 VCC.n1369 VCC.n1257 0.00318571
R13107 VCC.n1480 VCC.n1479 0.00318571
R13108 VCC.n1481 VCC.n1196 0.00318571
R13109 VCC.n1601 VCC.n1150 0.00318571
R13110 VCC.n1611 VCC.n1130 0.00318571
R13111 VCC.n1904 VCC.n1826 0.00318571
R13112 VCC.n1920 VCC.n1808 0.00318571
R13113 VCC.n2032 VCC.n2031 0.00318571
R13114 VCC.n2033 VCC.n1748 0.00318571
R13115 VCC.n2145 VCC.n1696 0.00318571
R13116 VCC.n2166 VCC.n1691 0.00318571
R13117 VCC.n2462 VCC.n2384 0.00318571
R13118 VCC.n2478 VCC.n2366 0.00318571
R13119 VCC.n2589 VCC.n2588 0.00318571
R13120 VCC.n2590 VCC.n2305 0.00318571
R13121 VCC.n2710 VCC.n2259 0.00318571
R13122 VCC.n2720 VCC.n2239 0.00318571
R13123 VCC.n3013 VCC.n2935 0.00318571
R13124 VCC.n3029 VCC.n2917 0.00318571
R13125 VCC.n3141 VCC.n3140 0.00318571
R13126 VCC.n3142 VCC.n2857 0.00318571
R13127 VCC.n3254 VCC.n2805 0.00318571
R13128 VCC.n3275 VCC.n2800 0.00318571
R13129 VCC.n3571 VCC.n3493 0.00318571
R13130 VCC.n3587 VCC.n3475 0.00318571
R13131 VCC.n3698 VCC.n3697 0.00318571
R13132 VCC.n3699 VCC.n3414 0.00318571
R13133 VCC.n3819 VCC.n3368 0.00318571
R13134 VCC.n3829 VCC.n3348 0.00318571
R13135 VCC.n4122 VCC.n4044 0.00318571
R13136 VCC.n4138 VCC.n4026 0.00318571
R13137 VCC.n4250 VCC.n4249 0.00318571
R13138 VCC.n4251 VCC.n3966 0.00318571
R13139 VCC.n4363 VCC.n3914 0.00318571
R13140 VCC.n4384 VCC.n3909 0.00318571
R13141 VCC.n4680 VCC.n4602 0.00318571
R13142 VCC.n4696 VCC.n4584 0.00318571
R13143 VCC.n4807 VCC.n4806 0.00318571
R13144 VCC.n4808 VCC.n4523 0.00318571
R13145 VCC.n4928 VCC.n4477 0.00318571
R13146 VCC.n4938 VCC.n4457 0.00318571
R13147 VCC.n5231 VCC.n5153 0.00318571
R13148 VCC.n5247 VCC.n5135 0.00318571
R13149 VCC.n5359 VCC.n5358 0.00318571
R13150 VCC.n5360 VCC.n5075 0.00318571
R13151 VCC.n5472 VCC.n5023 0.00318571
R13152 VCC.n5493 VCC.n5018 0.00318571
R13153 VCC.n5788 VCC.n5710 0.00318571
R13154 VCC.n5804 VCC.n5692 0.00318571
R13155 VCC.n5915 VCC.n5914 0.00318571
R13156 VCC.n5916 VCC.n5631 0.00318571
R13157 VCC.n6036 VCC.n5585 0.00318571
R13158 VCC.n6046 VCC.n5565 0.00318571
R13159 VCC.n6338 VCC.n6260 0.00318571
R13160 VCC.n6354 VCC.n6242 0.00318571
R13161 VCC.n6466 VCC.n6465 0.00318571
R13162 VCC.n6467 VCC.n6182 0.00318571
R13163 VCC.n6579 VCC.n6130 0.00318571
R13164 VCC.n6600 VCC.n6125 0.00318571
R13165 VCC.n6895 VCC.n6817 0.00318571
R13166 VCC.n6911 VCC.n6799 0.00318571
R13167 VCC.n7022 VCC.n7021 0.00318571
R13168 VCC.n7023 VCC.n6738 0.00318571
R13169 VCC.n7143 VCC.n6692 0.00318571
R13170 VCC.n7153 VCC.n6672 0.00318571
R13171 VCC.n7445 VCC.n7367 0.00318571
R13172 VCC.n7461 VCC.n7349 0.00318571
R13173 VCC.n7573 VCC.n7572 0.00318571
R13174 VCC.n7574 VCC.n7289 0.00318571
R13175 VCC.n7686 VCC.n7237 0.00318571
R13176 VCC.n7707 VCC.n7232 0.00318571
R13177 VCC.n8002 VCC.n7924 0.00318571
R13178 VCC.n8018 VCC.n7906 0.00318571
R13179 VCC.n8129 VCC.n8128 0.00318571
R13180 VCC.n8130 VCC.n7845 0.00318571
R13181 VCC.n8250 VCC.n7799 0.00318571
R13182 VCC.n8260 VCC.n7779 0.00318571
R13183 VCC.n8493 VCC.n8492 0.00318571
R13184 VCC.n8494 VCC.n8396 0.00318571
R13185 VCC.n8606 VCC.n8344 0.00318571
R13186 VCC.n8627 VCC.n8339 0.00318571
R13187 VCC.n220 VCC.n185 0.00317857
R13188 VCC.n262 VCC.n157 0.00317857
R13189 VCC.n305 VCC.n304 0.00317857
R13190 VCC.n310 VCC.n129 0.00317857
R13191 VCC.n216 VCC.n190 0.00317857
R13192 VCC.n219 VCC.n186 0.00317857
R13193 VCC.n261 VCC.n163 0.00317857
R13194 VCC.n306 VCC.n133 0.00317857
R13195 VCC.n309 VCC.n130 0.00317857
R13196 VCC.n332 VCC.n125 0.00317857
R13197 VCC.n343 VCC.n116 0.00317857
R13198 VCC.n343 VCC.n342 0.00317857
R13199 VCC.n105 VCC.n98 0.00317857
R13200 VCC.n383 VCC.n99 0.00317857
R13201 VCC.n389 VCC.n388 0.00317857
R13202 VCC.n440 VCC.n73 0.00317857
R13203 VCC.n440 VCC.n439 0.00317857
R13204 VCC.n445 VCC.n68 0.00317857
R13205 VCC.n319 VCC.n318 0.00317857
R13206 VCC.n344 VCC.n115 0.00317857
R13207 VCC.n382 VCC.n381 0.00317857
R13208 VCC.n441 VCC.n72 0.00317857
R13209 VCC.n444 VCC.n69 0.00317857
R13210 VCC.n458 VCC.n457 0.00317857
R13211 VCC.n463 VCC.n59 0.00317857
R13212 VCC.n508 VCC.n32 0.00317857
R13213 VCC.n517 VCC.n516 0.00317857
R13214 VCC.n534 VCC.n533 0.00317857
R13215 VCC.n12 VCC.n11 0.00317857
R13216 VCC.n12 VCC.n2 0.00317857
R13217 VCC.n459 VCC.n64 0.00317857
R13218 VCC.n465 VCC.n464 0.00317857
R13219 VCC.n507 VCC.n33 0.00317857
R13220 VCC.n535 VCC.n15 0.00317857
R13221 VCC.n539 VCC.n538 0.00317857
R13222 VCC.n772 VCC.n737 0.00317857
R13223 VCC.n814 VCC.n709 0.00317857
R13224 VCC.n857 VCC.n856 0.00317857
R13225 VCC.n862 VCC.n681 0.00317857
R13226 VCC.n768 VCC.n742 0.00317857
R13227 VCC.n771 VCC.n738 0.00317857
R13228 VCC.n813 VCC.n715 0.00317857
R13229 VCC.n858 VCC.n685 0.00317857
R13230 VCC.n861 VCC.n682 0.00317857
R13231 VCC.n884 VCC.n677 0.00317857
R13232 VCC.n895 VCC.n668 0.00317857
R13233 VCC.n895 VCC.n894 0.00317857
R13234 VCC.n657 VCC.n650 0.00317857
R13235 VCC.n935 VCC.n651 0.00317857
R13236 VCC.n941 VCC.n940 0.00317857
R13237 VCC.n992 VCC.n625 0.00317857
R13238 VCC.n992 VCC.n991 0.00317857
R13239 VCC.n997 VCC.n620 0.00317857
R13240 VCC.n871 VCC.n870 0.00317857
R13241 VCC.n896 VCC.n667 0.00317857
R13242 VCC.n934 VCC.n933 0.00317857
R13243 VCC.n993 VCC.n624 0.00317857
R13244 VCC.n996 VCC.n621 0.00317857
R13245 VCC.n1010 VCC.n1009 0.00317857
R13246 VCC.n1015 VCC.n611 0.00317857
R13247 VCC.n1060 VCC.n584 0.00317857
R13248 VCC.n1069 VCC.n1068 0.00317857
R13249 VCC.n1086 VCC.n1085 0.00317857
R13250 VCC.n1092 VCC.n1091 0.00317857
R13251 VCC.n1092 VCC.n556 0.00317857
R13252 VCC.n1011 VCC.n616 0.00317857
R13253 VCC.n1017 VCC.n1016 0.00317857
R13254 VCC.n1059 VCC.n585 0.00317857
R13255 VCC.n1087 VCC.n567 0.00317857
R13256 VCC.n1093 VCC.n1090 0.00317857
R13257 VCC.n1569 VCC.n1568 0.00317857
R13258 VCC.n1575 VCC.n1169 0.00317857
R13259 VCC.n1614 VCC.n1148 0.00317857
R13260 VCC.n1139 VCC.n1128 0.00317857
R13261 VCC.n1633 VCC.n1118 0.00317857
R13262 VCC.n1640 VCC.n1639 0.00317857
R13263 VCC.n1639 VCC.n1110 0.00317857
R13264 VCC.n1570 VCC.n1173 0.00317857
R13265 VCC.n1574 VCC.n1573 0.00317857
R13266 VCC.n1613 VCC.n1149 0.00317857
R13267 VCC.n1634 VCC.n1120 0.00317857
R13268 VCC.n1638 VCC.n1637 0.00317857
R13269 VCC.n1441 VCC.n1234 0.00317857
R13270 VCC.n1452 VCC.n1225 0.00317857
R13271 VCC.n1452 VCC.n1451 0.00317857
R13272 VCC.n1214 VCC.n1207 0.00317857
R13273 VCC.n1492 VCC.n1208 0.00317857
R13274 VCC.n1498 VCC.n1497 0.00317857
R13275 VCC.n1550 VCC.n1182 0.00317857
R13276 VCC.n1550 VCC.n1549 0.00317857
R13277 VCC.n1555 VCC.n1177 0.00317857
R13278 VCC.n1440 VCC.n1428 0.00317857
R13279 VCC.n1453 VCC.n1224 0.00317857
R13280 VCC.n1491 VCC.n1490 0.00317857
R13281 VCC.n1551 VCC.n1181 0.00317857
R13282 VCC.n1554 VCC.n1178 0.00317857
R13283 VCC.n1330 VCC.n1295 0.00317857
R13284 VCC.n1372 VCC.n1267 0.00317857
R13285 VCC.n1415 VCC.n1414 0.00317857
R13286 VCC.n1420 VCC.n1239 0.00317857
R13287 VCC.n1326 VCC.n1300 0.00317857
R13288 VCC.n1329 VCC.n1296 0.00317857
R13289 VCC.n1371 VCC.n1273 0.00317857
R13290 VCC.n1416 VCC.n1243 0.00317857
R13291 VCC.n1419 VCC.n1240 0.00317857
R13292 VCC.n1881 VCC.n1846 0.00317857
R13293 VCC.n1923 VCC.n1818 0.00317857
R13294 VCC.n1966 VCC.n1965 0.00317857
R13295 VCC.n1971 VCC.n1790 0.00317857
R13296 VCC.n1877 VCC.n1851 0.00317857
R13297 VCC.n1880 VCC.n1847 0.00317857
R13298 VCC.n1922 VCC.n1824 0.00317857
R13299 VCC.n1967 VCC.n1794 0.00317857
R13300 VCC.n1970 VCC.n1791 0.00317857
R13301 VCC.n1993 VCC.n1786 0.00317857
R13302 VCC.n2004 VCC.n1777 0.00317857
R13303 VCC.n2004 VCC.n2003 0.00317857
R13304 VCC.n1766 VCC.n1759 0.00317857
R13305 VCC.n2044 VCC.n1760 0.00317857
R13306 VCC.n2050 VCC.n2049 0.00317857
R13307 VCC.n2101 VCC.n1734 0.00317857
R13308 VCC.n2101 VCC.n2100 0.00317857
R13309 VCC.n2106 VCC.n1729 0.00317857
R13310 VCC.n1980 VCC.n1979 0.00317857
R13311 VCC.n2005 VCC.n1776 0.00317857
R13312 VCC.n2043 VCC.n2042 0.00317857
R13313 VCC.n2102 VCC.n1733 0.00317857
R13314 VCC.n2105 VCC.n1730 0.00317857
R13315 VCC.n2119 VCC.n2118 0.00317857
R13316 VCC.n2124 VCC.n1720 0.00317857
R13317 VCC.n2169 VCC.n1693 0.00317857
R13318 VCC.n2178 VCC.n2177 0.00317857
R13319 VCC.n2195 VCC.n2194 0.00317857
R13320 VCC.n2201 VCC.n2200 0.00317857
R13321 VCC.n2201 VCC.n1665 0.00317857
R13322 VCC.n2120 VCC.n1725 0.00317857
R13323 VCC.n2126 VCC.n2125 0.00317857
R13324 VCC.n2168 VCC.n1694 0.00317857
R13325 VCC.n2196 VCC.n1676 0.00317857
R13326 VCC.n2202 VCC.n2199 0.00317857
R13327 VCC.n2678 VCC.n2677 0.00317857
R13328 VCC.n2684 VCC.n2278 0.00317857
R13329 VCC.n2723 VCC.n2257 0.00317857
R13330 VCC.n2248 VCC.n2237 0.00317857
R13331 VCC.n2742 VCC.n2227 0.00317857
R13332 VCC.n2749 VCC.n2748 0.00317857
R13333 VCC.n2748 VCC.n2219 0.00317857
R13334 VCC.n2679 VCC.n2282 0.00317857
R13335 VCC.n2683 VCC.n2682 0.00317857
R13336 VCC.n2722 VCC.n2258 0.00317857
R13337 VCC.n2743 VCC.n2229 0.00317857
R13338 VCC.n2747 VCC.n2746 0.00317857
R13339 VCC.n2550 VCC.n2343 0.00317857
R13340 VCC.n2561 VCC.n2334 0.00317857
R13341 VCC.n2561 VCC.n2560 0.00317857
R13342 VCC.n2323 VCC.n2316 0.00317857
R13343 VCC.n2601 VCC.n2317 0.00317857
R13344 VCC.n2607 VCC.n2606 0.00317857
R13345 VCC.n2659 VCC.n2291 0.00317857
R13346 VCC.n2659 VCC.n2658 0.00317857
R13347 VCC.n2664 VCC.n2286 0.00317857
R13348 VCC.n2549 VCC.n2537 0.00317857
R13349 VCC.n2562 VCC.n2333 0.00317857
R13350 VCC.n2600 VCC.n2599 0.00317857
R13351 VCC.n2660 VCC.n2290 0.00317857
R13352 VCC.n2663 VCC.n2287 0.00317857
R13353 VCC.n2439 VCC.n2404 0.00317857
R13354 VCC.n2481 VCC.n2376 0.00317857
R13355 VCC.n2524 VCC.n2523 0.00317857
R13356 VCC.n2529 VCC.n2348 0.00317857
R13357 VCC.n2435 VCC.n2409 0.00317857
R13358 VCC.n2438 VCC.n2405 0.00317857
R13359 VCC.n2480 VCC.n2382 0.00317857
R13360 VCC.n2525 VCC.n2352 0.00317857
R13361 VCC.n2528 VCC.n2349 0.00317857
R13362 VCC.n2990 VCC.n2955 0.00317857
R13363 VCC.n3032 VCC.n2927 0.00317857
R13364 VCC.n3075 VCC.n3074 0.00317857
R13365 VCC.n3080 VCC.n2899 0.00317857
R13366 VCC.n2986 VCC.n2960 0.00317857
R13367 VCC.n2989 VCC.n2956 0.00317857
R13368 VCC.n3031 VCC.n2933 0.00317857
R13369 VCC.n3076 VCC.n2903 0.00317857
R13370 VCC.n3079 VCC.n2900 0.00317857
R13371 VCC.n3102 VCC.n2895 0.00317857
R13372 VCC.n3113 VCC.n2886 0.00317857
R13373 VCC.n3113 VCC.n3112 0.00317857
R13374 VCC.n2875 VCC.n2868 0.00317857
R13375 VCC.n3153 VCC.n2869 0.00317857
R13376 VCC.n3159 VCC.n3158 0.00317857
R13377 VCC.n3210 VCC.n2843 0.00317857
R13378 VCC.n3210 VCC.n3209 0.00317857
R13379 VCC.n3215 VCC.n2838 0.00317857
R13380 VCC.n3089 VCC.n3088 0.00317857
R13381 VCC.n3114 VCC.n2885 0.00317857
R13382 VCC.n3152 VCC.n3151 0.00317857
R13383 VCC.n3211 VCC.n2842 0.00317857
R13384 VCC.n3214 VCC.n2839 0.00317857
R13385 VCC.n3228 VCC.n3227 0.00317857
R13386 VCC.n3233 VCC.n2829 0.00317857
R13387 VCC.n3278 VCC.n2802 0.00317857
R13388 VCC.n3287 VCC.n3286 0.00317857
R13389 VCC.n3304 VCC.n3303 0.00317857
R13390 VCC.n3310 VCC.n3309 0.00317857
R13391 VCC.n3310 VCC.n2774 0.00317857
R13392 VCC.n3229 VCC.n2834 0.00317857
R13393 VCC.n3235 VCC.n3234 0.00317857
R13394 VCC.n3277 VCC.n2803 0.00317857
R13395 VCC.n3305 VCC.n2785 0.00317857
R13396 VCC.n3311 VCC.n3308 0.00317857
R13397 VCC.n3787 VCC.n3786 0.00317857
R13398 VCC.n3793 VCC.n3387 0.00317857
R13399 VCC.n3832 VCC.n3366 0.00317857
R13400 VCC.n3357 VCC.n3346 0.00317857
R13401 VCC.n3851 VCC.n3336 0.00317857
R13402 VCC.n3858 VCC.n3857 0.00317857
R13403 VCC.n3857 VCC.n3328 0.00317857
R13404 VCC.n3788 VCC.n3391 0.00317857
R13405 VCC.n3792 VCC.n3791 0.00317857
R13406 VCC.n3831 VCC.n3367 0.00317857
R13407 VCC.n3852 VCC.n3338 0.00317857
R13408 VCC.n3856 VCC.n3855 0.00317857
R13409 VCC.n3659 VCC.n3452 0.00317857
R13410 VCC.n3670 VCC.n3443 0.00317857
R13411 VCC.n3670 VCC.n3669 0.00317857
R13412 VCC.n3432 VCC.n3425 0.00317857
R13413 VCC.n3710 VCC.n3426 0.00317857
R13414 VCC.n3716 VCC.n3715 0.00317857
R13415 VCC.n3768 VCC.n3400 0.00317857
R13416 VCC.n3768 VCC.n3767 0.00317857
R13417 VCC.n3773 VCC.n3395 0.00317857
R13418 VCC.n3658 VCC.n3646 0.00317857
R13419 VCC.n3671 VCC.n3442 0.00317857
R13420 VCC.n3709 VCC.n3708 0.00317857
R13421 VCC.n3769 VCC.n3399 0.00317857
R13422 VCC.n3772 VCC.n3396 0.00317857
R13423 VCC.n3548 VCC.n3513 0.00317857
R13424 VCC.n3590 VCC.n3485 0.00317857
R13425 VCC.n3633 VCC.n3632 0.00317857
R13426 VCC.n3638 VCC.n3457 0.00317857
R13427 VCC.n3544 VCC.n3518 0.00317857
R13428 VCC.n3547 VCC.n3514 0.00317857
R13429 VCC.n3589 VCC.n3491 0.00317857
R13430 VCC.n3634 VCC.n3461 0.00317857
R13431 VCC.n3637 VCC.n3458 0.00317857
R13432 VCC.n4099 VCC.n4064 0.00317857
R13433 VCC.n4141 VCC.n4036 0.00317857
R13434 VCC.n4184 VCC.n4183 0.00317857
R13435 VCC.n4189 VCC.n4008 0.00317857
R13436 VCC.n4095 VCC.n4069 0.00317857
R13437 VCC.n4098 VCC.n4065 0.00317857
R13438 VCC.n4140 VCC.n4042 0.00317857
R13439 VCC.n4185 VCC.n4012 0.00317857
R13440 VCC.n4188 VCC.n4009 0.00317857
R13441 VCC.n4211 VCC.n4004 0.00317857
R13442 VCC.n4222 VCC.n3995 0.00317857
R13443 VCC.n4222 VCC.n4221 0.00317857
R13444 VCC.n3984 VCC.n3977 0.00317857
R13445 VCC.n4262 VCC.n3978 0.00317857
R13446 VCC.n4268 VCC.n4267 0.00317857
R13447 VCC.n4319 VCC.n3952 0.00317857
R13448 VCC.n4319 VCC.n4318 0.00317857
R13449 VCC.n4324 VCC.n3947 0.00317857
R13450 VCC.n4198 VCC.n4197 0.00317857
R13451 VCC.n4223 VCC.n3994 0.00317857
R13452 VCC.n4261 VCC.n4260 0.00317857
R13453 VCC.n4320 VCC.n3951 0.00317857
R13454 VCC.n4323 VCC.n3948 0.00317857
R13455 VCC.n4337 VCC.n4336 0.00317857
R13456 VCC.n4342 VCC.n3938 0.00317857
R13457 VCC.n4387 VCC.n3911 0.00317857
R13458 VCC.n4396 VCC.n4395 0.00317857
R13459 VCC.n4413 VCC.n4412 0.00317857
R13460 VCC.n4419 VCC.n4418 0.00317857
R13461 VCC.n4419 VCC.n3883 0.00317857
R13462 VCC.n4338 VCC.n3943 0.00317857
R13463 VCC.n4344 VCC.n4343 0.00317857
R13464 VCC.n4386 VCC.n3912 0.00317857
R13465 VCC.n4414 VCC.n3894 0.00317857
R13466 VCC.n4420 VCC.n4417 0.00317857
R13467 VCC.n4896 VCC.n4895 0.00317857
R13468 VCC.n4902 VCC.n4496 0.00317857
R13469 VCC.n4941 VCC.n4475 0.00317857
R13470 VCC.n4466 VCC.n4455 0.00317857
R13471 VCC.n4960 VCC.n4445 0.00317857
R13472 VCC.n4967 VCC.n4966 0.00317857
R13473 VCC.n4966 VCC.n4437 0.00317857
R13474 VCC.n4897 VCC.n4500 0.00317857
R13475 VCC.n4901 VCC.n4900 0.00317857
R13476 VCC.n4940 VCC.n4476 0.00317857
R13477 VCC.n4961 VCC.n4447 0.00317857
R13478 VCC.n4965 VCC.n4964 0.00317857
R13479 VCC.n4768 VCC.n4561 0.00317857
R13480 VCC.n4779 VCC.n4552 0.00317857
R13481 VCC.n4779 VCC.n4778 0.00317857
R13482 VCC.n4541 VCC.n4534 0.00317857
R13483 VCC.n4819 VCC.n4535 0.00317857
R13484 VCC.n4825 VCC.n4824 0.00317857
R13485 VCC.n4877 VCC.n4509 0.00317857
R13486 VCC.n4877 VCC.n4876 0.00317857
R13487 VCC.n4882 VCC.n4504 0.00317857
R13488 VCC.n4767 VCC.n4755 0.00317857
R13489 VCC.n4780 VCC.n4551 0.00317857
R13490 VCC.n4818 VCC.n4817 0.00317857
R13491 VCC.n4878 VCC.n4508 0.00317857
R13492 VCC.n4881 VCC.n4505 0.00317857
R13493 VCC.n4657 VCC.n4622 0.00317857
R13494 VCC.n4699 VCC.n4594 0.00317857
R13495 VCC.n4742 VCC.n4741 0.00317857
R13496 VCC.n4747 VCC.n4566 0.00317857
R13497 VCC.n4653 VCC.n4627 0.00317857
R13498 VCC.n4656 VCC.n4623 0.00317857
R13499 VCC.n4698 VCC.n4600 0.00317857
R13500 VCC.n4743 VCC.n4570 0.00317857
R13501 VCC.n4746 VCC.n4567 0.00317857
R13502 VCC.n5208 VCC.n5173 0.00317857
R13503 VCC.n5250 VCC.n5145 0.00317857
R13504 VCC.n5293 VCC.n5292 0.00317857
R13505 VCC.n5298 VCC.n5117 0.00317857
R13506 VCC.n5204 VCC.n5178 0.00317857
R13507 VCC.n5207 VCC.n5174 0.00317857
R13508 VCC.n5249 VCC.n5151 0.00317857
R13509 VCC.n5294 VCC.n5121 0.00317857
R13510 VCC.n5297 VCC.n5118 0.00317857
R13511 VCC.n5320 VCC.n5113 0.00317857
R13512 VCC.n5331 VCC.n5104 0.00317857
R13513 VCC.n5331 VCC.n5330 0.00317857
R13514 VCC.n5093 VCC.n5086 0.00317857
R13515 VCC.n5371 VCC.n5087 0.00317857
R13516 VCC.n5377 VCC.n5376 0.00317857
R13517 VCC.n5428 VCC.n5061 0.00317857
R13518 VCC.n5428 VCC.n5427 0.00317857
R13519 VCC.n5433 VCC.n5056 0.00317857
R13520 VCC.n5307 VCC.n5306 0.00317857
R13521 VCC.n5332 VCC.n5103 0.00317857
R13522 VCC.n5370 VCC.n5369 0.00317857
R13523 VCC.n5429 VCC.n5060 0.00317857
R13524 VCC.n5432 VCC.n5057 0.00317857
R13525 VCC.n5446 VCC.n5445 0.00317857
R13526 VCC.n5451 VCC.n5047 0.00317857
R13527 VCC.n5496 VCC.n5020 0.00317857
R13528 VCC.n5505 VCC.n5504 0.00317857
R13529 VCC.n5522 VCC.n5521 0.00317857
R13530 VCC.n5528 VCC.n5527 0.00317857
R13531 VCC.n5528 VCC.n4992 0.00317857
R13532 VCC.n5447 VCC.n5052 0.00317857
R13533 VCC.n5453 VCC.n5452 0.00317857
R13534 VCC.n5495 VCC.n5021 0.00317857
R13535 VCC.n5523 VCC.n5003 0.00317857
R13536 VCC.n5529 VCC.n5526 0.00317857
R13537 VCC.n6004 VCC.n6003 0.00317857
R13538 VCC.n6010 VCC.n5604 0.00317857
R13539 VCC.n6049 VCC.n5583 0.00317857
R13540 VCC.n5574 VCC.n5563 0.00317857
R13541 VCC.n6068 VCC.n5553 0.00317857
R13542 VCC.n6075 VCC.n6074 0.00317857
R13543 VCC.n6074 VCC.n5545 0.00317857
R13544 VCC.n6005 VCC.n5608 0.00317857
R13545 VCC.n6009 VCC.n6008 0.00317857
R13546 VCC.n6048 VCC.n5584 0.00317857
R13547 VCC.n6069 VCC.n5555 0.00317857
R13548 VCC.n6073 VCC.n6072 0.00317857
R13549 VCC.n5876 VCC.n5669 0.00317857
R13550 VCC.n5887 VCC.n5660 0.00317857
R13551 VCC.n5887 VCC.n5886 0.00317857
R13552 VCC.n5649 VCC.n5642 0.00317857
R13553 VCC.n5927 VCC.n5643 0.00317857
R13554 VCC.n5933 VCC.n5932 0.00317857
R13555 VCC.n5985 VCC.n5617 0.00317857
R13556 VCC.n5985 VCC.n5984 0.00317857
R13557 VCC.n5990 VCC.n5612 0.00317857
R13558 VCC.n5875 VCC.n5863 0.00317857
R13559 VCC.n5888 VCC.n5659 0.00317857
R13560 VCC.n5926 VCC.n5925 0.00317857
R13561 VCC.n5986 VCC.n5616 0.00317857
R13562 VCC.n5989 VCC.n5613 0.00317857
R13563 VCC.n5765 VCC.n5730 0.00317857
R13564 VCC.n5807 VCC.n5702 0.00317857
R13565 VCC.n5850 VCC.n5849 0.00317857
R13566 VCC.n5855 VCC.n5674 0.00317857
R13567 VCC.n5761 VCC.n5735 0.00317857
R13568 VCC.n5764 VCC.n5731 0.00317857
R13569 VCC.n5806 VCC.n5708 0.00317857
R13570 VCC.n5851 VCC.n5678 0.00317857
R13571 VCC.n5854 VCC.n5675 0.00317857
R13572 VCC.n6315 VCC.n6280 0.00317857
R13573 VCC.n6357 VCC.n6252 0.00317857
R13574 VCC.n6400 VCC.n6399 0.00317857
R13575 VCC.n6405 VCC.n6224 0.00317857
R13576 VCC.n6311 VCC.n6285 0.00317857
R13577 VCC.n6314 VCC.n6281 0.00317857
R13578 VCC.n6356 VCC.n6258 0.00317857
R13579 VCC.n6401 VCC.n6228 0.00317857
R13580 VCC.n6404 VCC.n6225 0.00317857
R13581 VCC.n6427 VCC.n6220 0.00317857
R13582 VCC.n6438 VCC.n6211 0.00317857
R13583 VCC.n6438 VCC.n6437 0.00317857
R13584 VCC.n6200 VCC.n6193 0.00317857
R13585 VCC.n6478 VCC.n6194 0.00317857
R13586 VCC.n6484 VCC.n6483 0.00317857
R13587 VCC.n6535 VCC.n6168 0.00317857
R13588 VCC.n6535 VCC.n6534 0.00317857
R13589 VCC.n6540 VCC.n6163 0.00317857
R13590 VCC.n6414 VCC.n6413 0.00317857
R13591 VCC.n6439 VCC.n6210 0.00317857
R13592 VCC.n6477 VCC.n6476 0.00317857
R13593 VCC.n6536 VCC.n6167 0.00317857
R13594 VCC.n6539 VCC.n6164 0.00317857
R13595 VCC.n6553 VCC.n6552 0.00317857
R13596 VCC.n6558 VCC.n6154 0.00317857
R13597 VCC.n6603 VCC.n6127 0.00317857
R13598 VCC.n6612 VCC.n6611 0.00317857
R13599 VCC.n6629 VCC.n6628 0.00317857
R13600 VCC.n6635 VCC.n6634 0.00317857
R13601 VCC.n6635 VCC.n6099 0.00317857
R13602 VCC.n6554 VCC.n6159 0.00317857
R13603 VCC.n6560 VCC.n6559 0.00317857
R13604 VCC.n6602 VCC.n6128 0.00317857
R13605 VCC.n6630 VCC.n6110 0.00317857
R13606 VCC.n6636 VCC.n6633 0.00317857
R13607 VCC.n7111 VCC.n7110 0.00317857
R13608 VCC.n7117 VCC.n6711 0.00317857
R13609 VCC.n7156 VCC.n6690 0.00317857
R13610 VCC.n6681 VCC.n6670 0.00317857
R13611 VCC.n7175 VCC.n6660 0.00317857
R13612 VCC.n7182 VCC.n7181 0.00317857
R13613 VCC.n7181 VCC.n6652 0.00317857
R13614 VCC.n7112 VCC.n6715 0.00317857
R13615 VCC.n7116 VCC.n7115 0.00317857
R13616 VCC.n7155 VCC.n6691 0.00317857
R13617 VCC.n7176 VCC.n6662 0.00317857
R13618 VCC.n7180 VCC.n7179 0.00317857
R13619 VCC.n6983 VCC.n6776 0.00317857
R13620 VCC.n6994 VCC.n6767 0.00317857
R13621 VCC.n6994 VCC.n6993 0.00317857
R13622 VCC.n6756 VCC.n6749 0.00317857
R13623 VCC.n7034 VCC.n6750 0.00317857
R13624 VCC.n7040 VCC.n7039 0.00317857
R13625 VCC.n7092 VCC.n6724 0.00317857
R13626 VCC.n7092 VCC.n7091 0.00317857
R13627 VCC.n7097 VCC.n6719 0.00317857
R13628 VCC.n6982 VCC.n6970 0.00317857
R13629 VCC.n6995 VCC.n6766 0.00317857
R13630 VCC.n7033 VCC.n7032 0.00317857
R13631 VCC.n7093 VCC.n6723 0.00317857
R13632 VCC.n7096 VCC.n6720 0.00317857
R13633 VCC.n6872 VCC.n6837 0.00317857
R13634 VCC.n6914 VCC.n6809 0.00317857
R13635 VCC.n6957 VCC.n6956 0.00317857
R13636 VCC.n6962 VCC.n6781 0.00317857
R13637 VCC.n6868 VCC.n6842 0.00317857
R13638 VCC.n6871 VCC.n6838 0.00317857
R13639 VCC.n6913 VCC.n6815 0.00317857
R13640 VCC.n6958 VCC.n6785 0.00317857
R13641 VCC.n6961 VCC.n6782 0.00317857
R13642 VCC.n7422 VCC.n7387 0.00317857
R13643 VCC.n7464 VCC.n7359 0.00317857
R13644 VCC.n7507 VCC.n7506 0.00317857
R13645 VCC.n7512 VCC.n7331 0.00317857
R13646 VCC.n7418 VCC.n7392 0.00317857
R13647 VCC.n7421 VCC.n7388 0.00317857
R13648 VCC.n7463 VCC.n7365 0.00317857
R13649 VCC.n7508 VCC.n7335 0.00317857
R13650 VCC.n7511 VCC.n7332 0.00317857
R13651 VCC.n7534 VCC.n7327 0.00317857
R13652 VCC.n7545 VCC.n7318 0.00317857
R13653 VCC.n7545 VCC.n7544 0.00317857
R13654 VCC.n7307 VCC.n7300 0.00317857
R13655 VCC.n7585 VCC.n7301 0.00317857
R13656 VCC.n7591 VCC.n7590 0.00317857
R13657 VCC.n7642 VCC.n7275 0.00317857
R13658 VCC.n7642 VCC.n7641 0.00317857
R13659 VCC.n7647 VCC.n7270 0.00317857
R13660 VCC.n7521 VCC.n7520 0.00317857
R13661 VCC.n7546 VCC.n7317 0.00317857
R13662 VCC.n7584 VCC.n7583 0.00317857
R13663 VCC.n7643 VCC.n7274 0.00317857
R13664 VCC.n7646 VCC.n7271 0.00317857
R13665 VCC.n7660 VCC.n7659 0.00317857
R13666 VCC.n7665 VCC.n7261 0.00317857
R13667 VCC.n7710 VCC.n7234 0.00317857
R13668 VCC.n7719 VCC.n7718 0.00317857
R13669 VCC.n7736 VCC.n7735 0.00317857
R13670 VCC.n7742 VCC.n7741 0.00317857
R13671 VCC.n7742 VCC.n7206 0.00317857
R13672 VCC.n7661 VCC.n7266 0.00317857
R13673 VCC.n7667 VCC.n7666 0.00317857
R13674 VCC.n7709 VCC.n7235 0.00317857
R13675 VCC.n7737 VCC.n7217 0.00317857
R13676 VCC.n7743 VCC.n7740 0.00317857
R13677 VCC.n8218 VCC.n8217 0.00317857
R13678 VCC.n8224 VCC.n7818 0.00317857
R13679 VCC.n8263 VCC.n7797 0.00317857
R13680 VCC.n7788 VCC.n7777 0.00317857
R13681 VCC.n8282 VCC.n7767 0.00317857
R13682 VCC.n8289 VCC.n8288 0.00317857
R13683 VCC.n8288 VCC.n7759 0.00317857
R13684 VCC.n8219 VCC.n7822 0.00317857
R13685 VCC.n8223 VCC.n8222 0.00317857
R13686 VCC.n8262 VCC.n7798 0.00317857
R13687 VCC.n8283 VCC.n7769 0.00317857
R13688 VCC.n8287 VCC.n8286 0.00317857
R13689 VCC.n8090 VCC.n7883 0.00317857
R13690 VCC.n8101 VCC.n7874 0.00317857
R13691 VCC.n8101 VCC.n8100 0.00317857
R13692 VCC.n7863 VCC.n7856 0.00317857
R13693 VCC.n8141 VCC.n7857 0.00317857
R13694 VCC.n8147 VCC.n8146 0.00317857
R13695 VCC.n8199 VCC.n7831 0.00317857
R13696 VCC.n8199 VCC.n8198 0.00317857
R13697 VCC.n8204 VCC.n7826 0.00317857
R13698 VCC.n8089 VCC.n8077 0.00317857
R13699 VCC.n8102 VCC.n7873 0.00317857
R13700 VCC.n8140 VCC.n8139 0.00317857
R13701 VCC.n8200 VCC.n7830 0.00317857
R13702 VCC.n8203 VCC.n7827 0.00317857
R13703 VCC.n7979 VCC.n7944 0.00317857
R13704 VCC.n8021 VCC.n7916 0.00317857
R13705 VCC.n8064 VCC.n8063 0.00317857
R13706 VCC.n8069 VCC.n7888 0.00317857
R13707 VCC.n7975 VCC.n7949 0.00317857
R13708 VCC.n7978 VCC.n7945 0.00317857
R13709 VCC.n8020 VCC.n7922 0.00317857
R13710 VCC.n8065 VCC.n7892 0.00317857
R13711 VCC.n8068 VCC.n7889 0.00317857
R13712 VCC.n8454 VCC.n8434 0.00317857
R13713 VCC.n8465 VCC.n8425 0.00317857
R13714 VCC.n8465 VCC.n8464 0.00317857
R13715 VCC.n8414 VCC.n8407 0.00317857
R13716 VCC.n8505 VCC.n8408 0.00317857
R13717 VCC.n8511 VCC.n8510 0.00317857
R13718 VCC.n8562 VCC.n8382 0.00317857
R13719 VCC.n8562 VCC.n8561 0.00317857
R13720 VCC.n8567 VCC.n8377 0.00317857
R13721 VCC.n8441 VCC.n8440 0.00317857
R13722 VCC.n8466 VCC.n8424 0.00317857
R13723 VCC.n8504 VCC.n8503 0.00317857
R13724 VCC.n8563 VCC.n8381 0.00317857
R13725 VCC.n8566 VCC.n8378 0.00317857
R13726 VCC.n8580 VCC.n8579 0.00317857
R13727 VCC.n8585 VCC.n8368 0.00317857
R13728 VCC.n8630 VCC.n8341 0.00317857
R13729 VCC.n8639 VCC.n8638 0.00317857
R13730 VCC.n8656 VCC.n8655 0.00317857
R13731 VCC.n8662 VCC.n8661 0.00317857
R13732 VCC.n8662 VCC.n8313 0.00317857
R13733 VCC.n8581 VCC.n8373 0.00317857
R13734 VCC.n8587 VCC.n8586 0.00317857
R13735 VCC.n8629 VCC.n8342 0.00317857
R13736 VCC.n8657 VCC.n8324 0.00317857
R13737 VCC.n8663 VCC.n8660 0.00317857
R13738 VCC.n215 VCC.n214 0.00228571
R13739 VCC.n222 VCC.n220 0.00228571
R13740 VCC.n162 VCC.n161 0.00228571
R13741 VCC.n278 VCC.n150 0.00228571
R13742 VCC.n352 VCC.n112 0.00228571
R13743 VCC.n478 VCC.n477 0.00228571
R13744 VCC.n489 VCC.n44 0.00228571
R13745 VCC.n501 VCC.n38 0.00228571
R13746 VCC.n522 VCC.n521 0.00228571
R13747 VCC.n502 VCC.n36 0.00228571
R13748 VCC.n767 VCC.n766 0.00228571
R13749 VCC.n774 VCC.n772 0.00228571
R13750 VCC.n714 VCC.n713 0.00228571
R13751 VCC.n830 VCC.n702 0.00228571
R13752 VCC.n904 VCC.n664 0.00228571
R13753 VCC.n1030 VCC.n1029 0.00228571
R13754 VCC.n1041 VCC.n596 0.00228571
R13755 VCC.n1053 VCC.n590 0.00228571
R13756 VCC.n1074 VCC.n1073 0.00228571
R13757 VCC.n1054 VCC.n588 0.00228571
R13758 VCC.n1596 VCC.n1595 0.00228571
R13759 VCC.n1592 VCC.n1588 0.00228571
R13760 VCC.n1605 VCC.n1146 0.00228571
R13761 VCC.n1624 VCC.n1134 0.00228571
R13762 VCC.n1607 VCC.n1606 0.00228571
R13763 VCC.n1461 VCC.n1221 0.00228571
R13764 VCC.n1325 VCC.n1324 0.00228571
R13765 VCC.n1332 VCC.n1330 0.00228571
R13766 VCC.n1272 VCC.n1271 0.00228571
R13767 VCC.n1388 VCC.n1260 0.00228571
R13768 VCC.n1876 VCC.n1875 0.00228571
R13769 VCC.n1883 VCC.n1881 0.00228571
R13770 VCC.n1823 VCC.n1822 0.00228571
R13771 VCC.n1939 VCC.n1811 0.00228571
R13772 VCC.n2013 VCC.n1773 0.00228571
R13773 VCC.n2139 VCC.n2138 0.00228571
R13774 VCC.n2150 VCC.n1705 0.00228571
R13775 VCC.n2162 VCC.n1699 0.00228571
R13776 VCC.n2183 VCC.n2182 0.00228571
R13777 VCC.n2163 VCC.n1697 0.00228571
R13778 VCC.n2705 VCC.n2704 0.00228571
R13779 VCC.n2701 VCC.n2697 0.00228571
R13780 VCC.n2714 VCC.n2255 0.00228571
R13781 VCC.n2733 VCC.n2243 0.00228571
R13782 VCC.n2716 VCC.n2715 0.00228571
R13783 VCC.n2570 VCC.n2330 0.00228571
R13784 VCC.n2434 VCC.n2433 0.00228571
R13785 VCC.n2441 VCC.n2439 0.00228571
R13786 VCC.n2381 VCC.n2380 0.00228571
R13787 VCC.n2497 VCC.n2369 0.00228571
R13788 VCC.n2985 VCC.n2984 0.00228571
R13789 VCC.n2992 VCC.n2990 0.00228571
R13790 VCC.n2932 VCC.n2931 0.00228571
R13791 VCC.n3048 VCC.n2920 0.00228571
R13792 VCC.n3122 VCC.n2882 0.00228571
R13793 VCC.n3248 VCC.n3247 0.00228571
R13794 VCC.n3259 VCC.n2814 0.00228571
R13795 VCC.n3271 VCC.n2808 0.00228571
R13796 VCC.n3292 VCC.n3291 0.00228571
R13797 VCC.n3272 VCC.n2806 0.00228571
R13798 VCC.n3814 VCC.n3813 0.00228571
R13799 VCC.n3810 VCC.n3806 0.00228571
R13800 VCC.n3823 VCC.n3364 0.00228571
R13801 VCC.n3842 VCC.n3352 0.00228571
R13802 VCC.n3825 VCC.n3824 0.00228571
R13803 VCC.n3679 VCC.n3439 0.00228571
R13804 VCC.n3543 VCC.n3542 0.00228571
R13805 VCC.n3550 VCC.n3548 0.00228571
R13806 VCC.n3490 VCC.n3489 0.00228571
R13807 VCC.n3606 VCC.n3478 0.00228571
R13808 VCC.n4094 VCC.n4093 0.00228571
R13809 VCC.n4101 VCC.n4099 0.00228571
R13810 VCC.n4041 VCC.n4040 0.00228571
R13811 VCC.n4157 VCC.n4029 0.00228571
R13812 VCC.n4231 VCC.n3991 0.00228571
R13813 VCC.n4357 VCC.n4356 0.00228571
R13814 VCC.n4368 VCC.n3923 0.00228571
R13815 VCC.n4380 VCC.n3917 0.00228571
R13816 VCC.n4401 VCC.n4400 0.00228571
R13817 VCC.n4381 VCC.n3915 0.00228571
R13818 VCC.n4923 VCC.n4922 0.00228571
R13819 VCC.n4919 VCC.n4915 0.00228571
R13820 VCC.n4932 VCC.n4473 0.00228571
R13821 VCC.n4951 VCC.n4461 0.00228571
R13822 VCC.n4934 VCC.n4933 0.00228571
R13823 VCC.n4788 VCC.n4548 0.00228571
R13824 VCC.n4652 VCC.n4651 0.00228571
R13825 VCC.n4659 VCC.n4657 0.00228571
R13826 VCC.n4599 VCC.n4598 0.00228571
R13827 VCC.n4715 VCC.n4587 0.00228571
R13828 VCC.n5203 VCC.n5202 0.00228571
R13829 VCC.n5210 VCC.n5208 0.00228571
R13830 VCC.n5150 VCC.n5149 0.00228571
R13831 VCC.n5266 VCC.n5138 0.00228571
R13832 VCC.n5340 VCC.n5100 0.00228571
R13833 VCC.n5466 VCC.n5465 0.00228571
R13834 VCC.n5477 VCC.n5032 0.00228571
R13835 VCC.n5489 VCC.n5026 0.00228571
R13836 VCC.n5510 VCC.n5509 0.00228571
R13837 VCC.n5490 VCC.n5024 0.00228571
R13838 VCC.n6031 VCC.n6030 0.00228571
R13839 VCC.n6027 VCC.n6023 0.00228571
R13840 VCC.n6040 VCC.n5581 0.00228571
R13841 VCC.n6059 VCC.n5569 0.00228571
R13842 VCC.n6042 VCC.n6041 0.00228571
R13843 VCC.n5896 VCC.n5656 0.00228571
R13844 VCC.n5760 VCC.n5759 0.00228571
R13845 VCC.n5767 VCC.n5765 0.00228571
R13846 VCC.n5707 VCC.n5706 0.00228571
R13847 VCC.n5823 VCC.n5695 0.00228571
R13848 VCC.n6310 VCC.n6309 0.00228571
R13849 VCC.n6317 VCC.n6315 0.00228571
R13850 VCC.n6257 VCC.n6256 0.00228571
R13851 VCC.n6373 VCC.n6245 0.00228571
R13852 VCC.n6447 VCC.n6207 0.00228571
R13853 VCC.n6573 VCC.n6572 0.00228571
R13854 VCC.n6584 VCC.n6139 0.00228571
R13855 VCC.n6596 VCC.n6133 0.00228571
R13856 VCC.n6617 VCC.n6616 0.00228571
R13857 VCC.n6597 VCC.n6131 0.00228571
R13858 VCC.n7138 VCC.n7137 0.00228571
R13859 VCC.n7134 VCC.n7130 0.00228571
R13860 VCC.n7147 VCC.n6688 0.00228571
R13861 VCC.n7166 VCC.n6676 0.00228571
R13862 VCC.n7149 VCC.n7148 0.00228571
R13863 VCC.n7003 VCC.n6763 0.00228571
R13864 VCC.n6867 VCC.n6866 0.00228571
R13865 VCC.n6874 VCC.n6872 0.00228571
R13866 VCC.n6814 VCC.n6813 0.00228571
R13867 VCC.n6930 VCC.n6802 0.00228571
R13868 VCC.n7417 VCC.n7416 0.00228571
R13869 VCC.n7424 VCC.n7422 0.00228571
R13870 VCC.n7364 VCC.n7363 0.00228571
R13871 VCC.n7480 VCC.n7352 0.00228571
R13872 VCC.n7554 VCC.n7314 0.00228571
R13873 VCC.n7680 VCC.n7679 0.00228571
R13874 VCC.n7691 VCC.n7246 0.00228571
R13875 VCC.n7703 VCC.n7240 0.00228571
R13876 VCC.n7724 VCC.n7723 0.00228571
R13877 VCC.n7704 VCC.n7238 0.00228571
R13878 VCC.n8245 VCC.n8244 0.00228571
R13879 VCC.n8241 VCC.n8237 0.00228571
R13880 VCC.n8254 VCC.n7795 0.00228571
R13881 VCC.n8273 VCC.n7783 0.00228571
R13882 VCC.n8256 VCC.n8255 0.00228571
R13883 VCC.n8110 VCC.n7870 0.00228571
R13884 VCC.n7974 VCC.n7973 0.00228571
R13885 VCC.n7981 VCC.n7979 0.00228571
R13886 VCC.n7921 VCC.n7920 0.00228571
R13887 VCC.n8037 VCC.n7909 0.00228571
R13888 VCC.n8474 VCC.n8421 0.00228571
R13889 VCC.n8600 VCC.n8599 0.00228571
R13890 VCC.n8611 VCC.n8353 0.00228571
R13891 VCC.n8623 VCC.n8347 0.00228571
R13892 VCC.n8644 VCC.n8643 0.00228571
R13893 VCC.n8624 VCC.n8345 0.00228571
R13894 VCC.n217 VCC.n188 0.00217857
R13895 VCC.n218 VCC.n173 0.00217857
R13896 VCC.n307 VCC.n131 0.00217857
R13897 VCC.n308 VCC.n127 0.00217857
R13898 VCC.n317 VCC.n316 0.00217857
R13899 VCC.n346 VCC.n114 0.00217857
R13900 VCC.n442 VCC.n70 0.00217857
R13901 VCC.n443 VCC.n66 0.00217857
R13902 VCC.n460 VCC.n62 0.00217857
R13903 VCC.n461 VCC.n49 0.00217857
R13904 VCC.n536 VCC.n13 0.00217857
R13905 VCC.n537 VCC.n0 0.00217857
R13906 VCC.n769 VCC.n740 0.00217857
R13907 VCC.n770 VCC.n725 0.00217857
R13908 VCC.n859 VCC.n683 0.00217857
R13909 VCC.n860 VCC.n679 0.00217857
R13910 VCC.n869 VCC.n868 0.00217857
R13911 VCC.n898 VCC.n666 0.00217857
R13912 VCC.n994 VCC.n622 0.00217857
R13913 VCC.n995 VCC.n618 0.00217857
R13914 VCC.n1012 VCC.n614 0.00217857
R13915 VCC.n1013 VCC.n601 0.00217857
R13916 VCC.n1088 VCC.n565 0.00217857
R13917 VCC.n1089 VCC.n554 0.00217857
R13918 VCC.n1327 VCC.n1298 0.00217857
R13919 VCC.n1328 VCC.n1283 0.00217857
R13920 VCC.n1417 VCC.n1241 0.00217857
R13921 VCC.n1418 VCC.n1237 0.00217857
R13922 VCC.n1427 VCC.n1426 0.00217857
R13923 VCC.n1455 VCC.n1223 0.00217857
R13924 VCC.n1552 VCC.n1179 0.00217857
R13925 VCC.n1553 VCC.n1175 0.00217857
R13926 VCC.n1571 VCC.n1171 0.00217857
R13927 VCC.n1572 VCC.n1154 0.00217857
R13928 VCC.n1635 VCC.n1126 0.00217857
R13929 VCC.n1636 VCC.n1108 0.00217857
R13930 VCC.n1878 VCC.n1849 0.00217857
R13931 VCC.n1879 VCC.n1834 0.00217857
R13932 VCC.n1968 VCC.n1792 0.00217857
R13933 VCC.n1969 VCC.n1788 0.00217857
R13934 VCC.n1978 VCC.n1977 0.00217857
R13935 VCC.n2007 VCC.n1775 0.00217857
R13936 VCC.n2103 VCC.n1731 0.00217857
R13937 VCC.n2104 VCC.n1727 0.00217857
R13938 VCC.n2121 VCC.n1723 0.00217857
R13939 VCC.n2122 VCC.n1710 0.00217857
R13940 VCC.n2197 VCC.n1674 0.00217857
R13941 VCC.n2198 VCC.n1663 0.00217857
R13942 VCC.n2436 VCC.n2407 0.00217857
R13943 VCC.n2437 VCC.n2392 0.00217857
R13944 VCC.n2526 VCC.n2350 0.00217857
R13945 VCC.n2527 VCC.n2346 0.00217857
R13946 VCC.n2536 VCC.n2535 0.00217857
R13947 VCC.n2564 VCC.n2332 0.00217857
R13948 VCC.n2661 VCC.n2288 0.00217857
R13949 VCC.n2662 VCC.n2284 0.00217857
R13950 VCC.n2680 VCC.n2280 0.00217857
R13951 VCC.n2681 VCC.n2263 0.00217857
R13952 VCC.n2744 VCC.n2235 0.00217857
R13953 VCC.n2745 VCC.n2217 0.00217857
R13954 VCC.n2987 VCC.n2958 0.00217857
R13955 VCC.n2988 VCC.n2943 0.00217857
R13956 VCC.n3077 VCC.n2901 0.00217857
R13957 VCC.n3078 VCC.n2897 0.00217857
R13958 VCC.n3087 VCC.n3086 0.00217857
R13959 VCC.n3116 VCC.n2884 0.00217857
R13960 VCC.n3212 VCC.n2840 0.00217857
R13961 VCC.n3213 VCC.n2836 0.00217857
R13962 VCC.n3230 VCC.n2832 0.00217857
R13963 VCC.n3231 VCC.n2819 0.00217857
R13964 VCC.n3306 VCC.n2783 0.00217857
R13965 VCC.n3307 VCC.n2772 0.00217857
R13966 VCC.n3545 VCC.n3516 0.00217857
R13967 VCC.n3546 VCC.n3501 0.00217857
R13968 VCC.n3635 VCC.n3459 0.00217857
R13969 VCC.n3636 VCC.n3455 0.00217857
R13970 VCC.n3645 VCC.n3644 0.00217857
R13971 VCC.n3673 VCC.n3441 0.00217857
R13972 VCC.n3770 VCC.n3397 0.00217857
R13973 VCC.n3771 VCC.n3393 0.00217857
R13974 VCC.n3789 VCC.n3389 0.00217857
R13975 VCC.n3790 VCC.n3372 0.00217857
R13976 VCC.n3853 VCC.n3344 0.00217857
R13977 VCC.n3854 VCC.n3326 0.00217857
R13978 VCC.n4096 VCC.n4067 0.00217857
R13979 VCC.n4097 VCC.n4052 0.00217857
R13980 VCC.n4186 VCC.n4010 0.00217857
R13981 VCC.n4187 VCC.n4006 0.00217857
R13982 VCC.n4196 VCC.n4195 0.00217857
R13983 VCC.n4225 VCC.n3993 0.00217857
R13984 VCC.n4321 VCC.n3949 0.00217857
R13985 VCC.n4322 VCC.n3945 0.00217857
R13986 VCC.n4339 VCC.n3941 0.00217857
R13987 VCC.n4340 VCC.n3928 0.00217857
R13988 VCC.n4415 VCC.n3892 0.00217857
R13989 VCC.n4416 VCC.n3881 0.00217857
R13990 VCC.n4654 VCC.n4625 0.00217857
R13991 VCC.n4655 VCC.n4610 0.00217857
R13992 VCC.n4744 VCC.n4568 0.00217857
R13993 VCC.n4745 VCC.n4564 0.00217857
R13994 VCC.n4754 VCC.n4753 0.00217857
R13995 VCC.n4782 VCC.n4550 0.00217857
R13996 VCC.n4879 VCC.n4506 0.00217857
R13997 VCC.n4880 VCC.n4502 0.00217857
R13998 VCC.n4898 VCC.n4498 0.00217857
R13999 VCC.n4899 VCC.n4481 0.00217857
R14000 VCC.n4962 VCC.n4453 0.00217857
R14001 VCC.n4963 VCC.n4435 0.00217857
R14002 VCC.n5205 VCC.n5176 0.00217857
R14003 VCC.n5206 VCC.n5161 0.00217857
R14004 VCC.n5295 VCC.n5119 0.00217857
R14005 VCC.n5296 VCC.n5115 0.00217857
R14006 VCC.n5305 VCC.n5304 0.00217857
R14007 VCC.n5334 VCC.n5102 0.00217857
R14008 VCC.n5430 VCC.n5058 0.00217857
R14009 VCC.n5431 VCC.n5054 0.00217857
R14010 VCC.n5448 VCC.n5050 0.00217857
R14011 VCC.n5449 VCC.n5037 0.00217857
R14012 VCC.n5524 VCC.n5001 0.00217857
R14013 VCC.n5525 VCC.n4990 0.00217857
R14014 VCC.n5762 VCC.n5733 0.00217857
R14015 VCC.n5763 VCC.n5718 0.00217857
R14016 VCC.n5852 VCC.n5676 0.00217857
R14017 VCC.n5853 VCC.n5672 0.00217857
R14018 VCC.n5862 VCC.n5861 0.00217857
R14019 VCC.n5890 VCC.n5658 0.00217857
R14020 VCC.n5987 VCC.n5614 0.00217857
R14021 VCC.n5988 VCC.n5610 0.00217857
R14022 VCC.n6006 VCC.n5606 0.00217857
R14023 VCC.n6007 VCC.n5589 0.00217857
R14024 VCC.n6070 VCC.n5561 0.00217857
R14025 VCC.n6071 VCC.n5543 0.00217857
R14026 VCC.n6312 VCC.n6283 0.00217857
R14027 VCC.n6313 VCC.n6268 0.00217857
R14028 VCC.n6402 VCC.n6226 0.00217857
R14029 VCC.n6403 VCC.n6222 0.00217857
R14030 VCC.n6412 VCC.n6411 0.00217857
R14031 VCC.n6441 VCC.n6209 0.00217857
R14032 VCC.n6537 VCC.n6165 0.00217857
R14033 VCC.n6538 VCC.n6161 0.00217857
R14034 VCC.n6555 VCC.n6157 0.00217857
R14035 VCC.n6556 VCC.n6144 0.00217857
R14036 VCC.n6631 VCC.n6108 0.00217857
R14037 VCC.n6632 VCC.n6097 0.00217857
R14038 VCC.n6869 VCC.n6840 0.00217857
R14039 VCC.n6870 VCC.n6825 0.00217857
R14040 VCC.n6959 VCC.n6783 0.00217857
R14041 VCC.n6960 VCC.n6779 0.00217857
R14042 VCC.n6969 VCC.n6968 0.00217857
R14043 VCC.n6997 VCC.n6765 0.00217857
R14044 VCC.n7094 VCC.n6721 0.00217857
R14045 VCC.n7095 VCC.n6717 0.00217857
R14046 VCC.n7113 VCC.n6713 0.00217857
R14047 VCC.n7114 VCC.n6696 0.00217857
R14048 VCC.n7177 VCC.n6668 0.00217857
R14049 VCC.n7178 VCC.n6650 0.00217857
R14050 VCC.n7419 VCC.n7390 0.00217857
R14051 VCC.n7420 VCC.n7375 0.00217857
R14052 VCC.n7509 VCC.n7333 0.00217857
R14053 VCC.n7510 VCC.n7329 0.00217857
R14054 VCC.n7519 VCC.n7518 0.00217857
R14055 VCC.n7548 VCC.n7316 0.00217857
R14056 VCC.n7644 VCC.n7272 0.00217857
R14057 VCC.n7645 VCC.n7268 0.00217857
R14058 VCC.n7662 VCC.n7264 0.00217857
R14059 VCC.n7663 VCC.n7251 0.00217857
R14060 VCC.n7738 VCC.n7215 0.00217857
R14061 VCC.n7739 VCC.n7204 0.00217857
R14062 VCC.n7976 VCC.n7947 0.00217857
R14063 VCC.n7977 VCC.n7932 0.00217857
R14064 VCC.n8066 VCC.n7890 0.00217857
R14065 VCC.n8067 VCC.n7886 0.00217857
R14066 VCC.n8076 VCC.n8075 0.00217857
R14067 VCC.n8104 VCC.n7872 0.00217857
R14068 VCC.n8201 VCC.n7828 0.00217857
R14069 VCC.n8202 VCC.n7824 0.00217857
R14070 VCC.n8220 VCC.n7820 0.00217857
R14071 VCC.n8221 VCC.n7803 0.00217857
R14072 VCC.n8284 VCC.n7775 0.00217857
R14073 VCC.n8285 VCC.n7757 0.00217857
R14074 VCC.n8439 VCC.n8438 0.00217857
R14075 VCC.n8468 VCC.n8423 0.00217857
R14076 VCC.n8564 VCC.n8379 0.00217857
R14077 VCC.n8565 VCC.n8375 0.00217857
R14078 VCC.n8582 VCC.n8371 0.00217857
R14079 VCC.n8583 VCC.n8358 0.00217857
R14080 VCC.n8658 VCC.n8322 0.00217857
R14081 VCC.n8659 VCC.n8311 0.00217857
R14082 VCC.n214 VCC.n193 0.00139286
R14083 VCC.n237 VCC.n236 0.00139286
R14084 VCC.n254 VCC.n253 0.00139286
R14085 VCC.n294 VCC.n129 0.00139286
R14086 VCC.n252 VCC.n167 0.00139286
R14087 VCC.n350 VCC.n104 0.00139286
R14088 VCC.n405 VCC.n90 0.00139286
R14089 VCC.n532 VCC.n19 0.00139286
R14090 VCC.n543 VCC.n8 0.00139286
R14091 VCC.n766 VCC.n745 0.00139286
R14092 VCC.n789 VCC.n788 0.00139286
R14093 VCC.n806 VCC.n805 0.00139286
R14094 VCC.n846 VCC.n681 0.00139286
R14095 VCC.n804 VCC.n719 0.00139286
R14096 VCC.n902 VCC.n656 0.00139286
R14097 VCC.n957 VCC.n642 0.00139286
R14098 VCC.n1084 VCC.n571 0.00139286
R14099 VCC.n1097 VCC.n562 0.00139286
R14100 VCC.n1647 VCC.n1646 0.00139286
R14101 VCC.n1125 VCC.n1122 0.00139286
R14102 VCC.n1459 VCC.n1213 0.00139286
R14103 VCC.n1514 VCC.n1199 0.00139286
R14104 VCC.n1324 VCC.n1303 0.00139286
R14105 VCC.n1347 VCC.n1346 0.00139286
R14106 VCC.n1364 VCC.n1363 0.00139286
R14107 VCC.n1404 VCC.n1239 0.00139286
R14108 VCC.n1362 VCC.n1277 0.00139286
R14109 VCC.n1875 VCC.n1854 0.00139286
R14110 VCC.n1898 VCC.n1897 0.00139286
R14111 VCC.n1915 VCC.n1914 0.00139286
R14112 VCC.n1955 VCC.n1790 0.00139286
R14113 VCC.n1913 VCC.n1828 0.00139286
R14114 VCC.n2011 VCC.n1765 0.00139286
R14115 VCC.n2066 VCC.n1751 0.00139286
R14116 VCC.n2193 VCC.n1680 0.00139286
R14117 VCC.n2206 VCC.n1671 0.00139286
R14118 VCC.n2756 VCC.n2755 0.00139286
R14119 VCC.n2234 VCC.n2231 0.00139286
R14120 VCC.n2568 VCC.n2322 0.00139286
R14121 VCC.n2623 VCC.n2308 0.00139286
R14122 VCC.n2433 VCC.n2412 0.00139286
R14123 VCC.n2456 VCC.n2455 0.00139286
R14124 VCC.n2473 VCC.n2472 0.00139286
R14125 VCC.n2513 VCC.n2348 0.00139286
R14126 VCC.n2471 VCC.n2386 0.00139286
R14127 VCC.n2984 VCC.n2963 0.00139286
R14128 VCC.n3007 VCC.n3006 0.00139286
R14129 VCC.n3024 VCC.n3023 0.00139286
R14130 VCC.n3064 VCC.n2899 0.00139286
R14131 VCC.n3022 VCC.n2937 0.00139286
R14132 VCC.n3120 VCC.n2874 0.00139286
R14133 VCC.n3175 VCC.n2860 0.00139286
R14134 VCC.n3302 VCC.n2789 0.00139286
R14135 VCC.n3315 VCC.n2780 0.00139286
R14136 VCC.n3865 VCC.n3864 0.00139286
R14137 VCC.n3343 VCC.n3340 0.00139286
R14138 VCC.n3677 VCC.n3431 0.00139286
R14139 VCC.n3732 VCC.n3417 0.00139286
R14140 VCC.n3542 VCC.n3521 0.00139286
R14141 VCC.n3565 VCC.n3564 0.00139286
R14142 VCC.n3582 VCC.n3581 0.00139286
R14143 VCC.n3622 VCC.n3457 0.00139286
R14144 VCC.n3580 VCC.n3495 0.00139286
R14145 VCC.n4093 VCC.n4072 0.00139286
R14146 VCC.n4116 VCC.n4115 0.00139286
R14147 VCC.n4133 VCC.n4132 0.00139286
R14148 VCC.n4173 VCC.n4008 0.00139286
R14149 VCC.n4131 VCC.n4046 0.00139286
R14150 VCC.n4229 VCC.n3983 0.00139286
R14151 VCC.n4284 VCC.n3969 0.00139286
R14152 VCC.n4411 VCC.n3898 0.00139286
R14153 VCC.n4424 VCC.n3889 0.00139286
R14154 VCC.n4974 VCC.n4973 0.00139286
R14155 VCC.n4452 VCC.n4449 0.00139286
R14156 VCC.n4786 VCC.n4540 0.00139286
R14157 VCC.n4841 VCC.n4526 0.00139286
R14158 VCC.n4651 VCC.n4630 0.00139286
R14159 VCC.n4674 VCC.n4673 0.00139286
R14160 VCC.n4691 VCC.n4690 0.00139286
R14161 VCC.n4731 VCC.n4566 0.00139286
R14162 VCC.n4689 VCC.n4604 0.00139286
R14163 VCC.n5202 VCC.n5181 0.00139286
R14164 VCC.n5225 VCC.n5224 0.00139286
R14165 VCC.n5242 VCC.n5241 0.00139286
R14166 VCC.n5282 VCC.n5117 0.00139286
R14167 VCC.n5240 VCC.n5155 0.00139286
R14168 VCC.n5338 VCC.n5092 0.00139286
R14169 VCC.n5393 VCC.n5078 0.00139286
R14170 VCC.n5520 VCC.n5007 0.00139286
R14171 VCC.n5533 VCC.n4998 0.00139286
R14172 VCC.n6082 VCC.n6081 0.00139286
R14173 VCC.n5560 VCC.n5557 0.00139286
R14174 VCC.n5894 VCC.n5648 0.00139286
R14175 VCC.n5949 VCC.n5634 0.00139286
R14176 VCC.n5759 VCC.n5738 0.00139286
R14177 VCC.n5782 VCC.n5781 0.00139286
R14178 VCC.n5799 VCC.n5798 0.00139286
R14179 VCC.n5839 VCC.n5674 0.00139286
R14180 VCC.n5797 VCC.n5712 0.00139286
R14181 VCC.n6309 VCC.n6288 0.00139286
R14182 VCC.n6332 VCC.n6331 0.00139286
R14183 VCC.n6349 VCC.n6348 0.00139286
R14184 VCC.n6389 VCC.n6224 0.00139286
R14185 VCC.n6347 VCC.n6262 0.00139286
R14186 VCC.n6445 VCC.n6199 0.00139286
R14187 VCC.n6500 VCC.n6185 0.00139286
R14188 VCC.n6627 VCC.n6114 0.00139286
R14189 VCC.n6640 VCC.n6105 0.00139286
R14190 VCC.n7189 VCC.n7188 0.00139286
R14191 VCC.n6667 VCC.n6664 0.00139286
R14192 VCC.n7001 VCC.n6755 0.00139286
R14193 VCC.n7056 VCC.n6741 0.00139286
R14194 VCC.n6866 VCC.n6845 0.00139286
R14195 VCC.n6889 VCC.n6888 0.00139286
R14196 VCC.n6906 VCC.n6905 0.00139286
R14197 VCC.n6946 VCC.n6781 0.00139286
R14198 VCC.n6904 VCC.n6819 0.00139286
R14199 VCC.n7416 VCC.n7395 0.00139286
R14200 VCC.n7439 VCC.n7438 0.00139286
R14201 VCC.n7456 VCC.n7455 0.00139286
R14202 VCC.n7496 VCC.n7331 0.00139286
R14203 VCC.n7454 VCC.n7369 0.00139286
R14204 VCC.n7552 VCC.n7306 0.00139286
R14205 VCC.n7607 VCC.n7292 0.00139286
R14206 VCC.n7734 VCC.n7221 0.00139286
R14207 VCC.n7747 VCC.n7212 0.00139286
R14208 VCC.n8296 VCC.n8295 0.00139286
R14209 VCC.n7774 VCC.n7771 0.00139286
R14210 VCC.n8108 VCC.n7862 0.00139286
R14211 VCC.n8163 VCC.n7848 0.00139286
R14212 VCC.n7973 VCC.n7952 0.00139286
R14213 VCC.n7996 VCC.n7995 0.00139286
R14214 VCC.n8013 VCC.n8012 0.00139286
R14215 VCC.n8053 VCC.n7888 0.00139286
R14216 VCC.n8011 VCC.n7926 0.00139286
R14217 VCC.n8472 VCC.n8413 0.00139286
R14218 VCC.n8527 VCC.n8399 0.00139286
R14219 VCC.n8654 VCC.n8328 0.00139286
R14220 VCC.n8667 VCC.n8319 0.00139286
R14221 VCC.n8677 VCC.n8310 0.00054824
R14222 VCC.n8679 VCC.n7203 0.00054824
R14223 VCC.n8681 VCC.n6096 0.00054824
R14224 VCC.n4989 VCC.n4988 0.00054824
R14225 VCC.n3880 VCC.n3879 0.00054824
R14226 VCC.n2771 VCC.n2770 0.00054824
R14227 VCC.n1662 VCC.n1661 0.00054824
R14228 VSS.n9340 VSS.n24 106073
R14229 VSS.n1003 VSS.n24 54262.5
R14230 VSS.n9340 VSS.n16 12274.8
R14231 VSS.n9340 VSS.n17 12232.2
R14232 VSS.n9340 VSS.n15 12232.2
R14233 VSS.n9341 VSS.n9340 12232.2
R14234 VSS.n9340 VSS.n18 12232.2
R14235 VSS.n9340 VSS.n14 12232.2
R14236 VSS.n9340 VSS.n19 12232.2
R14237 VSS.n9340 VSS.n13 12232.2
R14238 VSS.n9340 VSS.n20 12232.2
R14239 VSS.n9340 VSS.n12 12232.2
R14240 VSS.n9340 VSS.n21 12232.2
R14241 VSS.n9340 VSS.n11 12232.2
R14242 VSS.n9340 VSS.n22 12232.2
R14243 VSS.n9340 VSS.n23 12232.2
R14244 VSS.n9340 VSS.n10 12232.2
R14245 VSS.n9340 VSS.n9339 12232.2
R14246 VSS.n1004 VSS.n1003 6909.46
R14247 VSS.n8535 VSS.n1004 6909.46
R14248 VSS.n8535 VSS.n8534 6909.46
R14249 VSS.n8534 VSS.n8533 6909.46
R14250 VSS.n8533 VSS.n8532 6909.46
R14251 VSS.n8532 VSS.n8531 6909.46
R14252 VSS.n8531 VSS.n8530 6909.46
R14253 VSS.n8530 VSS.n8529 6909.46
R14254 VSS.n8529 VSS.n8528 6909.46
R14255 VSS.n8528 VSS.n8527 6909.46
R14256 VSS.n8527 VSS.n8526 6909.46
R14257 VSS.n8526 VSS.n8525 6909.46
R14258 VSS.n8525 VSS.n8524 6909.46
R14259 VSS.n8524 VSS.t85 6273.77
R14260 VSS.n7605 VSS.t49 4305.17
R14261 VSS.n8197 VSS.t300 4305.17
R14262 VSS.n1664 VSS.t312 4305.17
R14263 VSS.n2256 VSS.t91 4305.17
R14264 VSS.n3807 VSS.t246 4305.17
R14265 VSS.n4399 VSS.t17 4305.17
R14266 VSS.n4991 VSS.t122 4305.17
R14267 VSS.n5583 VSS.t275 4305.17
R14268 VSS.n6175 VSS.t105 4305.17
R14269 VSS.n6767 VSS.t283 4305.17
R14270 VSS.n7000 VSS.t204 4305.17
R14271 VSS.n3215 VSS.t57 4305.17
R14272 VSS.n9175 VSS.t141 4305.17
R14273 VSS.n9001 VSS.t6 4305.17
R14274 VSS.n819 VSS.t293 4305.17
R14275 VSS.n8477 VSS.n7055 3531.03
R14276 VSS.n7055 VSS.n7054 3531.03
R14277 VSS.n7054 VSS.n7053 3531.03
R14278 VSS.n7053 VSS.n7052 3531.03
R14279 VSS.n7052 VSS.n7051 3531.03
R14280 VSS.n7051 VSS.n7050 3531.03
R14281 VSS.n7050 VSS.n7049 3531.03
R14282 VSS.n7049 VSS.n7048 3531.03
R14283 VSS.n7048 VSS.n7047 3531.03
R14284 VSS.n7047 VSS.n191 3531.03
R14285 VSS.n9049 VSS.n24 3531.03
R14286 VSS.n9049 VSS.n9048 3531.03
R14287 VSS.n9048 VSS.n191 3531.03
R14288 VSS.n8477 VSS.n8476 3531.03
R14289 VSS.n7055 VSS.t163 3054.19
R14290 VSS.n7054 VSS.t23 3054.19
R14291 VSS.n7053 VSS.t198 3054.19
R14292 VSS.n7052 VSS.t238 3054.19
R14293 VSS.n7051 VSS.t166 3054.19
R14294 VSS.n7050 VSS.t208 3054.19
R14295 VSS.n7049 VSS.t185 3054.19
R14296 VSS.n7048 VSS.t297 3054.19
R14297 VSS.n7047 VSS.t201 3054.19
R14298 VSS.t58 VSS.n191 3054.19
R14299 VSS.n9049 VSS.t109 3054.19
R14300 VSS.n9048 VSS.t145 3054.19
R14301 VSS.t254 VSS.n24 3054.19
R14302 VSS.n8477 VSS.t287 3054.19
R14303 VSS.n8428 VSS.t133 2804.58
R14304 VSS.n8427 VSS.t134 2770.93
R14305 VSS.n8429 VSS.n8428 2671.38
R14306 VSS.t134 VSS.t74 2603.46
R14307 VSS.n9048 VSS.n192 2588.02
R14308 VSS.n7055 VSS.n1138 2588.02
R14309 VSS.n7054 VSS.n1711 2588.02
R14310 VSS.n7053 VSS.n2303 2588.02
R14311 VSS.n7052 VSS.n2304 2588.02
R14312 VSS.n7051 VSS.n2305 2588.02
R14313 VSS.n7050 VSS.n2306 2588.02
R14314 VSS.n7049 VSS.n2307 2588.02
R14315 VSS.n7048 VSS.n2308 2588.02
R14316 VSS.n7047 VSS.n2309 2588.02
R14317 VSS.n3090 VSS.n191 2588.02
R14318 VSS.n9050 VSS.n9049 2588.02
R14319 VSS.n957 VSS.n24 2588.02
R14320 VSS.n8478 VSS.n8477 2588.02
R14321 VSS.n7606 VSS.n7605 2406.66
R14322 VSS.n8198 VSS.n8197 2406.66
R14323 VSS.n1665 VSS.n1664 2406.66
R14324 VSS.n2257 VSS.n2256 2406.66
R14325 VSS.n3808 VSS.n3807 2406.66
R14326 VSS.n4400 VSS.n4399 2406.66
R14327 VSS.n4992 VSS.n4991 2406.66
R14328 VSS.n5584 VSS.n5583 2406.66
R14329 VSS.n6176 VSS.n6175 2406.66
R14330 VSS.n6768 VSS.n6767 2406.66
R14331 VSS.n7001 VSS.n7000 2406.66
R14332 VSS.n3216 VSS.n3215 2406.66
R14333 VSS.n9176 VSS.n9175 2406.66
R14334 VSS.n9002 VSS.n9001 2406.66
R14335 VSS.n820 VSS.n819 2406.66
R14336 VSS.t108 VSS.n8474 2349.66
R14337 VSS.t162 VSS.t108 2304.76
R14338 VSS.n7480 VSS.t124 1937.11
R14339 VSS.n7894 VSS.t284 1937.11
R14340 VSS.t70 VSS.n1710 1937.11
R14341 VSS.t138 VSS.n2302 1937.11
R14342 VSS.n3504 VSS.t174 1937.11
R14343 VSS.n4096 VSS.t247 1937.11
R14344 VSS.n4688 VSS.t169 1937.11
R14345 VSS.n5280 VSS.t129 1937.11
R14346 VSS.n5872 VSS.t95 1937.11
R14347 VSS.n6464 VSS.t190 1937.11
R14348 VSS.t235 VSS.n7046 1937.11
R14349 VSS.n2911 VSS.t153 1937.11
R14350 VSS.t261 VSS.n190 1937.11
R14351 VSS.t26 VSS.n9047 1937.11
R14352 VSS.n544 VSS.t220 1937.11
R14353 VSS.n8536 VSS.t42 1930.89
R14354 VSS.n1218 VSS.t214 1930.89
R14355 VSS.n1791 VSS.t242 1930.89
R14356 VSS.n3585 VSS.t90 1930.89
R14357 VSS.n4177 VSS.t179 1930.89
R14358 VSS.n4769 VSS.t264 1930.89
R14359 VSS.n5361 VSS.t211 1930.89
R14360 VSS.n5953 VSS.t184 1930.89
R14361 VSS.n6545 VSS.t130 1930.89
R14362 VSS.n2389 VSS.t315 1930.89
R14363 VSS.n2986 VSS.t135 1930.89
R14364 VSS.t156 VSS.n437 1930.89
R14365 VSS.t159 VSS.n1002 1930.89
R14366 VSS.t84 VSS.n8523 1930.89
R14367 VSS.n7605 VSS.n7604 1896.55
R14368 VSS.n8197 VSS.n8196 1896.55
R14369 VSS.n1664 VSS.n1663 1896.55
R14370 VSS.n2256 VSS.n2255 1896.55
R14371 VSS.n3807 VSS.n3806 1896.55
R14372 VSS.n4399 VSS.n4398 1896.55
R14373 VSS.n4991 VSS.n4990 1896.55
R14374 VSS.n5583 VSS.n5582 1896.55
R14375 VSS.n6175 VSS.n6174 1896.55
R14376 VSS.n6767 VSS.n6766 1896.55
R14377 VSS.n7000 VSS.n6999 1896.55
R14378 VSS.n3215 VSS.n3214 1896.55
R14379 VSS.n9175 VSS.n9174 1896.55
R14380 VSS.n9001 VSS.n9000 1896.55
R14381 VSS.n819 VSS.n818 1896.55
R14382 VSS.t284 VSS.t223 1892.74
R14383 VSS.t42 VSS.t7 1892.74
R14384 VSS.t214 VSS.t51 1892.74
R14385 VSS.t163 VSS.t70 1892.74
R14386 VSS.t242 VSS.t67 1892.74
R14387 VSS.t23 VSS.t138 1892.74
R14388 VSS.t90 VSS.t63 1892.74
R14389 VSS.t174 VSS.t198 1892.74
R14390 VSS.t179 VSS.t148 1892.74
R14391 VSS.t247 VSS.t238 1892.74
R14392 VSS.t264 VSS.t64 1892.74
R14393 VSS.t169 VSS.t166 1892.74
R14394 VSS.t211 VSS.t81 1892.74
R14395 VSS.t129 VSS.t208 1892.74
R14396 VSS.t184 VSS.t294 1892.74
R14397 VSS.t95 VSS.t185 1892.74
R14398 VSS.t130 VSS.t191 1892.74
R14399 VSS.t190 VSS.t297 1892.74
R14400 VSS.t315 VSS.t232 1892.74
R14401 VSS.t201 VSS.t235 1892.74
R14402 VSS.t135 VSS.t215 1892.74
R14403 VSS.t153 VSS.t58 1892.74
R14404 VSS.t308 VSS.t156 1892.74
R14405 VSS.t109 VSS.t261 1892.74
R14406 VSS.t145 VSS.t26 1892.74
R14407 VSS.t267 VSS.t159 1892.74
R14408 VSS.t220 VSS.t254 1892.74
R14409 VSS.t18 VSS.t84 1892.74
R14410 VSS.t124 VSS.t287 1892.74
R14411 VSS.n7604 VSS.t50 1791.5
R14412 VSS.n8196 VSS.t303 1791.5
R14413 VSS.n1663 VSS.t311 1791.5
R14414 VSS.n2255 VSS.t94 1791.5
R14415 VSS.n3806 VSS.t243 1791.5
R14416 VSS.n4398 VSS.t14 1791.5
R14417 VSS.n4990 VSS.t123 1791.5
R14418 VSS.n5582 VSS.t274 1791.5
R14419 VSS.n6174 VSS.t104 1791.5
R14420 VSS.n6766 VSS.t280 1791.5
R14421 VSS.n6999 VSS.t207 1791.5
R14422 VSS.n3214 VSS.t54 1791.5
R14423 VSS.n9174 VSS.t144 1791.5
R14424 VSS.n9000 VSS.t3 1791.5
R14425 VSS.n818 VSS.t292 1791.5
R14426 VSS.t50 VSS.t77 1683.22
R14427 VSS.t303 VSS.t224 1683.22
R14428 VSS.t311 VSS.t112 1683.22
R14429 VSS.t94 VSS.t175 1683.22
R14430 VSS.t243 VSS.t250 1683.22
R14431 VSS.t14 VSS.t229 1683.22
R14432 VSS.t123 VSS.t116 1683.22
R14433 VSS.t274 VSS.t304 1683.22
R14434 VSS.t104 VSS.t276 1683.22
R14435 VSS.t280 VSS.t101 1683.22
R14436 VSS.t207 VSS.t194 1683.22
R14437 VSS.t54 VSS.t30 1683.22
R14438 VSS.t144 VSS.t38 1683.22
R14439 VSS.t3 VSS.t37 1683.22
R14440 VSS.t292 VSS.t260 1683.22
R14441 VSS.t74 VSS.n8426 1560.55
R14442 VSS.n8475 VSS.t162 1331.97
R14443 VSS.n8475 VSS.t223 1093.85
R14444 VSS.t7 VSS.n8535 1093.85
R14445 VSS.n8525 VSS.t51 1093.85
R14446 VSS.n8526 VSS.t67 1093.85
R14447 VSS.n8527 VSS.t63 1093.85
R14448 VSS.n8528 VSS.t148 1093.85
R14449 VSS.n8529 VSS.t64 1093.85
R14450 VSS.n8530 VSS.t81 1093.85
R14451 VSS.n8531 VSS.t294 1093.85
R14452 VSS.n8532 VSS.t191 1093.85
R14453 VSS.n8533 VSS.t232 1093.85
R14454 VSS.n8534 VSS.t215 1093.85
R14455 VSS.n1004 VSS.t308 1093.85
R14456 VSS.n1003 VSS.t267 1093.85
R14457 VSS.n8524 VSS.t18 1093.85
R14458 VSS.t77 VSS.n7603 1045.79
R14459 VSS.t224 VSS.n8195 1045.79
R14460 VSS.t112 VSS.n1662 1045.79
R14461 VSS.t175 VSS.n2254 1045.79
R14462 VSS.t250 VSS.n3805 1045.79
R14463 VSS.t229 VSS.n4397 1045.79
R14464 VSS.t116 VSS.n4989 1045.79
R14465 VSS.t304 VSS.n5581 1045.79
R14466 VSS.t276 VSS.n6173 1045.79
R14467 VSS.t101 VSS.n6765 1045.79
R14468 VSS.t194 VSS.n6998 1045.79
R14469 VSS.t30 VSS.n3213 1045.79
R14470 VSS.t38 VSS.n9173 1045.79
R14471 VSS.t37 VSS.n8999 1045.79
R14472 VSS.t260 VSS.n817 1045.79
R14473 VSS.n8476 VSS.n7056 1017.62
R14474 VSS.n8476 VSS.n8475 772.908
R14475 VSS.n7975 VSS.t241 758.37
R14476 VSS.t241 VSS.t85 746.255
R14477 VSS.n7603 VSS.n7602 590.341
R14478 VSS.n7344 VSS.n17 590.341
R14479 VSS.n8195 VSS.n8194 590.341
R14480 VSS.n7758 VSS.n15 590.341
R14481 VSS.n8999 VSS.n8998 590.341
R14482 VSS.n8899 VSS.n10 590.341
R14483 VSS.n1662 VSS.n1661 590.341
R14484 VSS.n9341 VSS.n6 590.341
R14485 VSS.n2254 VSS.n2253 590.341
R14486 VSS.n2158 VSS.n18 590.341
R14487 VSS.n3805 VSS.n3804 590.341
R14488 VSS.n3369 VSS.n14 590.341
R14489 VSS.n4397 VSS.n4396 590.341
R14490 VSS.n3961 VSS.n19 590.341
R14491 VSS.n4989 VSS.n4988 590.341
R14492 VSS.n4553 VSS.n13 590.341
R14493 VSS.n5581 VSS.n5580 590.341
R14494 VSS.n5145 VSS.n20 590.341
R14495 VSS.n6173 VSS.n6172 590.341
R14496 VSS.n5737 VSS.n12 590.341
R14497 VSS.n6765 VSS.n6764 590.341
R14498 VSS.n6329 VSS.n21 590.341
R14499 VSS.n6998 VSS.n6997 590.341
R14500 VSS.n2756 VSS.n11 590.341
R14501 VSS.n3213 VSS.n3212 590.341
R14502 VSS.n2776 VSS.n22 590.341
R14503 VSS.n9173 VSS.n9172 590.341
R14504 VSS.n43 VSS.n23 590.341
R14505 VSS.n817 VSS.n816 590.341
R14506 VSS.n9339 VSS.n9338 590.341
R14507 VSS.n8426 VSS.n8425 590.341
R14508 VSS.n7324 VSS.n16 590.341
R14509 VSS.n7479 VSS.n7468 585
R14510 VSS.n7481 VSS.n7468 585
R14511 VSS.n7467 VSS.n7466 585
R14512 VSS.n7508 VSS.n7467 585
R14513 VSS.n7528 VSS.n7527 585
R14514 VSS.n7529 VSS.n7528 585
R14515 VSS.n7434 VSS.n7433 585
R14516 VSS.n7433 VSS.n7432 585
R14517 VSS.n7563 VSS.n7562 585
R14518 VSS.n7562 VSS.t71 585
R14519 VSS.n7581 VSS.n7580 585
R14520 VSS.n7582 VSS.n7581 585
R14521 VSS.n7452 VSS.n7450 585
R14522 VSS.n7531 VSS.n7452 585
R14523 VSS.n7451 VSS.n7449 585
R14524 VSS.n7530 VSS.n7451 585
R14525 VSS.n7511 VSS.n7510 585
R14526 VSS.n7510 VSS.n7509 585
R14527 VSS.n7431 VSS.n7430 585
R14528 VSS.n7561 VSS.n7431 585
R14529 VSS.n7416 VSS.n7415 585
R14530 VSS.n7583 VSS.n7416 585
R14531 VSS.n7484 VSS.n7483 585
R14532 VSS.n7483 VSS.n7482 585
R14533 VSS.n7594 VSS.n7590 585
R14534 VSS.n7598 VSS.n7590 585
R14535 VSS.n7642 VSS.n7641 585
R14536 VSS.n7643 VSS.n7642 585
R14537 VSS.n7393 VSS.n7391 585
R14538 VSS.n7645 VSS.n7393 585
R14539 VSS.n7698 VSS.n7697 585
R14540 VSS.n7697 VSS.n7696 585
R14541 VSS.n7359 VSS.n7358 585
R14542 VSS.t313 VSS.n7359 585
R14543 VSS.n7739 VSS.n7738 585
R14544 VSS.n7740 VSS.n7739 585
R14545 VSS.n7737 VSS.n7345 585
R14546 VSS.n7741 VSS.n7345 585
R14547 VSS.n7718 VSS.n7717 585
R14548 VSS.n7717 VSS.n7716 585
R14549 VSS.n7699 VSS.n7361 585
R14550 VSS.n7361 VSS.n7360 585
R14551 VSS.n7396 VSS.n7395 585
R14552 VSS.n7395 VSS.n7394 585
R14553 VSS.n7648 VSS.n7647 585
R14554 VSS.n7647 VSS.n7646 585
R14555 VSS.n7742 VSS.n7346 585
R14556 VSS.n7585 VSS.n7584 585
R14557 VSS.n7596 VSS.n7595 585
R14558 VSS.n7597 VSS.n7596 585
R14559 VSS.n7893 VSS.n7882 585
R14560 VSS.n7895 VSS.n7882 585
R14561 VSS.n7881 VSS.n7880 585
R14562 VSS.n8100 VSS.n7881 585
R14563 VSS.n8120 VSS.n8119 585
R14564 VSS.n8121 VSS.n8120 585
R14565 VSS.n7848 VSS.n7847 585
R14566 VSS.n7847 VSS.n7846 585
R14567 VSS.n8155 VSS.n8154 585
R14568 VSS.n8154 VSS.t125 585
R14569 VSS.n8173 VSS.n8172 585
R14570 VSS.n8174 VSS.n8173 585
R14571 VSS.n7866 VSS.n7864 585
R14572 VSS.n8123 VSS.n7866 585
R14573 VSS.n7865 VSS.n7863 585
R14574 VSS.n8122 VSS.n7865 585
R14575 VSS.n8103 VSS.n8102 585
R14576 VSS.n8102 VSS.n8101 585
R14577 VSS.n7845 VSS.n7844 585
R14578 VSS.n8153 VSS.n7845 585
R14579 VSS.n7830 VSS.n7829 585
R14580 VSS.n8175 VSS.n7830 585
R14581 VSS.n7898 VSS.n7897 585
R14582 VSS.n7897 VSS.n7896 585
R14583 VSS.n8186 VSS.n8182 585
R14584 VSS.n8190 VSS.n8182 585
R14585 VSS.n8234 VSS.n8233 585
R14586 VSS.n8235 VSS.n8234 585
R14587 VSS.n7807 VSS.n7805 585
R14588 VSS.n8237 VSS.n7807 585
R14589 VSS.n8290 VSS.n8289 585
R14590 VSS.n8289 VSS.n8288 585
R14591 VSS.n7773 VSS.n7772 585
R14592 VSS.t47 VSS.n7773 585
R14593 VSS.n8331 VSS.n8330 585
R14594 VSS.n8332 VSS.n8331 585
R14595 VSS.n8329 VSS.n7759 585
R14596 VSS.n8333 VSS.n7759 585
R14597 VSS.n8310 VSS.n8309 585
R14598 VSS.n8309 VSS.n8308 585
R14599 VSS.n8291 VSS.n7775 585
R14600 VSS.n7775 VSS.n7774 585
R14601 VSS.n7810 VSS.n7809 585
R14602 VSS.n7809 VSS.n7808 585
R14603 VSS.n8240 VSS.n8239 585
R14604 VSS.n8239 VSS.n8238 585
R14605 VSS.n8334 VSS.n7760 585
R14606 VSS.n8177 VSS.n8176 585
R14607 VSS.n8188 VSS.n8187 585
R14608 VSS.n8189 VSS.n8188 585
R14609 VSS.n271 VSS.n270 585
R14610 VSS.n8537 VSS.n271 585
R14611 VSS.n8563 VSS.n8562 585
R14612 VSS.n8564 VSS.n8563 585
R14613 VSS.n256 VSS.n254 585
R14614 VSS.n8568 VSS.n256 585
R14615 VSS.n226 VSS.n224 585
R14616 VSS.n8599 VSS.n226 585
R14617 VSS.n204 VSS.n203 585
R14618 VSS.n8600 VSS.n203 585
R14619 VSS.n212 VSS.n202 585
R14620 VSS.n8631 VSS.n202 585
R14621 VSS.n8597 VSS.n8596 585
R14622 VSS.n8598 VSS.n8597 585
R14623 VSS.n8566 VSS.n236 585
R14624 VSS.n8567 VSS.n8566 585
R14625 VSS.n8561 VSS.n255 585
R14626 VSS.n8565 VSS.n255 585
R14627 VSS.n233 VSS.n232 585
R14628 VSS.n8601 VSS.n233 585
R14629 VSS.n8633 VSS.n201 585
R14630 VSS.n8633 VSS.n8632 585
R14631 VSS.n8540 VSS.n8539 585
R14632 VSS.n8539 VSS.n8538 585
R14633 VSS.n1383 VSS.n1382 585
R14634 VSS.n1382 VSS.n1381 585
R14635 VSS.n1406 VSS.n1405 585
R14636 VSS.n1407 VSS.n1406 585
R14637 VSS.n1412 VSS.n1375 585
R14638 VSS.n1375 VSS.n1374 585
R14639 VSS.n1420 VSS.n1371 585
R14640 VSS.n1371 VSS.n1370 585
R14641 VSS.n1435 VSS.n1434 585
R14642 VSS.n1434 VSS.t139 585
R14643 VSS.n1447 VSS.n1446 585
R14644 VSS.n1448 VSS.n1447 585
R14645 VSS.n1419 VSS.n1418 585
R14646 VSS.n1418 VSS.n1417 585
R14647 VSS.n1414 VSS.n1413 585
R14648 VSS.n1415 VSS.n1414 585
R14649 VSS.n1404 VSS.n1378 585
R14650 VSS.n1408 VSS.n1378 585
R14651 VSS.n1369 VSS.n1368 585
R14652 VSS.n1433 VSS.n1369 585
R14653 VSS.n1360 VSS.n1359 585
R14654 VSS.n1449 VSS.n1360 585
R14655 VSS.n1141 VSS.n1140 585
R14656 VSS.n1140 VSS.n1139 585
R14657 VSS.n1457 VSS.n1454 585
R14658 VSS.n1657 VSS.n1454 585
R14659 VSS.n1484 VSS.n1483 585
R14660 VSS.n1641 VSS.n1484 585
R14661 VSS.n1628 VSS.n1627 585
R14662 VSS.n1627 VSS.n1626 585
R14663 VSS.n1580 VSS.n1579 585
R14664 VSS.n1581 VSS.n1580 585
R14665 VSS.n1588 VSS.n1587 585
R14666 VSS.t92 VSS.n1588 585
R14667 VSS.n1569 VSS.n1567 585
R14668 VSS.n1590 VSS.n1569 585
R14669 VSS.n1566 VSS.n7 585
R14670 VSS.n9 VSS.n7 585
R14671 VSS.n1586 VSS.n1568 585
R14672 VSS.n1589 VSS.n1568 585
R14673 VSS.n1583 VSS.n1537 585
R14674 VSS.n1583 VSS.n1582 585
R14675 VSS.n1644 VSS.n1643 585
R14676 VSS.n1643 VSS.n1642 585
R14677 VSS.n1629 VSS.n1486 585
R14678 VSS.n1486 VSS.n1485 585
R14679 VSS.n9342 VSS.n8 585
R14680 VSS.n1451 VSS.n1450 585
R14681 VSS.n1655 VSS.n1654 585
R14682 VSS.n1656 VSS.n1655 585
R14683 VSS.n1217 VSS.n1216 585
R14684 VSS.n1219 VSS.n1217 585
R14685 VSS.n1245 VSS.n1244 585
R14686 VSS.n1246 VSS.n1245 585
R14687 VSS.n1202 VSS.n1200 585
R14688 VSS.n1250 VSS.n1202 585
R14689 VSS.n1172 VSS.n1170 585
R14690 VSS.n1281 VSS.n1172 585
R14691 VSS.n1150 VSS.n1149 585
R14692 VSS.n1282 VSS.n1149 585
R14693 VSS.n1158 VSS.n1148 585
R14694 VSS.n1313 VSS.n1148 585
R14695 VSS.n1279 VSS.n1278 585
R14696 VSS.n1280 VSS.n1279 585
R14697 VSS.n1248 VSS.n1182 585
R14698 VSS.n1249 VSS.n1248 585
R14699 VSS.n1243 VSS.n1201 585
R14700 VSS.n1247 VSS.n1201 585
R14701 VSS.n1179 VSS.n1178 585
R14702 VSS.n1283 VSS.n1179 585
R14703 VSS.n1315 VSS.n1147 585
R14704 VSS.n1315 VSS.n1314 585
R14705 VSS.n1222 VSS.n1221 585
R14706 VSS.n1221 VSS.n1220 585
R14707 VSS.n1956 VSS.n1955 585
R14708 VSS.n1955 VSS.n1954 585
R14709 VSS.n1979 VSS.n1978 585
R14710 VSS.n1980 VSS.n1979 585
R14711 VSS.n1985 VSS.n1948 585
R14712 VSS.n1948 VSS.n1947 585
R14713 VSS.n1993 VSS.n1944 585
R14714 VSS.n1944 VSS.n1943 585
R14715 VSS.n2008 VSS.n2007 585
R14716 VSS.n2007 VSS.t172 585
R14717 VSS.n2020 VSS.n2019 585
R14718 VSS.n2021 VSS.n2020 585
R14719 VSS.n1992 VSS.n1991 585
R14720 VSS.n1991 VSS.n1990 585
R14721 VSS.n1987 VSS.n1986 585
R14722 VSS.n1988 VSS.n1987 585
R14723 VSS.n1977 VSS.n1951 585
R14724 VSS.n1981 VSS.n1951 585
R14725 VSS.n1942 VSS.n1941 585
R14726 VSS.n2006 VSS.n1942 585
R14727 VSS.n1933 VSS.n1932 585
R14728 VSS.n2022 VSS.n1933 585
R14729 VSS.n1714 VSS.n1713 585
R14730 VSS.n1713 VSS.n1712 585
R14731 VSS.n2030 VSS.n2027 585
R14732 VSS.n2249 VSS.n2027 585
R14733 VSS.n2057 VSS.n2056 585
R14734 VSS.n2233 VSS.n2057 585
R14735 VSS.n2220 VSS.n2219 585
R14736 VSS.n2219 VSS.n2218 585
R14737 VSS.n2140 VSS.n2139 585
R14738 VSS.n2141 VSS.n2140 585
R14739 VSS.n2148 VSS.n2147 585
R14740 VSS.t244 VSS.n2148 585
R14741 VSS.n2129 VSS.n2127 585
R14742 VSS.n2182 VSS.n2129 585
R14743 VSS.n2180 VSS.n2179 585
R14744 VSS.n2181 VSS.n2180 585
R14745 VSS.n2146 VSS.n2128 585
R14746 VSS.n2149 VSS.n2128 585
R14747 VSS.n2143 VSS.n2110 585
R14748 VSS.n2143 VSS.n2142 585
R14749 VSS.n2236 VSS.n2235 585
R14750 VSS.n2235 VSS.n2234 585
R14751 VSS.n2221 VSS.n2059 585
R14752 VSS.n2059 VSS.n2058 585
R14753 VSS.n2157 VSS.n2156 585
R14754 VSS.n2024 VSS.n2023 585
R14755 VSS.n2247 VSS.n2246 585
R14756 VSS.n2248 VSS.n2247 585
R14757 VSS.n1790 VSS.n1789 585
R14758 VSS.n1792 VSS.n1790 585
R14759 VSS.n1818 VSS.n1817 585
R14760 VSS.n1819 VSS.n1818 585
R14761 VSS.n1775 VSS.n1773 585
R14762 VSS.n1823 VSS.n1775 585
R14763 VSS.n1745 VSS.n1743 585
R14764 VSS.n1854 VSS.n1745 585
R14765 VSS.n1723 VSS.n1722 585
R14766 VSS.n1855 VSS.n1722 585
R14767 VSS.n1731 VSS.n1721 585
R14768 VSS.n1886 VSS.n1721 585
R14769 VSS.n1852 VSS.n1851 585
R14770 VSS.n1853 VSS.n1852 585
R14771 VSS.n1821 VSS.n1755 585
R14772 VSS.n1822 VSS.n1821 585
R14773 VSS.n1816 VSS.n1774 585
R14774 VSS.n1820 VSS.n1774 585
R14775 VSS.n1752 VSS.n1751 585
R14776 VSS.n1856 VSS.n1752 585
R14777 VSS.n1888 VSS.n1720 585
R14778 VSS.n1888 VSS.n1887 585
R14779 VSS.n1795 VSS.n1794 585
R14780 VSS.n1794 VSS.n1793 585
R14781 VSS.n3503 VSS.n3492 585
R14782 VSS.n3505 VSS.n3492 585
R14783 VSS.n3491 VSS.n3490 585
R14784 VSS.n3710 VSS.n3491 585
R14785 VSS.n3730 VSS.n3729 585
R14786 VSS.n3731 VSS.n3730 585
R14787 VSS.n3458 VSS.n3457 585
R14788 VSS.n3457 VSS.n3456 585
R14789 VSS.n3765 VSS.n3764 585
R14790 VSS.n3764 VSS.t248 585
R14791 VSS.n3783 VSS.n3782 585
R14792 VSS.n3784 VSS.n3783 585
R14793 VSS.n3476 VSS.n3474 585
R14794 VSS.n3733 VSS.n3476 585
R14795 VSS.n3475 VSS.n3473 585
R14796 VSS.n3732 VSS.n3475 585
R14797 VSS.n3713 VSS.n3712 585
R14798 VSS.n3712 VSS.n3711 585
R14799 VSS.n3455 VSS.n3454 585
R14800 VSS.n3763 VSS.n3455 585
R14801 VSS.n3440 VSS.n3439 585
R14802 VSS.n3785 VSS.n3440 585
R14803 VSS.n3508 VSS.n3507 585
R14804 VSS.n3507 VSS.n3506 585
R14805 VSS.n3796 VSS.n3792 585
R14806 VSS.n3800 VSS.n3792 585
R14807 VSS.n3844 VSS.n3843 585
R14808 VSS.n3845 VSS.n3844 585
R14809 VSS.n3417 VSS.n3415 585
R14810 VSS.n3847 VSS.n3417 585
R14811 VSS.n3900 VSS.n3899 585
R14812 VSS.n3899 VSS.n3898 585
R14813 VSS.n3383 VSS.n3382 585
R14814 VSS.t15 VSS.n3383 585
R14815 VSS.n3942 VSS.n3941 585
R14816 VSS.n3943 VSS.n3942 585
R14817 VSS.n3940 VSS.n3370 585
R14818 VSS.n3944 VSS.n3370 585
R14819 VSS.n3920 VSS.n3919 585
R14820 VSS.n3919 VSS.n3918 585
R14821 VSS.n3901 VSS.n3385 585
R14822 VSS.n3385 VSS.n3384 585
R14823 VSS.n3420 VSS.n3419 585
R14824 VSS.n3419 VSS.n3418 585
R14825 VSS.n3850 VSS.n3849 585
R14826 VSS.n3849 VSS.n3848 585
R14827 VSS.n3945 VSS.n3371 585
R14828 VSS.n3787 VSS.n3786 585
R14829 VSS.n3798 VSS.n3797 585
R14830 VSS.n3799 VSS.n3798 585
R14831 VSS.n3584 VSS.n3583 585
R14832 VSS.n3586 VSS.n3584 585
R14833 VSS.n3612 VSS.n3611 585
R14834 VSS.n3613 VSS.n3612 585
R14835 VSS.n3569 VSS.n3567 585
R14836 VSS.n3617 VSS.n3569 585
R14837 VSS.n3539 VSS.n3537 585
R14838 VSS.n3648 VSS.n3539 585
R14839 VSS.n3517 VSS.n3516 585
R14840 VSS.n3649 VSS.n3516 585
R14841 VSS.n3525 VSS.n3515 585
R14842 VSS.n3680 VSS.n3515 585
R14843 VSS.n3646 VSS.n3645 585
R14844 VSS.n3647 VSS.n3646 585
R14845 VSS.n3615 VSS.n3549 585
R14846 VSS.n3616 VSS.n3615 585
R14847 VSS.n3610 VSS.n3568 585
R14848 VSS.n3614 VSS.n3568 585
R14849 VSS.n3546 VSS.n3545 585
R14850 VSS.n3650 VSS.n3546 585
R14851 VSS.n3682 VSS.n3514 585
R14852 VSS.n3682 VSS.n3681 585
R14853 VSS.n3589 VSS.n3588 585
R14854 VSS.n3588 VSS.n3587 585
R14855 VSS.n4095 VSS.n4084 585
R14856 VSS.n4097 VSS.n4084 585
R14857 VSS.n4083 VSS.n4082 585
R14858 VSS.n4302 VSS.n4083 585
R14859 VSS.n4322 VSS.n4321 585
R14860 VSS.n4323 VSS.n4322 585
R14861 VSS.n4050 VSS.n4049 585
R14862 VSS.n4049 VSS.n4048 585
R14863 VSS.n4357 VSS.n4356 585
R14864 VSS.n4356 VSS.t170 585
R14865 VSS.n4375 VSS.n4374 585
R14866 VSS.n4376 VSS.n4375 585
R14867 VSS.n4068 VSS.n4066 585
R14868 VSS.n4325 VSS.n4068 585
R14869 VSS.n4067 VSS.n4065 585
R14870 VSS.n4324 VSS.n4067 585
R14871 VSS.n4305 VSS.n4304 585
R14872 VSS.n4304 VSS.n4303 585
R14873 VSS.n4047 VSS.n4046 585
R14874 VSS.n4355 VSS.n4047 585
R14875 VSS.n4032 VSS.n4031 585
R14876 VSS.n4377 VSS.n4032 585
R14877 VSS.n4100 VSS.n4099 585
R14878 VSS.n4099 VSS.n4098 585
R14879 VSS.n4388 VSS.n4384 585
R14880 VSS.n4392 VSS.n4384 585
R14881 VSS.n4436 VSS.n4435 585
R14882 VSS.n4437 VSS.n4436 585
R14883 VSS.n4009 VSS.n4007 585
R14884 VSS.n4439 VSS.n4009 585
R14885 VSS.n4492 VSS.n4491 585
R14886 VSS.n4491 VSS.n4490 585
R14887 VSS.n3975 VSS.n3974 585
R14888 VSS.t120 VSS.n3975 585
R14889 VSS.n4534 VSS.n4533 585
R14890 VSS.n4535 VSS.n4534 585
R14891 VSS.n4532 VSS.n3962 585
R14892 VSS.n4536 VSS.n3962 585
R14893 VSS.n4512 VSS.n4511 585
R14894 VSS.n4511 VSS.n4510 585
R14895 VSS.n4493 VSS.n3977 585
R14896 VSS.n3977 VSS.n3976 585
R14897 VSS.n4012 VSS.n4011 585
R14898 VSS.n4011 VSS.n4010 585
R14899 VSS.n4442 VSS.n4441 585
R14900 VSS.n4441 VSS.n4440 585
R14901 VSS.n4537 VSS.n3963 585
R14902 VSS.n4379 VSS.n4378 585
R14903 VSS.n4390 VSS.n4389 585
R14904 VSS.n4391 VSS.n4390 585
R14905 VSS.n4176 VSS.n4175 585
R14906 VSS.n4178 VSS.n4176 585
R14907 VSS.n4204 VSS.n4203 585
R14908 VSS.n4205 VSS.n4204 585
R14909 VSS.n4161 VSS.n4159 585
R14910 VSS.n4209 VSS.n4161 585
R14911 VSS.n4131 VSS.n4129 585
R14912 VSS.n4240 VSS.n4131 585
R14913 VSS.n4109 VSS.n4108 585
R14914 VSS.n4241 VSS.n4108 585
R14915 VSS.n4117 VSS.n4107 585
R14916 VSS.n4272 VSS.n4107 585
R14917 VSS.n4238 VSS.n4237 585
R14918 VSS.n4239 VSS.n4238 585
R14919 VSS.n4207 VSS.n4141 585
R14920 VSS.n4208 VSS.n4207 585
R14921 VSS.n4202 VSS.n4160 585
R14922 VSS.n4206 VSS.n4160 585
R14923 VSS.n4138 VSS.n4137 585
R14924 VSS.n4242 VSS.n4138 585
R14925 VSS.n4274 VSS.n4106 585
R14926 VSS.n4274 VSS.n4273 585
R14927 VSS.n4181 VSS.n4180 585
R14928 VSS.n4180 VSS.n4179 585
R14929 VSS.n4687 VSS.n4676 585
R14930 VSS.n4689 VSS.n4676 585
R14931 VSS.n4675 VSS.n4674 585
R14932 VSS.n4894 VSS.n4675 585
R14933 VSS.n4914 VSS.n4913 585
R14934 VSS.n4915 VSS.n4914 585
R14935 VSS.n4642 VSS.n4641 585
R14936 VSS.n4641 VSS.n4640 585
R14937 VSS.n4949 VSS.n4948 585
R14938 VSS.n4948 VSS.t127 585
R14939 VSS.n4967 VSS.n4966 585
R14940 VSS.n4968 VSS.n4967 585
R14941 VSS.n4660 VSS.n4658 585
R14942 VSS.n4917 VSS.n4660 585
R14943 VSS.n4659 VSS.n4657 585
R14944 VSS.n4916 VSS.n4659 585
R14945 VSS.n4897 VSS.n4896 585
R14946 VSS.n4896 VSS.n4895 585
R14947 VSS.n4639 VSS.n4638 585
R14948 VSS.n4947 VSS.n4639 585
R14949 VSS.n4624 VSS.n4623 585
R14950 VSS.n4969 VSS.n4624 585
R14951 VSS.n4692 VSS.n4691 585
R14952 VSS.n4691 VSS.n4690 585
R14953 VSS.n4980 VSS.n4976 585
R14954 VSS.n4984 VSS.n4976 585
R14955 VSS.n5028 VSS.n5027 585
R14956 VSS.n5029 VSS.n5028 585
R14957 VSS.n4601 VSS.n4599 585
R14958 VSS.n5031 VSS.n4601 585
R14959 VSS.n5084 VSS.n5083 585
R14960 VSS.n5083 VSS.n5082 585
R14961 VSS.n4567 VSS.n4566 585
R14962 VSS.t272 VSS.n4567 585
R14963 VSS.n5126 VSS.n5125 585
R14964 VSS.n5127 VSS.n5126 585
R14965 VSS.n5124 VSS.n4554 585
R14966 VSS.n5128 VSS.n4554 585
R14967 VSS.n5104 VSS.n5103 585
R14968 VSS.n5103 VSS.n5102 585
R14969 VSS.n5085 VSS.n4569 585
R14970 VSS.n4569 VSS.n4568 585
R14971 VSS.n4604 VSS.n4603 585
R14972 VSS.n4603 VSS.n4602 585
R14973 VSS.n5034 VSS.n5033 585
R14974 VSS.n5033 VSS.n5032 585
R14975 VSS.n5129 VSS.n4555 585
R14976 VSS.n4971 VSS.n4970 585
R14977 VSS.n4982 VSS.n4981 585
R14978 VSS.n4983 VSS.n4982 585
R14979 VSS.n4768 VSS.n4767 585
R14980 VSS.n4770 VSS.n4768 585
R14981 VSS.n4796 VSS.n4795 585
R14982 VSS.n4797 VSS.n4796 585
R14983 VSS.n4753 VSS.n4751 585
R14984 VSS.n4801 VSS.n4753 585
R14985 VSS.n4723 VSS.n4721 585
R14986 VSS.n4832 VSS.n4723 585
R14987 VSS.n4701 VSS.n4700 585
R14988 VSS.n4833 VSS.n4700 585
R14989 VSS.n4709 VSS.n4699 585
R14990 VSS.n4864 VSS.n4699 585
R14991 VSS.n4830 VSS.n4829 585
R14992 VSS.n4831 VSS.n4830 585
R14993 VSS.n4799 VSS.n4733 585
R14994 VSS.n4800 VSS.n4799 585
R14995 VSS.n4794 VSS.n4752 585
R14996 VSS.n4798 VSS.n4752 585
R14997 VSS.n4730 VSS.n4729 585
R14998 VSS.n4834 VSS.n4730 585
R14999 VSS.n4866 VSS.n4698 585
R15000 VSS.n4866 VSS.n4865 585
R15001 VSS.n4773 VSS.n4772 585
R15002 VSS.n4772 VSS.n4771 585
R15003 VSS.n5279 VSS.n5268 585
R15004 VSS.n5281 VSS.n5268 585
R15005 VSS.n5267 VSS.n5266 585
R15006 VSS.n5486 VSS.n5267 585
R15007 VSS.n5506 VSS.n5505 585
R15008 VSS.n5507 VSS.n5506 585
R15009 VSS.n5234 VSS.n5233 585
R15010 VSS.n5233 VSS.n5232 585
R15011 VSS.n5541 VSS.n5540 585
R15012 VSS.n5540 VSS.t96 585
R15013 VSS.n5559 VSS.n5558 585
R15014 VSS.n5560 VSS.n5559 585
R15015 VSS.n5252 VSS.n5250 585
R15016 VSS.n5509 VSS.n5252 585
R15017 VSS.n5251 VSS.n5249 585
R15018 VSS.n5508 VSS.n5251 585
R15019 VSS.n5489 VSS.n5488 585
R15020 VSS.n5488 VSS.n5487 585
R15021 VSS.n5231 VSS.n5230 585
R15022 VSS.n5539 VSS.n5231 585
R15023 VSS.n5216 VSS.n5215 585
R15024 VSS.n5561 VSS.n5216 585
R15025 VSS.n5284 VSS.n5283 585
R15026 VSS.n5283 VSS.n5282 585
R15027 VSS.n5572 VSS.n5568 585
R15028 VSS.n5576 VSS.n5568 585
R15029 VSS.n5620 VSS.n5619 585
R15030 VSS.n5621 VSS.n5620 585
R15031 VSS.n5193 VSS.n5191 585
R15032 VSS.n5623 VSS.n5193 585
R15033 VSS.n5676 VSS.n5675 585
R15034 VSS.n5675 VSS.n5674 585
R15035 VSS.n5159 VSS.n5158 585
R15036 VSS.t106 VSS.n5159 585
R15037 VSS.n5718 VSS.n5717 585
R15038 VSS.n5719 VSS.n5718 585
R15039 VSS.n5716 VSS.n5146 585
R15040 VSS.n5720 VSS.n5146 585
R15041 VSS.n5696 VSS.n5695 585
R15042 VSS.n5695 VSS.n5694 585
R15043 VSS.n5677 VSS.n5161 585
R15044 VSS.n5161 VSS.n5160 585
R15045 VSS.n5196 VSS.n5195 585
R15046 VSS.n5195 VSS.n5194 585
R15047 VSS.n5626 VSS.n5625 585
R15048 VSS.n5625 VSS.n5624 585
R15049 VSS.n5721 VSS.n5147 585
R15050 VSS.n5563 VSS.n5562 585
R15051 VSS.n5574 VSS.n5573 585
R15052 VSS.n5575 VSS.n5574 585
R15053 VSS.n5360 VSS.n5359 585
R15054 VSS.n5362 VSS.n5360 585
R15055 VSS.n5388 VSS.n5387 585
R15056 VSS.n5389 VSS.n5388 585
R15057 VSS.n5345 VSS.n5343 585
R15058 VSS.n5393 VSS.n5345 585
R15059 VSS.n5315 VSS.n5313 585
R15060 VSS.n5424 VSS.n5315 585
R15061 VSS.n5293 VSS.n5292 585
R15062 VSS.n5425 VSS.n5292 585
R15063 VSS.n5301 VSS.n5291 585
R15064 VSS.n5456 VSS.n5291 585
R15065 VSS.n5422 VSS.n5421 585
R15066 VSS.n5423 VSS.n5422 585
R15067 VSS.n5391 VSS.n5325 585
R15068 VSS.n5392 VSS.n5391 585
R15069 VSS.n5386 VSS.n5344 585
R15070 VSS.n5390 VSS.n5344 585
R15071 VSS.n5322 VSS.n5321 585
R15072 VSS.n5426 VSS.n5322 585
R15073 VSS.n5458 VSS.n5290 585
R15074 VSS.n5458 VSS.n5457 585
R15075 VSS.n5365 VSS.n5364 585
R15076 VSS.n5364 VSS.n5363 585
R15077 VSS.n5871 VSS.n5860 585
R15078 VSS.n5873 VSS.n5860 585
R15079 VSS.n5859 VSS.n5858 585
R15080 VSS.n6078 VSS.n5859 585
R15081 VSS.n6098 VSS.n6097 585
R15082 VSS.n6099 VSS.n6098 585
R15083 VSS.n5826 VSS.n5825 585
R15084 VSS.n5825 VSS.n5824 585
R15085 VSS.n6133 VSS.n6132 585
R15086 VSS.n6132 VSS.t188 585
R15087 VSS.n6151 VSS.n6150 585
R15088 VSS.n6152 VSS.n6151 585
R15089 VSS.n5844 VSS.n5842 585
R15090 VSS.n6101 VSS.n5844 585
R15091 VSS.n5843 VSS.n5841 585
R15092 VSS.n6100 VSS.n5843 585
R15093 VSS.n6081 VSS.n6080 585
R15094 VSS.n6080 VSS.n6079 585
R15095 VSS.n5823 VSS.n5822 585
R15096 VSS.n6131 VSS.n5823 585
R15097 VSS.n5808 VSS.n5807 585
R15098 VSS.n6153 VSS.n5808 585
R15099 VSS.n5876 VSS.n5875 585
R15100 VSS.n5875 VSS.n5874 585
R15101 VSS.n6164 VSS.n6160 585
R15102 VSS.n6168 VSS.n6160 585
R15103 VSS.n6212 VSS.n6211 585
R15104 VSS.n6213 VSS.n6212 585
R15105 VSS.n5785 VSS.n5783 585
R15106 VSS.n6215 VSS.n5785 585
R15107 VSS.n6268 VSS.n6267 585
R15108 VSS.n6267 VSS.n6266 585
R15109 VSS.n5751 VSS.n5750 585
R15110 VSS.t281 VSS.n5751 585
R15111 VSS.n6310 VSS.n6309 585
R15112 VSS.n6311 VSS.n6310 585
R15113 VSS.n6308 VSS.n5738 585
R15114 VSS.n6312 VSS.n5738 585
R15115 VSS.n6288 VSS.n6287 585
R15116 VSS.n6287 VSS.n6286 585
R15117 VSS.n6269 VSS.n5753 585
R15118 VSS.n5753 VSS.n5752 585
R15119 VSS.n5788 VSS.n5787 585
R15120 VSS.n5787 VSS.n5786 585
R15121 VSS.n6218 VSS.n6217 585
R15122 VSS.n6217 VSS.n6216 585
R15123 VSS.n6313 VSS.n5739 585
R15124 VSS.n6155 VSS.n6154 585
R15125 VSS.n6166 VSS.n6165 585
R15126 VSS.n6167 VSS.n6166 585
R15127 VSS.n5952 VSS.n5951 585
R15128 VSS.n5954 VSS.n5952 585
R15129 VSS.n5980 VSS.n5979 585
R15130 VSS.n5981 VSS.n5980 585
R15131 VSS.n5937 VSS.n5935 585
R15132 VSS.n5985 VSS.n5937 585
R15133 VSS.n5907 VSS.n5905 585
R15134 VSS.n6016 VSS.n5907 585
R15135 VSS.n5885 VSS.n5884 585
R15136 VSS.n6017 VSS.n5884 585
R15137 VSS.n5893 VSS.n5883 585
R15138 VSS.n6048 VSS.n5883 585
R15139 VSS.n6014 VSS.n6013 585
R15140 VSS.n6015 VSS.n6014 585
R15141 VSS.n5983 VSS.n5917 585
R15142 VSS.n5984 VSS.n5983 585
R15143 VSS.n5978 VSS.n5936 585
R15144 VSS.n5982 VSS.n5936 585
R15145 VSS.n5914 VSS.n5913 585
R15146 VSS.n6018 VSS.n5914 585
R15147 VSS.n6050 VSS.n5882 585
R15148 VSS.n6050 VSS.n6049 585
R15149 VSS.n5957 VSS.n5956 585
R15150 VSS.n5956 VSS.n5955 585
R15151 VSS.n6463 VSS.n6452 585
R15152 VSS.n6465 VSS.n6452 585
R15153 VSS.n6451 VSS.n6450 585
R15154 VSS.n6670 VSS.n6451 585
R15155 VSS.n6690 VSS.n6689 585
R15156 VSS.n6691 VSS.n6690 585
R15157 VSS.n6418 VSS.n6417 585
R15158 VSS.n6417 VSS.n6416 585
R15159 VSS.n6725 VSS.n6724 585
R15160 VSS.n6724 VSS.t236 585
R15161 VSS.n6743 VSS.n6742 585
R15162 VSS.n6744 VSS.n6743 585
R15163 VSS.n6436 VSS.n6434 585
R15164 VSS.n6693 VSS.n6436 585
R15165 VSS.n6435 VSS.n6433 585
R15166 VSS.n6692 VSS.n6435 585
R15167 VSS.n6673 VSS.n6672 585
R15168 VSS.n6672 VSS.n6671 585
R15169 VSS.n6415 VSS.n6414 585
R15170 VSS.n6723 VSS.n6415 585
R15171 VSS.n6400 VSS.n6399 585
R15172 VSS.n6745 VSS.n6400 585
R15173 VSS.n6468 VSS.n6467 585
R15174 VSS.n6467 VSS.n6466 585
R15175 VSS.n6756 VSS.n6752 585
R15176 VSS.n6760 VSS.n6752 585
R15177 VSS.n6804 VSS.n6803 585
R15178 VSS.n6805 VSS.n6804 585
R15179 VSS.n6377 VSS.n6375 585
R15180 VSS.n6807 VSS.n6377 585
R15181 VSS.n6860 VSS.n6859 585
R15182 VSS.n6859 VSS.n6858 585
R15183 VSS.n6343 VSS.n6342 585
R15184 VSS.t205 VSS.n6343 585
R15185 VSS.n6902 VSS.n6901 585
R15186 VSS.n6903 VSS.n6902 585
R15187 VSS.n6900 VSS.n6330 585
R15188 VSS.n6904 VSS.n6330 585
R15189 VSS.n6880 VSS.n6879 585
R15190 VSS.n6879 VSS.n6878 585
R15191 VSS.n6861 VSS.n6345 585
R15192 VSS.n6345 VSS.n6344 585
R15193 VSS.n6380 VSS.n6379 585
R15194 VSS.n6379 VSS.n6378 585
R15195 VSS.n6810 VSS.n6809 585
R15196 VSS.n6809 VSS.n6808 585
R15197 VSS.n6905 VSS.n6331 585
R15198 VSS.n6747 VSS.n6746 585
R15199 VSS.n6758 VSS.n6757 585
R15200 VSS.n6759 VSS.n6758 585
R15201 VSS.n6544 VSS.n6543 585
R15202 VSS.n6546 VSS.n6544 585
R15203 VSS.n6572 VSS.n6571 585
R15204 VSS.n6573 VSS.n6572 585
R15205 VSS.n6529 VSS.n6527 585
R15206 VSS.n6577 VSS.n6529 585
R15207 VSS.n6499 VSS.n6497 585
R15208 VSS.n6608 VSS.n6499 585
R15209 VSS.n6477 VSS.n6476 585
R15210 VSS.n6609 VSS.n6476 585
R15211 VSS.n6485 VSS.n6475 585
R15212 VSS.n6640 VSS.n6475 585
R15213 VSS.n6606 VSS.n6605 585
R15214 VSS.n6607 VSS.n6606 585
R15215 VSS.n6575 VSS.n6509 585
R15216 VSS.n6576 VSS.n6575 585
R15217 VSS.n6570 VSS.n6528 585
R15218 VSS.n6574 VSS.n6528 585
R15219 VSS.n6506 VSS.n6505 585
R15220 VSS.n6610 VSS.n6506 585
R15221 VSS.n6642 VSS.n6474 585
R15222 VSS.n6642 VSS.n6641 585
R15223 VSS.n6549 VSS.n6548 585
R15224 VSS.n6548 VSS.n6547 585
R15225 VSS.n2554 VSS.n2553 585
R15226 VSS.n2553 VSS.n2552 585
R15227 VSS.n2577 VSS.n2576 585
R15228 VSS.n2578 VSS.n2577 585
R15229 VSS.n2583 VSS.n2546 585
R15230 VSS.n2546 VSS.n2545 585
R15231 VSS.n2591 VSS.n2542 585
R15232 VSS.n2542 VSS.n2541 585
R15233 VSS.n2606 VSS.n2605 585
R15234 VSS.n2605 VSS.t151 585
R15235 VSS.n2618 VSS.n2617 585
R15236 VSS.n2619 VSS.n2618 585
R15237 VSS.n2590 VSS.n2589 585
R15238 VSS.n2589 VSS.n2588 585
R15239 VSS.n2585 VSS.n2584 585
R15240 VSS.n2586 VSS.n2585 585
R15241 VSS.n2575 VSS.n2549 585
R15242 VSS.n2579 VSS.n2549 585
R15243 VSS.n2540 VSS.n2539 585
R15244 VSS.n2604 VSS.n2540 585
R15245 VSS.n2531 VSS.n2530 585
R15246 VSS.n2620 VSS.n2531 585
R15247 VSS.n2312 VSS.n2311 585
R15248 VSS.n2311 VSS.n2310 585
R15249 VSS.n2628 VSS.n2625 585
R15250 VSS.n6993 VSS.n2625 585
R15251 VSS.n2655 VSS.n2654 585
R15252 VSS.n6977 VSS.n2655 585
R15253 VSS.n6964 VSS.n6963 585
R15254 VSS.n6963 VSS.n6962 585
R15255 VSS.n2738 VSS.n2737 585
R15256 VSS.n2739 VSS.n2738 585
R15257 VSS.n2746 VSS.n2745 585
R15258 VSS.t55 VSS.n2746 585
R15259 VSS.n2727 VSS.n2725 585
R15260 VSS.n6926 VSS.n2727 585
R15261 VSS.n6924 VSS.n6923 585
R15262 VSS.n6925 VSS.n6924 585
R15263 VSS.n2744 VSS.n2726 585
R15264 VSS.n2747 VSS.n2726 585
R15265 VSS.n2741 VSS.n2708 585
R15266 VSS.n2741 VSS.n2740 585
R15267 VSS.n6980 VSS.n6979 585
R15268 VSS.n6979 VSS.n6978 585
R15269 VSS.n6965 VSS.n2657 585
R15270 VSS.n2657 VSS.n2656 585
R15271 VSS.n2755 VSS.n2754 585
R15272 VSS.n2622 VSS.n2621 585
R15273 VSS.n6991 VSS.n6990 585
R15274 VSS.n6992 VSS.n6991 585
R15275 VSS.n2388 VSS.n2387 585
R15276 VSS.n2390 VSS.n2388 585
R15277 VSS.n2416 VSS.n2415 585
R15278 VSS.n2417 VSS.n2416 585
R15279 VSS.n2373 VSS.n2371 585
R15280 VSS.n2421 VSS.n2373 585
R15281 VSS.n2343 VSS.n2341 585
R15282 VSS.n2452 VSS.n2343 585
R15283 VSS.n2321 VSS.n2320 585
R15284 VSS.n2453 VSS.n2320 585
R15285 VSS.n2329 VSS.n2319 585
R15286 VSS.n2484 VSS.n2319 585
R15287 VSS.n2450 VSS.n2449 585
R15288 VSS.n2451 VSS.n2450 585
R15289 VSS.n2419 VSS.n2353 585
R15290 VSS.n2420 VSS.n2419 585
R15291 VSS.n2414 VSS.n2372 585
R15292 VSS.n2418 VSS.n2372 585
R15293 VSS.n2350 VSS.n2349 585
R15294 VSS.n2454 VSS.n2350 585
R15295 VSS.n2486 VSS.n2318 585
R15296 VSS.n2486 VSS.n2485 585
R15297 VSS.n2393 VSS.n2392 585
R15298 VSS.n2392 VSS.n2391 585
R15299 VSS.n2910 VSS.n2899 585
R15300 VSS.n2912 VSS.n2899 585
R15301 VSS.n2898 VSS.n2897 585
R15302 VSS.n3118 VSS.n2898 585
R15303 VSS.n3138 VSS.n3137 585
R15304 VSS.n3139 VSS.n3138 585
R15305 VSS.n2865 VSS.n2864 585
R15306 VSS.n2864 VSS.n2863 585
R15307 VSS.n3173 VSS.n3172 585
R15308 VSS.n3172 VSS.t24 585
R15309 VSS.n3191 VSS.n3190 585
R15310 VSS.n3192 VSS.n3191 585
R15311 VSS.n2883 VSS.n2881 585
R15312 VSS.n3141 VSS.n2883 585
R15313 VSS.n2882 VSS.n2880 585
R15314 VSS.n3140 VSS.n2882 585
R15315 VSS.n3121 VSS.n3120 585
R15316 VSS.n3120 VSS.n3119 585
R15317 VSS.n2862 VSS.n2861 585
R15318 VSS.n3171 VSS.n2862 585
R15319 VSS.n2847 VSS.n2846 585
R15320 VSS.n3193 VSS.n2847 585
R15321 VSS.n2915 VSS.n2914 585
R15322 VSS.n2914 VSS.n2913 585
R15323 VSS.n3204 VSS.n3200 585
R15324 VSS.n3208 VSS.n3200 585
R15325 VSS.n3252 VSS.n3251 585
R15326 VSS.n3253 VSS.n3252 585
R15327 VSS.n2824 VSS.n2822 585
R15328 VSS.n3255 VSS.n2824 585
R15329 VSS.n3308 VSS.n3307 585
R15330 VSS.n3307 VSS.n3306 585
R15331 VSS.n2790 VSS.n2789 585
R15332 VSS.t4 VSS.n2790 585
R15333 VSS.n3350 VSS.n3349 585
R15334 VSS.n3351 VSS.n3350 585
R15335 VSS.n3348 VSS.n2777 585
R15336 VSS.n3352 VSS.n2777 585
R15337 VSS.n3328 VSS.n3327 585
R15338 VSS.n3327 VSS.n3326 585
R15339 VSS.n3309 VSS.n2792 585
R15340 VSS.n2792 VSS.n2791 585
R15341 VSS.n2827 VSS.n2826 585
R15342 VSS.n2826 VSS.n2825 585
R15343 VSS.n3258 VSS.n3257 585
R15344 VSS.n3257 VSS.n3256 585
R15345 VSS.n3353 VSS.n2778 585
R15346 VSS.n3195 VSS.n3194 585
R15347 VSS.n3206 VSS.n3205 585
R15348 VSS.n3207 VSS.n3206 585
R15349 VSS.n2985 VSS.n2974 585
R15350 VSS.n2987 VSS.n2974 585
R15351 VSS.n2973 VSS.n2972 585
R15352 VSS.n3013 VSS.n2973 585
R15353 VSS.n3033 VSS.n3032 585
R15354 VSS.n3034 VSS.n3033 585
R15355 VSS.n2940 VSS.n2939 585
R15356 VSS.n2939 VSS.n2938 585
R15357 VSS.n3069 VSS.n3068 585
R15358 VSS.n3068 VSS.n3067 585
R15359 VSS.n3087 VSS.n3086 585
R15360 VSS.n3088 VSS.n3087 585
R15361 VSS.n2960 VSS.n2958 585
R15362 VSS.n3036 VSS.n2960 585
R15363 VSS.n2959 VSS.n2957 585
R15364 VSS.n3035 VSS.n2959 585
R15365 VSS.n3016 VSS.n3015 585
R15366 VSS.n3015 VSS.n3014 585
R15367 VSS.n2937 VSS.n2936 585
R15368 VSS.n3066 VSS.n2937 585
R15369 VSS.n2922 VSS.n2921 585
R15370 VSS.n3089 VSS.n2922 585
R15371 VSS.n2990 VSS.n2989 585
R15372 VSS.n2989 VSS.n2988 585
R15373 VSS.n186 VSS.n166 585
R15374 VSS.n184 VSS.n166 585
R15375 VSS.n165 VSS.n164 585
R15376 VSS.n9078 VSS.n165 585
R15377 VSS.n9098 VSS.n9097 585
R15378 VSS.n9099 VSS.n9098 585
R15379 VSS.n132 VSS.n131 585
R15380 VSS.n131 VSS.n130 585
R15381 VSS.n9133 VSS.n9132 585
R15382 VSS.n9132 VSS.t218 585
R15383 VSS.n9151 VSS.n9150 585
R15384 VSS.n9152 VSS.n9151 585
R15385 VSS.n150 VSS.n148 585
R15386 VSS.n9101 VSS.n150 585
R15387 VSS.n149 VSS.n147 585
R15388 VSS.n9100 VSS.n149 585
R15389 VSS.n9081 VSS.n9080 585
R15390 VSS.n9080 VSS.n9079 585
R15391 VSS.n129 VSS.n128 585
R15392 VSS.n9131 VSS.n129 585
R15393 VSS.n114 VSS.n113 585
R15394 VSS.n9153 VSS.n114 585
R15395 VSS.n188 VSS.n187 585
R15396 VSS.n188 VSS.n185 585
R15397 VSS.n9164 VSS.n9160 585
R15398 VSS.n9168 VSS.n9160 585
R15399 VSS.n9212 VSS.n9211 585
R15400 VSS.n9213 VSS.n9212 585
R15401 VSS.n91 VSS.n89 585
R15402 VSS.n9215 VSS.n91 585
R15403 VSS.n9268 VSS.n9267 585
R15404 VSS.n9267 VSS.n9266 585
R15405 VSS.n57 VSS.n56 585
R15406 VSS.t290 VSS.n57 585
R15407 VSS.n9310 VSS.n9309 585
R15408 VSS.n9311 VSS.n9310 585
R15409 VSS.n9308 VSS.n44 585
R15410 VSS.n9312 VSS.n44 585
R15411 VSS.n9288 VSS.n9287 585
R15412 VSS.n9287 VSS.n9286 585
R15413 VSS.n9269 VSS.n59 585
R15414 VSS.n59 VSS.n58 585
R15415 VSS.n94 VSS.n93 585
R15416 VSS.n93 VSS.n92 585
R15417 VSS.n9218 VSS.n9217 585
R15418 VSS.n9217 VSS.n9216 585
R15419 VSS.n9313 VSS.n45 585
R15420 VSS.n9155 VSS.n9154 585
R15421 VSS.n9166 VSS.n9165 585
R15422 VSS.n9167 VSS.n9166 585
R15423 VSS.n342 VSS.n341 585
R15424 VSS.n343 VSS.n342 585
R15425 VSS.n347 VSS.n346 585
R15426 VSS.n346 VSS.n345 585
R15427 VSS.n323 VSS.n322 585
R15428 VSS.n358 VSS.n323 585
R15429 VSS.n319 VSS.n318 585
R15430 VSS.n367 VSS.n319 585
R15431 VSS.n382 VSS.n381 585
R15432 VSS.n383 VSS.n382 585
R15433 VSS.n387 VSS.n386 585
R15434 VSS.n386 VSS.n385 585
R15435 VSS.n365 VSS.n364 585
R15436 VSS.n366 VSS.n365 585
R15437 VSS.n361 VSS.n360 585
R15438 VSS.n360 VSS.n359 585
R15439 VSS.n348 VSS.n325 585
R15440 VSS.n325 VSS.n324 585
R15441 VSS.n378 VSS.n315 585
R15442 VSS.n315 VSS.n314 585
R15443 VSS.n182 VSS.n181 585
R15444 VSS.n183 VSS.n182 585
R15445 VSS.n274 VSS.n273 585
R15446 VSS.n273 VSS.n272 585
R15447 VSS.n8701 VSS.n8700 585
R15448 VSS.n8700 VSS.n8699 585
R15449 VSS.n8724 VSS.n8723 585
R15450 VSS.n8725 VSS.n8724 585
R15451 VSS.n8730 VSS.n8693 585
R15452 VSS.n8693 VSS.n8692 585
R15453 VSS.n8738 VSS.n8689 585
R15454 VSS.n8689 VSS.n8688 585
R15455 VSS.n8753 VSS.n8752 585
R15456 VSS.n8752 VSS.t262 585
R15457 VSS.n8765 VSS.n8764 585
R15458 VSS.n8766 VSS.n8765 585
R15459 VSS.n8737 VSS.n8736 585
R15460 VSS.n8736 VSS.n8735 585
R15461 VSS.n8732 VSS.n8731 585
R15462 VSS.n8733 VSS.n8732 585
R15463 VSS.n8722 VSS.n8696 585
R15464 VSS.n8726 VSS.n8696 585
R15465 VSS.n8687 VSS.n8686 585
R15466 VSS.n8751 VSS.n8687 585
R15467 VSS.n8678 VSS.n8677 585
R15468 VSS.n8767 VSS.n8678 585
R15469 VSS.n195 VSS.n194 585
R15470 VSS.n194 VSS.n193 585
R15471 VSS.n8775 VSS.n8772 585
R15472 VSS.n8994 VSS.n8772 585
R15473 VSS.n8829 VSS.n8825 585
R15474 VSS.n8833 VSS.n8825 585
R15475 VSS.n8844 VSS.n8843 585
R15476 VSS.n8845 VSS.n8844 585
R15477 VSS.n8956 VSS.n8955 585
R15478 VSS.n8957 VSS.n8956 585
R15479 VSS.n8905 VSS.n8903 585
R15480 VSS.t142 VSS.n8903 585
R15481 VSS.n8919 VSS.n8918 585
R15482 VSS.n8920 VSS.n8919 585
R15483 VSS.n8917 VSS.n8900 585
R15484 VSS.n8921 VSS.n8900 585
R15485 VSS.n8915 VSS.n8883 585
R15486 VSS.n8915 VSS.n8914 585
R15487 VSS.n8954 VSS.n8848 585
R15488 VSS.n8848 VSS.n8847 585
R15489 VSS.n8831 VSS.n8830 585
R15490 VSS.n8832 VSS.n8831 585
R15491 VSS.n8836 VSS.n8807 585
R15492 VSS.n8836 VSS.n8824 585
R15493 VSS.n8922 VSS.n8901 585
R15494 VSS.n8769 VSS.n8768 585
R15495 VSS.n8992 VSS.n8991 585
R15496 VSS.n8993 VSS.n8992 585
R15497 VSS.n548 VSS.n547 585
R15498 VSS.n547 VSS.n546 585
R15499 VSS.n569 VSS.n568 585
R15500 VSS.n570 VSS.n569 585
R15501 VSS.n575 VSS.n535 585
R15502 VSS.n535 VSS.n534 585
R15503 VSS.n583 VSS.n531 585
R15504 VSS.n531 VSS.n530 585
R15505 VSS.n598 VSS.n597 585
R15506 VSS.n597 VSS.t27 585
R15507 VSS.n610 VSS.n609 585
R15508 VSS.n611 VSS.n610 585
R15509 VSS.n582 VSS.n581 585
R15510 VSS.n581 VSS.n580 585
R15511 VSS.n577 VSS.n576 585
R15512 VSS.n578 VSS.n577 585
R15513 VSS.n567 VSS.n538 585
R15514 VSS.n571 VSS.n538 585
R15515 VSS.n529 VSS.n528 585
R15516 VSS.n596 VSS.n529 585
R15517 VSS.n520 VSS.n519 585
R15518 VSS.n612 VSS.n520 585
R15519 VSS.n542 VSS.n541 585
R15520 VSS.n545 VSS.n542 585
R15521 VSS.n746 VSS.n745 585
R15522 VSS.n745 VSS.n744 585
R15523 VSS.n784 VSS.n649 585
R15524 VSS.n649 VSS.n648 585
R15525 VSS.n783 VSS.n782 585
R15526 VSS.n782 VSS.n781 585
R15527 VSS.n799 VSS.n798 585
R15528 VSS.n798 VSS.n797 585
R15529 VSS.n614 VSS.n613 585
R15530 VSS.n620 VSS.n617 585
R15531 VSS.n812 VSS.n617 585
R15532 VSS.n810 VSS.n809 585
R15533 VSS.n811 VSS.n810 585
R15534 VSS.n647 VSS.n646 585
R15535 VSS.n796 VSS.n647 585
R15536 VSS.n741 VSS.n700 585
R15537 VSS.n741 VSS.n729 585
R15538 VSS.n740 VSS.n738 585
R15539 VSS.n740 VSS.n739 585
R15540 VSS.n728 VSS.n727 585
R15541 VSS.t102 VSS.n728 585
R15542 VSS.n9330 VSS.n29 585
R15543 VSS.n9334 VSS.n29 585
R15544 VSS.n9332 VSS.n9331 585
R15545 VSS.n9333 VSS.n9332 585
R15546 VSS.n26 VSS.n25 585
R15547 VSS.n891 VSS.n890 585
R15548 VSS.n890 VSS.n889 585
R15549 VSS.n912 VSS.n911 585
R15550 VSS.n913 VSS.n912 585
R15551 VSS.n918 VSS.n883 585
R15552 VSS.n883 VSS.n882 585
R15553 VSS.n926 VSS.n878 585
R15554 VSS.n878 VSS.n877 585
R15555 VSS.n942 VSS.n941 585
R15556 VSS.n941 VSS.n940 585
R15557 VSS.n954 VSS.n953 585
R15558 VSS.n955 VSS.n954 585
R15559 VSS.n925 VSS.n924 585
R15560 VSS.n924 VSS.n923 585
R15561 VSS.n920 VSS.n919 585
R15562 VSS.n921 VSS.n920 585
R15563 VSS.n910 VSS.n886 585
R15564 VSS.n914 VSS.n886 585
R15565 VSS.n876 VSS.n875 585
R15566 VSS.n939 VSS.n876 585
R15567 VSS.n867 VSS.n866 585
R15568 VSS.n956 VSS.n867 585
R15569 VSS.n440 VSS.n439 585
R15570 VSS.n439 VSS.n438 585
R15571 VSS.n1072 VSS.n1071 585
R15572 VSS.n1071 VSS.n1070 585
R15573 VSS.n1093 VSS.n1092 585
R15574 VSS.n1094 VSS.n1093 585
R15575 VSS.n1099 VSS.n1064 585
R15576 VSS.n1064 VSS.n1063 585
R15577 VSS.n1107 VSS.n1059 585
R15578 VSS.n1059 VSS.n1058 585
R15579 VSS.n1123 VSS.n1122 585
R15580 VSS.n1122 VSS.n1121 585
R15581 VSS.n1135 VSS.n1134 585
R15582 VSS.n1136 VSS.n1135 585
R15583 VSS.n1106 VSS.n1105 585
R15584 VSS.n1105 VSS.n1104 585
R15585 VSS.n1101 VSS.n1100 585
R15586 VSS.n1102 VSS.n1101 585
R15587 VSS.n1091 VSS.n1067 585
R15588 VSS.n1095 VSS.n1067 585
R15589 VSS.n1057 VSS.n1056 585
R15590 VSS.n1120 VSS.n1057 585
R15591 VSS.n1048 VSS.n1047 585
R15592 VSS.n1137 VSS.n1048 585
R15593 VSS.n1007 VSS.n1006 585
R15594 VSS.n1006 VSS.n1005 585
R15595 VSS.n7974 VSS.n7973 585
R15596 VSS.n7976 VSS.n7974 585
R15597 VSS.n8002 VSS.n8001 585
R15598 VSS.n8003 VSS.n8002 585
R15599 VSS.n7959 VSS.n7957 585
R15600 VSS.n8007 VSS.n7959 585
R15601 VSS.n7929 VSS.n7927 585
R15602 VSS.n8038 VSS.n7929 585
R15603 VSS.n7907 VSS.n7906 585
R15604 VSS.n8039 VSS.n7906 585
R15605 VSS.n7915 VSS.n7905 585
R15606 VSS.n8070 VSS.n7905 585
R15607 VSS.n8036 VSS.n8035 585
R15608 VSS.n8037 VSS.n8036 585
R15609 VSS.n8005 VSS.n7939 585
R15610 VSS.n8006 VSS.n8005 585
R15611 VSS.n8000 VSS.n7958 585
R15612 VSS.n8004 VSS.n7958 585
R15613 VSS.n7936 VSS.n7935 585
R15614 VSS.n8040 VSS.n7936 585
R15615 VSS.n8072 VSS.n7904 585
R15616 VSS.n8072 VSS.n8071 585
R15617 VSS.n7979 VSS.n7978 585
R15618 VSS.n7978 VSS.n7977 585
R15619 VSS.n7122 VSS.n7121 585
R15620 VSS.n7121 VSS.n7120 585
R15621 VSS.n7145 VSS.n7144 585
R15622 VSS.n7146 VSS.n7145 585
R15623 VSS.n7151 VSS.n7114 585
R15624 VSS.n7114 VSS.n7113 585
R15625 VSS.n7159 VSS.n7110 585
R15626 VSS.n7110 VSS.n7109 585
R15627 VSS.n7174 VSS.n7173 585
R15628 VSS.n7173 VSS.t285 585
R15629 VSS.n7186 VSS.n7185 585
R15630 VSS.n7187 VSS.n7186 585
R15631 VSS.n7158 VSS.n7157 585
R15632 VSS.n7157 VSS.n7156 585
R15633 VSS.n7153 VSS.n7152 585
R15634 VSS.n7154 VSS.n7153 585
R15635 VSS.n7143 VSS.n7117 585
R15636 VSS.n7147 VSS.n7117 585
R15637 VSS.n7108 VSS.n7107 585
R15638 VSS.n7172 VSS.n7108 585
R15639 VSS.n7099 VSS.n7098 585
R15640 VSS.n7188 VSS.n7099 585
R15641 VSS.n7059 VSS.n7058 585
R15642 VSS.n7058 VSS.n7057 585
R15643 VSS.n7196 VSS.n7193 585
R15644 VSS.n8421 VSS.n7193 585
R15645 VSS.n7223 VSS.n7222 585
R15646 VSS.n8405 VSS.n7223 585
R15647 VSS.n8392 VSS.n8391 585
R15648 VSS.n8391 VSS.n8390 585
R15649 VSS.n7306 VSS.n7305 585
R15650 VSS.n7307 VSS.n7306 585
R15651 VSS.n7314 VSS.n7313 585
R15652 VSS.t301 VSS.n7314 585
R15653 VSS.n7295 VSS.n7293 585
R15654 VSS.n8354 VSS.n7295 585
R15655 VSS.n8352 VSS.n8351 585
R15656 VSS.n8353 VSS.n8352 585
R15657 VSS.n7312 VSS.n7294 585
R15658 VSS.n7315 VSS.n7294 585
R15659 VSS.n7309 VSS.n7276 585
R15660 VSS.n7309 VSS.n7308 585
R15661 VSS.n8408 VSS.n8407 585
R15662 VSS.n8407 VSS.n8406 585
R15663 VSS.n8393 VSS.n7225 585
R15664 VSS.n7225 VSS.n7224 585
R15665 VSS.n7323 VSS.n7322 585
R15666 VSS.n7190 VSS.n7189 585
R15667 VSS.n8419 VSS.n8418 585
R15668 VSS.n8420 VSS.n8419 585
R15669 VSS.n8422 VSS.n8421 403.461
R15670 VSS.n8404 VSS.n7224 403.461
R15671 VSS.n7308 VSS.n7296 403.461
R15672 VSS.n8355 VSS.n7315 403.461
R15673 VSS.n8353 VSS.n7316 403.461
R15674 VSS.n7148 VSS.n7147 396.599
R15675 VSS.n7155 VSS.n7154 396.599
R15676 VSS.n7156 VSS.n7155 396.599
R15677 VSS.n7172 VSS.n7171 396.599
R15678 VSS.n7187 VSS.n7100 396.599
R15679 VSS.n8389 VSS.n8388 395.849
R15680 VSS.n8388 VSS.n7242 395.849
R15681 VSS.n7599 VSS.n7598 338.954
R15682 VSS.n7646 VSS.n7644 338.954
R15683 VSS.n7715 VSS.n7360 338.954
R15684 VSS.n7716 VSS.n7347 338.954
R15685 VSS.n7743 VSS.n7741 338.954
R15686 VSS.n8191 VSS.n8190 338.954
R15687 VSS.n8238 VSS.n8236 338.954
R15688 VSS.n8307 VSS.n7774 338.954
R15689 VSS.n8308 VSS.n7761 338.954
R15690 VSS.n8335 VSS.n8333 338.954
R15691 VSS.n1658 VSS.n1657 338.954
R15692 VSS.n1640 VSS.n1485 338.954
R15693 VSS.n1582 VSS.n1570 338.954
R15694 VSS.n1591 VSS.n1589 338.954
R15695 VSS.n9343 VSS.n9 338.954
R15696 VSS.n2250 VSS.n2249 338.954
R15697 VSS.n2232 VSS.n2058 338.954
R15698 VSS.n2142 VSS.n2130 338.954
R15699 VSS.n2183 VSS.n2149 338.954
R15700 VSS.n2181 VSS.n2150 338.954
R15701 VSS.n3801 VSS.n3800 338.954
R15702 VSS.n3848 VSS.n3846 338.954
R15703 VSS.n3917 VSS.n3384 338.954
R15704 VSS.n3918 VSS.n3372 338.954
R15705 VSS.n3946 VSS.n3944 338.954
R15706 VSS.n4393 VSS.n4392 338.954
R15707 VSS.n4440 VSS.n4438 338.954
R15708 VSS.n4509 VSS.n3976 338.954
R15709 VSS.n4510 VSS.n3964 338.954
R15710 VSS.n4538 VSS.n4536 338.954
R15711 VSS.n4985 VSS.n4984 338.954
R15712 VSS.n5032 VSS.n5030 338.954
R15713 VSS.n5101 VSS.n4568 338.954
R15714 VSS.n5102 VSS.n4556 338.954
R15715 VSS.n5130 VSS.n5128 338.954
R15716 VSS.n5577 VSS.n5576 338.954
R15717 VSS.n5624 VSS.n5622 338.954
R15718 VSS.n5693 VSS.n5160 338.954
R15719 VSS.n5694 VSS.n5148 338.954
R15720 VSS.n5722 VSS.n5720 338.954
R15721 VSS.n6169 VSS.n6168 338.954
R15722 VSS.n6216 VSS.n6214 338.954
R15723 VSS.n6285 VSS.n5752 338.954
R15724 VSS.n6286 VSS.n5740 338.954
R15725 VSS.n6314 VSS.n6312 338.954
R15726 VSS.n6761 VSS.n6760 338.954
R15727 VSS.n6808 VSS.n6806 338.954
R15728 VSS.n6877 VSS.n6344 338.954
R15729 VSS.n6878 VSS.n6332 338.954
R15730 VSS.n6906 VSS.n6904 338.954
R15731 VSS.n6994 VSS.n6993 338.954
R15732 VSS.n6976 VSS.n2656 338.954
R15733 VSS.n2740 VSS.n2728 338.954
R15734 VSS.n6927 VSS.n2747 338.954
R15735 VSS.n6925 VSS.n2748 338.954
R15736 VSS.n3209 VSS.n3208 338.954
R15737 VSS.n3256 VSS.n3254 338.954
R15738 VSS.n3325 VSS.n2791 338.954
R15739 VSS.n3326 VSS.n2779 338.954
R15740 VSS.n3354 VSS.n3352 338.954
R15741 VSS.n9169 VSS.n9168 338.954
R15742 VSS.n9216 VSS.n9214 338.954
R15743 VSS.n9285 VSS.n58 338.954
R15744 VSS.n9286 VSS.n46 338.954
R15745 VSS.n9314 VSS.n9312 338.954
R15746 VSS.n8995 VSS.n8994 338.954
R15747 VSS.n8834 VSS.n8824 338.954
R15748 VSS.n8913 VSS.n8847 338.954
R15749 VSS.n8914 VSS.n8902 338.954
R15750 VSS.n8923 VSS.n8921 338.954
R15751 VSS.n813 VSS.n812 338.954
R15752 VSS.n795 VSS.n648 338.954
R15753 VSS.n743 VSS.n729 338.954
R15754 VSS.n744 VSS.n30 338.954
R15755 VSS.n9335 VSS.n9334 338.954
R15756 VSS.n7694 VSS.n7372 332.558
R15757 VSS.n7695 VSS.n7694 332.558
R15758 VSS.n8286 VSS.n7786 332.558
R15759 VSS.n8287 VSS.n8286 332.558
R15760 VSS.n1625 VSS.n1624 332.558
R15761 VSS.n1624 VSS.n1503 332.558
R15762 VSS.n2217 VSS.n2216 332.558
R15763 VSS.n2216 VSS.n2076 332.558
R15764 VSS.n3896 VSS.n3396 332.558
R15765 VSS.n3897 VSS.n3896 332.558
R15766 VSS.n4488 VSS.n3988 332.558
R15767 VSS.n4489 VSS.n4488 332.558
R15768 VSS.n5080 VSS.n4580 332.558
R15769 VSS.n5081 VSS.n5080 332.558
R15770 VSS.n5672 VSS.n5172 332.558
R15771 VSS.n5673 VSS.n5672 332.558
R15772 VSS.n6264 VSS.n5764 332.558
R15773 VSS.n6265 VSS.n6264 332.558
R15774 VSS.n6856 VSS.n6356 332.558
R15775 VSS.n6857 VSS.n6856 332.558
R15776 VSS.n6961 VSS.n6960 332.558
R15777 VSS.n6960 VSS.n2674 332.558
R15778 VSS.n3304 VSS.n2803 332.558
R15779 VSS.n3305 VSS.n3304 332.558
R15780 VSS.n9264 VSS.n70 332.558
R15781 VSS.n9265 VSS.n9264 332.558
R15782 VSS.n8959 VSS.n8846 332.558
R15783 VSS.n8959 VSS.n8958 332.558
R15784 VSS.n780 VSS.n779 332.558
R15785 VSS.n779 VSS.n666 332.558
R15786 VSS.n7509 VSS.n7453 329.38
R15787 VSS.n7532 VSS.n7530 329.38
R15788 VSS.n7532 VSS.n7531 329.38
R15789 VSS.n7561 VSS.n7560 329.38
R15790 VSS.n7582 VSS.n7417 329.38
R15791 VSS.n8101 VSS.n7867 329.38
R15792 VSS.n8124 VSS.n8122 329.38
R15793 VSS.n8124 VSS.n8123 329.38
R15794 VSS.n8153 VSS.n8152 329.38
R15795 VSS.n8174 VSS.n7831 329.38
R15796 VSS.n8569 VSS.n8565 329.38
R15797 VSS.n8567 VSS.n234 329.38
R15798 VSS.n8598 VSS.n234 329.38
R15799 VSS.n8602 VSS.n8601 329.38
R15800 VSS.n8631 VSS.n8630 329.38
R15801 VSS.n1409 VSS.n1408 329.38
R15802 VSS.n1416 VSS.n1415 329.38
R15803 VSS.n1417 VSS.n1416 329.38
R15804 VSS.n1433 VSS.n1432 329.38
R15805 VSS.n1448 VSS.n1361 329.38
R15806 VSS.n1251 VSS.n1247 329.38
R15807 VSS.n1249 VSS.n1180 329.38
R15808 VSS.n1280 VSS.n1180 329.38
R15809 VSS.n1284 VSS.n1283 329.38
R15810 VSS.n1313 VSS.n1312 329.38
R15811 VSS.n1982 VSS.n1981 329.38
R15812 VSS.n1989 VSS.n1988 329.38
R15813 VSS.n1990 VSS.n1989 329.38
R15814 VSS.n2006 VSS.n2005 329.38
R15815 VSS.n2021 VSS.n1934 329.38
R15816 VSS.n1824 VSS.n1820 329.38
R15817 VSS.n1822 VSS.n1753 329.38
R15818 VSS.n1853 VSS.n1753 329.38
R15819 VSS.n1857 VSS.n1856 329.38
R15820 VSS.n1886 VSS.n1885 329.38
R15821 VSS.n3711 VSS.n3477 329.38
R15822 VSS.n3734 VSS.n3732 329.38
R15823 VSS.n3734 VSS.n3733 329.38
R15824 VSS.n3763 VSS.n3762 329.38
R15825 VSS.n3784 VSS.n3441 329.38
R15826 VSS.n3618 VSS.n3614 329.38
R15827 VSS.n3616 VSS.n3547 329.38
R15828 VSS.n3647 VSS.n3547 329.38
R15829 VSS.n3651 VSS.n3650 329.38
R15830 VSS.n3680 VSS.n3679 329.38
R15831 VSS.n4303 VSS.n4069 329.38
R15832 VSS.n4326 VSS.n4324 329.38
R15833 VSS.n4326 VSS.n4325 329.38
R15834 VSS.n4355 VSS.n4354 329.38
R15835 VSS.n4376 VSS.n4033 329.38
R15836 VSS.n4210 VSS.n4206 329.38
R15837 VSS.n4208 VSS.n4139 329.38
R15838 VSS.n4239 VSS.n4139 329.38
R15839 VSS.n4243 VSS.n4242 329.38
R15840 VSS.n4272 VSS.n4271 329.38
R15841 VSS.n4895 VSS.n4661 329.38
R15842 VSS.n4918 VSS.n4916 329.38
R15843 VSS.n4918 VSS.n4917 329.38
R15844 VSS.n4947 VSS.n4946 329.38
R15845 VSS.n4968 VSS.n4625 329.38
R15846 VSS.n4802 VSS.n4798 329.38
R15847 VSS.n4800 VSS.n4731 329.38
R15848 VSS.n4831 VSS.n4731 329.38
R15849 VSS.n4835 VSS.n4834 329.38
R15850 VSS.n4864 VSS.n4863 329.38
R15851 VSS.n5487 VSS.n5253 329.38
R15852 VSS.n5510 VSS.n5508 329.38
R15853 VSS.n5510 VSS.n5509 329.38
R15854 VSS.n5539 VSS.n5538 329.38
R15855 VSS.n5560 VSS.n5217 329.38
R15856 VSS.n5394 VSS.n5390 329.38
R15857 VSS.n5392 VSS.n5323 329.38
R15858 VSS.n5423 VSS.n5323 329.38
R15859 VSS.n5427 VSS.n5426 329.38
R15860 VSS.n5456 VSS.n5455 329.38
R15861 VSS.n6079 VSS.n5845 329.38
R15862 VSS.n6102 VSS.n6100 329.38
R15863 VSS.n6102 VSS.n6101 329.38
R15864 VSS.n6131 VSS.n6130 329.38
R15865 VSS.n6152 VSS.n5809 329.38
R15866 VSS.n5986 VSS.n5982 329.38
R15867 VSS.n5984 VSS.n5915 329.38
R15868 VSS.n6015 VSS.n5915 329.38
R15869 VSS.n6019 VSS.n6018 329.38
R15870 VSS.n6048 VSS.n6047 329.38
R15871 VSS.n6671 VSS.n6437 329.38
R15872 VSS.n6694 VSS.n6692 329.38
R15873 VSS.n6694 VSS.n6693 329.38
R15874 VSS.n6723 VSS.n6722 329.38
R15875 VSS.n6744 VSS.n6401 329.38
R15876 VSS.n6578 VSS.n6574 329.38
R15877 VSS.n6576 VSS.n6507 329.38
R15878 VSS.n6607 VSS.n6507 329.38
R15879 VSS.n6611 VSS.n6610 329.38
R15880 VSS.n6640 VSS.n6639 329.38
R15881 VSS.n2580 VSS.n2579 329.38
R15882 VSS.n2587 VSS.n2586 329.38
R15883 VSS.n2588 VSS.n2587 329.38
R15884 VSS.n2604 VSS.n2603 329.38
R15885 VSS.n2619 VSS.n2532 329.38
R15886 VSS.n2422 VSS.n2418 329.38
R15887 VSS.n2420 VSS.n2351 329.38
R15888 VSS.n2451 VSS.n2351 329.38
R15889 VSS.n2455 VSS.n2454 329.38
R15890 VSS.n2484 VSS.n2483 329.38
R15891 VSS.n3119 VSS.n2884 329.38
R15892 VSS.n3142 VSS.n3140 329.38
R15893 VSS.n3142 VSS.n3141 329.38
R15894 VSS.n3171 VSS.n3170 329.38
R15895 VSS.n3192 VSS.n2848 329.38
R15896 VSS.n3014 VSS.n2961 329.38
R15897 VSS.n3037 VSS.n3035 329.38
R15898 VSS.n3037 VSS.n3036 329.38
R15899 VSS.n3066 VSS.n3065 329.38
R15900 VSS.n3088 VSS.n2923 329.38
R15901 VSS.n9079 VSS.n151 329.38
R15902 VSS.n9102 VSS.n9100 329.38
R15903 VSS.n9102 VSS.n9101 329.38
R15904 VSS.n9131 VSS.n9130 329.38
R15905 VSS.n9152 VSS.n115 329.38
R15906 VSS.n357 VSS.n324 329.38
R15907 VSS.n359 VSS.n320 329.38
R15908 VSS.n366 VSS.n320 329.38
R15909 VSS.n368 VSS.n314 329.38
R15910 VSS.n385 VSS.n384 329.38
R15911 VSS.n8727 VSS.n8726 329.38
R15912 VSS.n8734 VSS.n8733 329.38
R15913 VSS.n8735 VSS.n8734 329.38
R15914 VSS.n8751 VSS.n8750 329.38
R15915 VSS.n8766 VSS.n8679 329.38
R15916 VSS.n572 VSS.n571 329.38
R15917 VSS.n579 VSS.n578 329.38
R15918 VSS.n580 VSS.n579 329.38
R15919 VSS.n596 VSS.n595 329.38
R15920 VSS.n611 VSS.n521 329.38
R15921 VSS.n915 VSS.n914 329.38
R15922 VSS.n922 VSS.n921 329.38
R15923 VSS.n923 VSS.n922 329.38
R15924 VSS.n939 VSS.n938 329.38
R15925 VSS.n955 VSS.n868 329.38
R15926 VSS.n1096 VSS.n1095 329.38
R15927 VSS.n1103 VSS.n1102 329.38
R15928 VSS.n1104 VSS.n1103 329.38
R15929 VSS.n1120 VSS.n1119 329.38
R15930 VSS.n1136 VSS.n1049 329.38
R15931 VSS.t75 VSS.n7194 304.498
R15932 VSS.n7693 VSS.n7692 292.5
R15933 VSS.n7694 VSS.n7693 292.5
R15934 VSS.n8285 VSS.n8284 292.5
R15935 VSS.n8286 VSS.n8285 292.5
R15936 VSS.n1623 VSS.n1622 292.5
R15937 VSS.n1624 VSS.n1623 292.5
R15938 VSS.n2215 VSS.n2214 292.5
R15939 VSS.n2216 VSS.n2215 292.5
R15940 VSS.n3895 VSS.n3894 292.5
R15941 VSS.n3896 VSS.n3895 292.5
R15942 VSS.n4487 VSS.n4486 292.5
R15943 VSS.n4488 VSS.n4487 292.5
R15944 VSS.n5079 VSS.n5078 292.5
R15945 VSS.n5080 VSS.n5079 292.5
R15946 VSS.n5671 VSS.n5670 292.5
R15947 VSS.n5672 VSS.n5671 292.5
R15948 VSS.n6263 VSS.n6262 292.5
R15949 VSS.n6264 VSS.n6263 292.5
R15950 VSS.n6855 VSS.n6854 292.5
R15951 VSS.n6856 VSS.n6855 292.5
R15952 VSS.n6959 VSS.n6958 292.5
R15953 VSS.n6960 VSS.n6959 292.5
R15954 VSS.n3303 VSS.n3302 292.5
R15955 VSS.n3304 VSS.n3303 292.5
R15956 VSS.n9263 VSS.n9262 292.5
R15957 VSS.n9264 VSS.n9263 292.5
R15958 VSS.n8961 VSS.n8960 292.5
R15959 VSS.n8960 VSS.n8959 292.5
R15960 VSS.n778 VSS.n777 292.5
R15961 VSS.n779 VSS.n778 292.5
R15962 VSS.n8387 VSS.n8386 292.5
R15963 VSS.n8388 VSS.n8387 292.5
R15964 VSS.n7602 VSS.n7601 290.906
R15965 VSS.n7745 VSS.n7344 290.906
R15966 VSS.n8194 VSS.n8193 290.906
R15967 VSS.n8337 VSS.n7758 290.906
R15968 VSS.n8998 VSS.n8997 290.906
R15969 VSS.n8925 VSS.n8899 290.906
R15970 VSS.n1661 VSS.n1660 290.906
R15971 VSS.n9345 VSS.n6 290.906
R15972 VSS.n2253 VSS.n2252 290.906
R15973 VSS.n2159 VSS.n2158 290.906
R15974 VSS.n3804 VSS.n3803 290.906
R15975 VSS.n3948 VSS.n3369 290.906
R15976 VSS.n4396 VSS.n4395 290.906
R15977 VSS.n4540 VSS.n3961 290.906
R15978 VSS.n4988 VSS.n4987 290.906
R15979 VSS.n5132 VSS.n4553 290.906
R15980 VSS.n5580 VSS.n5579 290.906
R15981 VSS.n5724 VSS.n5145 290.906
R15982 VSS.n6172 VSS.n6171 290.906
R15983 VSS.n6316 VSS.n5737 290.906
R15984 VSS.n6764 VSS.n6763 290.906
R15985 VSS.n6908 VSS.n6329 290.906
R15986 VSS.n6997 VSS.n6996 290.906
R15987 VSS.n2757 VSS.n2756 290.906
R15988 VSS.n3212 VSS.n3211 290.906
R15989 VSS.n3356 VSS.n2776 290.906
R15990 VSS.n9172 VSS.n9171 290.906
R15991 VSS.n9316 VSS.n43 290.906
R15992 VSS.n816 VSS.n815 290.906
R15993 VSS.n9338 VSS.n9337 290.906
R15994 VSS.n8425 VSS.n8424 290.906
R15995 VSS.n7325 VSS.n7324 290.906
R15996 VSS.n8427 VSS.t73 269.807
R15997 VSS.n7591 VSS.t78 255.815
R15998 VSS.n8183 VSS.t225 255.815
R15999 VSS.t113 VSS.n1455 255.815
R16000 VSS.t176 VSS.n2028 255.815
R16001 VSS.n3793 VSS.t251 255.815
R16002 VSS.n4385 VSS.t230 255.815
R16003 VSS.n4977 VSS.t117 255.815
R16004 VSS.n5569 VSS.t305 255.815
R16005 VSS.n6161 VSS.t277 255.815
R16006 VSS.n6753 VSS.t98 255.815
R16007 VSS.t195 VSS.n2626 255.815
R16008 VSS.n3201 VSS.t31 255.815
R16009 VSS.n9161 VSS.t39 255.815
R16010 VSS.t34 VSS.n8773 255.815
R16011 VSS.t257 VSS.n618 255.815
R16012 VSS.t160 VSS.n7118 239.457
R16013 VSS.n7507 VSS.t288 198.87
R16014 VSS.n8099 VSS.t221 198.87
R16015 VSS.t164 VSS.n1379 198.87
R16016 VSS.t21 VSS.n1952 198.87
R16017 VSS.n3709 VSS.t199 198.87
R16018 VSS.n4301 VSS.t239 198.87
R16019 VSS.n4893 VSS.t167 198.87
R16020 VSS.n5485 VSS.t209 198.87
R16021 VSS.n6077 VSS.t186 198.87
R16022 VSS.n6669 VSS.t298 198.87
R16023 VSS.t202 VSS.n2550 198.87
R16024 VSS.n3117 VSS.t59 198.87
R16025 VSS.n9077 VSS.t110 198.87
R16026 VSS.t146 VSS.n8697 198.87
R16027 VSS.t255 VSS.n539 198.87
R16028 VSS.t8 VSS.n257 192.655
R16029 VSS.t52 VSS.n1203 192.655
R16030 VSS.t68 VSS.n1776 192.655
R16031 VSS.t61 VSS.n3570 192.655
R16032 VSS.t149 VSS.n4162 192.655
R16033 VSS.t65 VSS.n4754 192.655
R16034 VSS.t82 VSS.n5346 192.655
R16035 VSS.t295 VSS.n5938 192.655
R16036 VSS.t192 VSS.n6530 192.655
R16037 VSS.t233 VSS.n2374 192.655
R16038 VSS.n3012 VSS.t216 192.655
R16039 VSS.n344 VSS.t309 192.655
R16040 VSS.t268 VSS.n887 192.655
R16041 VSS.t19 VSS.n1068 192.655
R16042 VSS.n7604 VSS.t80 188.758
R16043 VSS.n8196 VSS.t227 188.758
R16044 VSS.n1663 VSS.t115 188.758
R16045 VSS.n2255 VSS.t178 188.758
R16046 VSS.n3806 VSS.t253 188.758
R16047 VSS.n4398 VSS.t228 188.758
R16048 VSS.n4990 VSS.t119 188.758
R16049 VSS.n5582 VSS.t307 188.758
R16050 VSS.n6174 VSS.t279 188.758
R16051 VSS.n6766 VSS.t100 188.758
R16052 VSS.n6999 VSS.t197 188.758
R16053 VSS.n3214 VSS.t33 188.758
R16054 VSS.n9174 VSS.t41 188.758
R16055 VSS.n9000 VSS.t36 188.758
R16056 VSS.n818 VSS.t259 188.758
R16057 VSS.n7120 VSS.t160 157.143
R16058 VSS.n8537 VSS.t8 136.724
R16059 VSS.n1219 VSS.t52 136.724
R16060 VSS.n1792 VSS.t68 136.724
R16061 VSS.n3586 VSS.t61 136.724
R16062 VSS.n4178 VSS.t149 136.724
R16063 VSS.n4770 VSS.t65 136.724
R16064 VSS.n5362 VSS.t82 136.724
R16065 VSS.n5954 VSS.t295 136.724
R16066 VSS.n6546 VSS.t192 136.724
R16067 VSS.n2390 VSS.t233 136.724
R16068 VSS.n2987 VSS.t216 136.724
R16069 VSS.t309 VSS.n343 136.724
R16070 VSS.n889 VSS.t268 136.724
R16071 VSS.n1070 VSS.t19 136.724
R16072 VSS.n7481 VSS.t288 130.508
R16073 VSS.n7895 VSS.t221 130.508
R16074 VSS.n1381 VSS.t164 130.508
R16075 VSS.n1954 VSS.t21 130.508
R16076 VSS.n3505 VSS.t199 130.508
R16077 VSS.n4097 VSS.t239 130.508
R16078 VSS.n4689 VSS.t167 130.508
R16079 VSS.n5281 VSS.t209 130.508
R16080 VSS.n5873 VSS.t186 130.508
R16081 VSS.n6465 VSS.t298 130.508
R16082 VSS.n2552 VSS.t202 130.508
R16083 VSS.n2912 VSS.t59 130.508
R16084 VSS.n184 VSS.t110 130.508
R16085 VSS.n8699 VSS.t146 130.508
R16086 VSS.n546 VSS.t255 130.508
R16087 VSS.n8008 VSS.n8004 128.415
R16088 VSS.n8006 VSS.n7937 128.415
R16089 VSS.n8037 VSS.n7937 128.415
R16090 VSS.n8041 VSS.n8040 128.415
R16091 VSS.n8070 VSS.n8069 128.415
R16092 VSS.n8390 VSS.n8389 121.799
R16093 VSS.n7307 VSS.n7242 121.799
R16094 VSS.n7154 VSS.n7113 112.246
R16095 VSS.n7156 VSS.n7109 112.246
R16096 VSS.n8405 VSS.n8404 106.575
R16097 VSS.t301 VSS.n7296 106.575
R16098 VSS.n7645 VSS.n7372 102.326
R16099 VSS.n7696 VSS.n7695 102.326
R16100 VSS.n8237 VSS.n7786 102.326
R16101 VSS.n8288 VSS.n8287 102.326
R16102 VSS.n1626 VSS.n1625 102.326
R16103 VSS.n1581 VSS.n1503 102.326
R16104 VSS.n2218 VSS.n2217 102.326
R16105 VSS.n2141 VSS.n2076 102.326
R16106 VSS.n3847 VSS.n3396 102.326
R16107 VSS.n3898 VSS.n3897 102.326
R16108 VSS.n4439 VSS.n3988 102.326
R16109 VSS.n4490 VSS.n4489 102.326
R16110 VSS.n5031 VSS.n4580 102.326
R16111 VSS.n5082 VSS.n5081 102.326
R16112 VSS.n5623 VSS.n5172 102.326
R16113 VSS.n5674 VSS.n5673 102.326
R16114 VSS.n6215 VSS.n5764 102.326
R16115 VSS.n6266 VSS.n6265 102.326
R16116 VSS.n6807 VSS.n6356 102.326
R16117 VSS.n6858 VSS.n6857 102.326
R16118 VSS.n6962 VSS.n6961 102.326
R16119 VSS.n2739 VSS.n2674 102.326
R16120 VSS.n3255 VSS.n2803 102.326
R16121 VSS.n3306 VSS.n3305 102.326
R16122 VSS.n9215 VSS.n70 102.326
R16123 VSS.n9266 VSS.n9265 102.326
R16124 VSS.n8846 VSS.n8845 102.326
R16125 VSS.n8958 VSS.n8957 102.326
R16126 VSS.n781 VSS.n780 102.326
R16127 VSS.n739 VSS.n666 102.326
R16128 VSS.n8406 VSS.t75 98.9624
R16129 VSS.n7147 VSS.n7146 97.2794
R16130 VSS.t285 VSS.n7172 97.2794
R16131 VSS.n7530 VSS.n7529 93.2208
R16132 VSS.n7531 VSS.n7432 93.2208
R16133 VSS.n8122 VSS.n8121 93.2208
R16134 VSS.n8123 VSS.n7846 93.2208
R16135 VSS.n8568 VSS.n8567 93.2208
R16136 VSS.n8599 VSS.n8598 93.2208
R16137 VSS.n1415 VSS.n1374 93.2208
R16138 VSS.n1417 VSS.n1370 93.2208
R16139 VSS.n1250 VSS.n1249 93.2208
R16140 VSS.n1281 VSS.n1280 93.2208
R16141 VSS.n1988 VSS.n1947 93.2208
R16142 VSS.n1990 VSS.n1943 93.2208
R16143 VSS.n1823 VSS.n1822 93.2208
R16144 VSS.n1854 VSS.n1853 93.2208
R16145 VSS.n3732 VSS.n3731 93.2208
R16146 VSS.n3733 VSS.n3456 93.2208
R16147 VSS.n3617 VSS.n3616 93.2208
R16148 VSS.n3648 VSS.n3647 93.2208
R16149 VSS.n4324 VSS.n4323 93.2208
R16150 VSS.n4325 VSS.n4048 93.2208
R16151 VSS.n4209 VSS.n4208 93.2208
R16152 VSS.n4240 VSS.n4239 93.2208
R16153 VSS.n4916 VSS.n4915 93.2208
R16154 VSS.n4917 VSS.n4640 93.2208
R16155 VSS.n4801 VSS.n4800 93.2208
R16156 VSS.n4832 VSS.n4831 93.2208
R16157 VSS.n5508 VSS.n5507 93.2208
R16158 VSS.n5509 VSS.n5232 93.2208
R16159 VSS.n5393 VSS.n5392 93.2208
R16160 VSS.n5424 VSS.n5423 93.2208
R16161 VSS.n6100 VSS.n6099 93.2208
R16162 VSS.n6101 VSS.n5824 93.2208
R16163 VSS.n5985 VSS.n5984 93.2208
R16164 VSS.n6016 VSS.n6015 93.2208
R16165 VSS.n6692 VSS.n6691 93.2208
R16166 VSS.n6693 VSS.n6416 93.2208
R16167 VSS.n6577 VSS.n6576 93.2208
R16168 VSS.n6608 VSS.n6607 93.2208
R16169 VSS.n2586 VSS.n2545 93.2208
R16170 VSS.n2588 VSS.n2541 93.2208
R16171 VSS.n2421 VSS.n2420 93.2208
R16172 VSS.n2452 VSS.n2451 93.2208
R16173 VSS.n3140 VSS.n3139 93.2208
R16174 VSS.n3141 VSS.n2863 93.2208
R16175 VSS.n3035 VSS.n3034 93.2208
R16176 VSS.n3036 VSS.n2938 93.2208
R16177 VSS.n9100 VSS.n9099 93.2208
R16178 VSS.n9101 VSS.n130 93.2208
R16179 VSS.n359 VSS.n358 93.2208
R16180 VSS.n367 VSS.n366 93.2208
R16181 VSS.n8733 VSS.n8692 93.2208
R16182 VSS.n8735 VSS.n8688 93.2208
R16183 VSS.n578 VSS.n534 93.2208
R16184 VSS.n580 VSS.n530 93.2208
R16185 VSS.n921 VSS.n882 93.2208
R16186 VSS.n923 VSS.n877 93.2208
R16187 VSS.n1102 VSS.n1063 93.2208
R16188 VSS.n1104 VSS.n1058 93.2208
R16189 VSS.n8420 VSS.n7194 91.35
R16190 VSS.n8355 VSS.n8354 91.35
R16191 VSS.n7644 VSS.n7643 89.5354
R16192 VSS.t313 VSS.n7715 89.5354
R16193 VSS.n8236 VSS.n8235 89.5354
R16194 VSS.t47 VSS.n8307 89.5354
R16195 VSS.n1641 VSS.n1640 89.5354
R16196 VSS.t92 VSS.n1570 89.5354
R16197 VSS.n2233 VSS.n2232 89.5354
R16198 VSS.t244 VSS.n2130 89.5354
R16199 VSS.n3846 VSS.n3845 89.5354
R16200 VSS.t15 VSS.n3917 89.5354
R16201 VSS.n4438 VSS.n4437 89.5354
R16202 VSS.t120 VSS.n4509 89.5354
R16203 VSS.n5030 VSS.n5029 89.5354
R16204 VSS.t272 VSS.n5101 89.5354
R16205 VSS.n5622 VSS.n5621 89.5354
R16206 VSS.t106 VSS.n5693 89.5354
R16207 VSS.n6214 VSS.n6213 89.5354
R16208 VSS.t281 VSS.n6285 89.5354
R16209 VSS.n6806 VSS.n6805 89.5354
R16210 VSS.t205 VSS.n6877 89.5354
R16211 VSS.n6977 VSS.n6976 89.5354
R16212 VSS.t55 VSS.n2728 89.5354
R16213 VSS.n3254 VSS.n3253 89.5354
R16214 VSS.t4 VSS.n3325 89.5354
R16215 VSS.n9214 VSS.n9213 89.5354
R16216 VSS.t290 VSS.n9285 89.5354
R16217 VSS.n8834 VSS.n8833 89.5354
R16218 VSS.t142 VSS.n8913 89.5354
R16219 VSS.n796 VSS.n795 89.5354
R16220 VSS.t102 VSS.n743 89.5354
R16221 VSS.t78 VSS.n7394 83.14
R16222 VSS.t225 VSS.n7808 83.14
R16223 VSS.n1642 VSS.t113 83.14
R16224 VSS.n2234 VSS.t176 83.14
R16225 VSS.t251 VSS.n3418 83.14
R16226 VSS.t230 VSS.n4010 83.14
R16227 VSS.t117 VSS.n4602 83.14
R16228 VSS.t305 VSS.n5194 83.14
R16229 VSS.t277 VSS.n5786 83.14
R16230 VSS.t98 VSS.n6378 83.14
R16231 VSS.n6978 VSS.t195 83.14
R16232 VSS.t31 VSS.n2825 83.14
R16233 VSS.t39 VSS.n92 83.14
R16234 VSS.n8832 VSS.t34 83.14
R16235 VSS.n797 VSS.t257 83.14
R16236 VSS.n7120 VSS.n7057 82.3134
R16237 VSS.n7188 VSS.n7187 82.3134
R16238 VSS.n7600 VSS.n7590 81.5708
R16239 VSS.n7592 VSS.n7395 81.5708
R16240 VSS.n7647 VSS.n7392 81.5708
R16241 VSS.n7714 VSS.n7361 81.5708
R16242 VSS.n7717 VSS.n7348 81.5708
R16243 VSS.n7744 VSS.n7345 81.5708
R16244 VSS.n8192 VSS.n8182 81.5708
R16245 VSS.n8184 VSS.n7809 81.5708
R16246 VSS.n8239 VSS.n7806 81.5708
R16247 VSS.n8306 VSS.n7775 81.5708
R16248 VSS.n8309 VSS.n7762 81.5708
R16249 VSS.n8336 VSS.n7759 81.5708
R16250 VSS.n8996 VSS.n8772 81.5708
R16251 VSS.n8831 VSS.n8774 81.5708
R16252 VSS.n8836 VSS.n8835 81.5708
R16253 VSS.n8912 VSS.n8848 81.5708
R16254 VSS.n8916 VSS.n8915 81.5708
R16255 VSS.n8924 VSS.n8900 81.5708
R16256 VSS.n1659 VSS.n1454 81.5708
R16257 VSS.n1643 VSS.n1456 81.5708
R16258 VSS.n1639 VSS.n1486 81.5708
R16259 VSS.n1584 VSS.n1583 81.5708
R16260 VSS.n1592 VSS.n1568 81.5708
R16261 VSS.n9344 VSS.n7 81.5708
R16262 VSS.n2251 VSS.n2027 81.5708
R16263 VSS.n2235 VSS.n2029 81.5708
R16264 VSS.n2231 VSS.n2059 81.5708
R16265 VSS.n2144 VSS.n2143 81.5708
R16266 VSS.n2184 VSS.n2128 81.5708
R16267 VSS.n2180 VSS.n2151 81.5708
R16268 VSS.n3802 VSS.n3792 81.5708
R16269 VSS.n3794 VSS.n3419 81.5708
R16270 VSS.n3849 VSS.n3416 81.5708
R16271 VSS.n3916 VSS.n3385 81.5708
R16272 VSS.n3919 VSS.n3373 81.5708
R16273 VSS.n3947 VSS.n3370 81.5708
R16274 VSS.n4394 VSS.n4384 81.5708
R16275 VSS.n4386 VSS.n4011 81.5708
R16276 VSS.n4441 VSS.n4008 81.5708
R16277 VSS.n4508 VSS.n3977 81.5708
R16278 VSS.n4511 VSS.n3965 81.5708
R16279 VSS.n4539 VSS.n3962 81.5708
R16280 VSS.n4986 VSS.n4976 81.5708
R16281 VSS.n4978 VSS.n4603 81.5708
R16282 VSS.n5033 VSS.n4600 81.5708
R16283 VSS.n5100 VSS.n4569 81.5708
R16284 VSS.n5103 VSS.n4557 81.5708
R16285 VSS.n5131 VSS.n4554 81.5708
R16286 VSS.n5578 VSS.n5568 81.5708
R16287 VSS.n5570 VSS.n5195 81.5708
R16288 VSS.n5625 VSS.n5192 81.5708
R16289 VSS.n5692 VSS.n5161 81.5708
R16290 VSS.n5695 VSS.n5149 81.5708
R16291 VSS.n5723 VSS.n5146 81.5708
R16292 VSS.n6170 VSS.n6160 81.5708
R16293 VSS.n6162 VSS.n5787 81.5708
R16294 VSS.n6217 VSS.n5784 81.5708
R16295 VSS.n6284 VSS.n5753 81.5708
R16296 VSS.n6287 VSS.n5741 81.5708
R16297 VSS.n6315 VSS.n5738 81.5708
R16298 VSS.n6762 VSS.n6752 81.5708
R16299 VSS.n6754 VSS.n6379 81.5708
R16300 VSS.n6809 VSS.n6376 81.5708
R16301 VSS.n6876 VSS.n6345 81.5708
R16302 VSS.n6879 VSS.n6333 81.5708
R16303 VSS.n6907 VSS.n6330 81.5708
R16304 VSS.n6995 VSS.n2625 81.5708
R16305 VSS.n6979 VSS.n2627 81.5708
R16306 VSS.n6975 VSS.n2657 81.5708
R16307 VSS.n2742 VSS.n2741 81.5708
R16308 VSS.n6928 VSS.n2726 81.5708
R16309 VSS.n6924 VSS.n2749 81.5708
R16310 VSS.n3210 VSS.n3200 81.5708
R16311 VSS.n3202 VSS.n2826 81.5708
R16312 VSS.n3257 VSS.n2823 81.5708
R16313 VSS.n3324 VSS.n2792 81.5708
R16314 VSS.n3327 VSS.n2780 81.5708
R16315 VSS.n3355 VSS.n2777 81.5708
R16316 VSS.n9170 VSS.n9160 81.5708
R16317 VSS.n9162 VSS.n93 81.5708
R16318 VSS.n9217 VSS.n90 81.5708
R16319 VSS.n9284 VSS.n59 81.5708
R16320 VSS.n9287 VSS.n47 81.5708
R16321 VSS.n9315 VSS.n44 81.5708
R16322 VSS.n814 VSS.n617 81.5708
R16323 VSS.n798 VSS.n619 81.5708
R16324 VSS.n794 VSS.n649 81.5708
R16325 VSS.n742 VSS.n741 81.5708
R16326 VSS.n745 VSS.n31 81.5708
R16327 VSS.n9336 VSS.n29 81.5708
R16328 VSS.n8423 VSS.n7193 81.5708
R16329 VSS.n8407 VSS.n7195 81.5708
R16330 VSS.n8403 VSS.n7225 81.5708
R16331 VSS.n7310 VSS.n7309 81.5708
R16332 VSS.n8356 VSS.n7294 81.5708
R16333 VSS.n8352 VSS.n7317 81.5708
R16334 VSS.n7509 VSS.n7508 80.7915
R16335 VSS.t71 VSS.n7561 80.7915
R16336 VSS.n8101 VSS.n8100 80.7915
R16337 VSS.t125 VSS.n8153 80.7915
R16338 VSS.n8565 VSS.n8564 80.7915
R16339 VSS.n8601 VSS.n8600 80.7915
R16340 VSS.n1408 VSS.n1407 80.7915
R16341 VSS.t139 VSS.n1433 80.7915
R16342 VSS.n1247 VSS.n1246 80.7915
R16343 VSS.n1283 VSS.n1282 80.7915
R16344 VSS.n1981 VSS.n1980 80.7915
R16345 VSS.t172 VSS.n2006 80.7915
R16346 VSS.n1820 VSS.n1819 80.7915
R16347 VSS.n1856 VSS.n1855 80.7915
R16348 VSS.n3711 VSS.n3710 80.7915
R16349 VSS.t248 VSS.n3763 80.7915
R16350 VSS.n3614 VSS.n3613 80.7915
R16351 VSS.n3650 VSS.n3649 80.7915
R16352 VSS.n4303 VSS.n4302 80.7915
R16353 VSS.t170 VSS.n4355 80.7915
R16354 VSS.n4206 VSS.n4205 80.7915
R16355 VSS.n4242 VSS.n4241 80.7915
R16356 VSS.n4895 VSS.n4894 80.7915
R16357 VSS.t127 VSS.n4947 80.7915
R16358 VSS.n4798 VSS.n4797 80.7915
R16359 VSS.n4834 VSS.n4833 80.7915
R16360 VSS.n5487 VSS.n5486 80.7915
R16361 VSS.t96 VSS.n5539 80.7915
R16362 VSS.n5390 VSS.n5389 80.7915
R16363 VSS.n5426 VSS.n5425 80.7915
R16364 VSS.n6079 VSS.n6078 80.7915
R16365 VSS.t188 VSS.n6131 80.7915
R16366 VSS.n5982 VSS.n5981 80.7915
R16367 VSS.n6018 VSS.n6017 80.7915
R16368 VSS.n6671 VSS.n6670 80.7915
R16369 VSS.t236 VSS.n6723 80.7915
R16370 VSS.n6574 VSS.n6573 80.7915
R16371 VSS.n6610 VSS.n6609 80.7915
R16372 VSS.n2579 VSS.n2578 80.7915
R16373 VSS.t151 VSS.n2604 80.7915
R16374 VSS.n2418 VSS.n2417 80.7915
R16375 VSS.n2454 VSS.n2453 80.7915
R16376 VSS.n3119 VSS.n3118 80.7915
R16377 VSS.t24 VSS.n3171 80.7915
R16378 VSS.n3014 VSS.n3013 80.7915
R16379 VSS.n3067 VSS.n3066 80.7915
R16380 VSS.n9079 VSS.n9078 80.7915
R16381 VSS.t218 VSS.n9131 80.7915
R16382 VSS.n345 VSS.n324 80.7915
R16383 VSS.n383 VSS.n314 80.7915
R16384 VSS.n8726 VSS.n8725 80.7915
R16385 VSS.t262 VSS.n8751 80.7915
R16386 VSS.n571 VSS.n570 80.7915
R16387 VSS.t27 VSS.n596 80.7915
R16388 VSS.n914 VSS.n913 80.7915
R16389 VSS.n940 VSS.n939 80.7915
R16390 VSS.n1095 VSS.n1094 80.7915
R16391 VSS.n1121 VSS.n1120 80.7915
R16392 VSS.n7693 VSS.n7373 80.0317
R16393 VSS.n7693 VSS.n7371 80.0317
R16394 VSS.n8285 VSS.n7787 80.0317
R16395 VSS.n8285 VSS.n7785 80.0317
R16396 VSS.n8960 VSS.n8822 80.0317
R16397 VSS.n8960 VSS.n8823 80.0317
R16398 VSS.n1623 VSS.n1502 80.0317
R16399 VSS.n1623 VSS.n1504 80.0317
R16400 VSS.n2215 VSS.n2075 80.0317
R16401 VSS.n2215 VSS.n2077 80.0317
R16402 VSS.n3895 VSS.n3397 80.0317
R16403 VSS.n3895 VSS.n3395 80.0317
R16404 VSS.n4487 VSS.n3989 80.0317
R16405 VSS.n4487 VSS.n3987 80.0317
R16406 VSS.n5079 VSS.n4581 80.0317
R16407 VSS.n5079 VSS.n4579 80.0317
R16408 VSS.n5671 VSS.n5173 80.0317
R16409 VSS.n5671 VSS.n5171 80.0317
R16410 VSS.n6263 VSS.n5765 80.0317
R16411 VSS.n6263 VSS.n5763 80.0317
R16412 VSS.n6855 VSS.n6357 80.0317
R16413 VSS.n6855 VSS.n6355 80.0317
R16414 VSS.n6959 VSS.n2673 80.0317
R16415 VSS.n6959 VSS.n2675 80.0317
R16416 VSS.n3303 VSS.n2804 80.0317
R16417 VSS.n3303 VSS.n2802 80.0317
R16418 VSS.n9263 VSS.n71 80.0317
R16419 VSS.n9263 VSS.n69 80.0317
R16420 VSS.n778 VSS.n665 80.0317
R16421 VSS.n778 VSS.n667 80.0317
R16422 VSS.n8387 VSS.n7241 80.0317
R16423 VSS.n8387 VSS.n7243 80.0317
R16424 VSS.n7597 VSS.n7591 76.7447
R16425 VSS.n7740 VSS.n7347 76.7447
R16426 VSS.n8189 VSS.n8183 76.7447
R16427 VSS.n8332 VSS.n7761 76.7447
R16428 VSS.n1656 VSS.n1455 76.7447
R16429 VSS.n1591 VSS.n1590 76.7447
R16430 VSS.n2248 VSS.n2028 76.7447
R16431 VSS.n2183 VSS.n2182 76.7447
R16432 VSS.n3799 VSS.n3793 76.7447
R16433 VSS.n3943 VSS.n3372 76.7447
R16434 VSS.n4391 VSS.n4385 76.7447
R16435 VSS.n4535 VSS.n3964 76.7447
R16436 VSS.n4983 VSS.n4977 76.7447
R16437 VSS.n5127 VSS.n4556 76.7447
R16438 VSS.n5575 VSS.n5569 76.7447
R16439 VSS.n5719 VSS.n5148 76.7447
R16440 VSS.n6167 VSS.n6161 76.7447
R16441 VSS.n6311 VSS.n5740 76.7447
R16442 VSS.n6759 VSS.n6753 76.7447
R16443 VSS.n6903 VSS.n6332 76.7447
R16444 VSS.n6992 VSS.n2626 76.7447
R16445 VSS.n6927 VSS.n6926 76.7447
R16446 VSS.n3207 VSS.n3201 76.7447
R16447 VSS.n3351 VSS.n2779 76.7447
R16448 VSS.n9167 VSS.n9161 76.7447
R16449 VSS.n9311 VSS.n46 76.7447
R16450 VSS.n8993 VSS.n8773 76.7447
R16451 VSS.n8920 VSS.n8902 76.7447
R16452 VSS.n811 VSS.n618 76.7447
R16453 VSS.n9333 VSS.n30 76.7447
R16454 VSS.n8422 VSS.n7189 76.1251
R16455 VSS.n7322 VSS.n7316 76.1251
R16456 VSS.t86 VSS.n7960 75.1106
R16457 VSS.n7121 VSS.n7119 74.5791
R16458 VSS.n7149 VSS.n7117 74.5791
R16459 VSS.n7153 VSS.n7112 74.5791
R16460 VSS.n7157 VSS.n7112 74.5791
R16461 VSS.n7170 VSS.n7108 74.5791
R16462 VSS.n7186 VSS.n7101 74.5791
R16463 VSS.n7974 VSS.n7961 74.5791
R16464 VSS.n8009 VSS.n7958 74.5791
R16465 VSS.n8005 VSS.n7938 74.5791
R16466 VSS.n8036 VSS.n7938 74.5791
R16467 VSS.n8042 VSS.n7936 74.5791
R16468 VSS.n8068 VSS.n7905 74.5791
R16469 VSS.n1071 VSS.n1069 74.5791
R16470 VSS.n1097 VSS.n1067 74.5791
R16471 VSS.n1101 VSS.n1062 74.5791
R16472 VSS.n1105 VSS.n1062 74.5791
R16473 VSS.n1118 VSS.n1057 74.5791
R16474 VSS.n1135 VSS.n1050 74.5791
R16475 VSS.n890 VSS.n888 74.5791
R16476 VSS.n916 VSS.n886 74.5791
R16477 VSS.n920 VSS.n881 74.5791
R16478 VSS.n924 VSS.n881 74.5791
R16479 VSS.n937 VSS.n876 74.5791
R16480 VSS.n954 VSS.n869 74.5791
R16481 VSS.n7506 VSS.n7468 74.5791
R16482 VSS.n7510 VSS.n7454 74.5791
R16483 VSS.n7533 VSS.n7451 74.5791
R16484 VSS.n7533 VSS.n7452 74.5791
R16485 VSS.n7559 VSS.n7431 74.5791
R16486 VSS.n7581 VSS.n7418 74.5791
R16487 VSS.n8098 VSS.n7882 74.5791
R16488 VSS.n8102 VSS.n7868 74.5791
R16489 VSS.n8125 VSS.n7865 74.5791
R16490 VSS.n8125 VSS.n7866 74.5791
R16491 VSS.n8151 VSS.n7845 74.5791
R16492 VSS.n8173 VSS.n7832 74.5791
R16493 VSS.n8700 VSS.n8698 74.5791
R16494 VSS.n8728 VSS.n8696 74.5791
R16495 VSS.n8732 VSS.n8691 74.5791
R16496 VSS.n8736 VSS.n8691 74.5791
R16497 VSS.n8749 VSS.n8687 74.5791
R16498 VSS.n8765 VSS.n8680 74.5791
R16499 VSS.n271 VSS.n258 74.5791
R16500 VSS.n8570 VSS.n255 74.5791
R16501 VSS.n8566 VSS.n235 74.5791
R16502 VSS.n8597 VSS.n235 74.5791
R16503 VSS.n8603 VSS.n233 74.5791
R16504 VSS.n8629 VSS.n202 74.5791
R16505 VSS.n1217 VSS.n1204 74.5791
R16506 VSS.n1252 VSS.n1201 74.5791
R16507 VSS.n1248 VSS.n1181 74.5791
R16508 VSS.n1279 VSS.n1181 74.5791
R16509 VSS.n1285 VSS.n1179 74.5791
R16510 VSS.n1311 VSS.n1148 74.5791
R16511 VSS.n1382 VSS.n1380 74.5791
R16512 VSS.n1410 VSS.n1378 74.5791
R16513 VSS.n1414 VSS.n1373 74.5791
R16514 VSS.n1418 VSS.n1373 74.5791
R16515 VSS.n1431 VSS.n1369 74.5791
R16516 VSS.n1447 VSS.n1362 74.5791
R16517 VSS.n1790 VSS.n1777 74.5791
R16518 VSS.n1825 VSS.n1774 74.5791
R16519 VSS.n1821 VSS.n1754 74.5791
R16520 VSS.n1852 VSS.n1754 74.5791
R16521 VSS.n1858 VSS.n1752 74.5791
R16522 VSS.n1884 VSS.n1721 74.5791
R16523 VSS.n1955 VSS.n1953 74.5791
R16524 VSS.n1983 VSS.n1951 74.5791
R16525 VSS.n1987 VSS.n1946 74.5791
R16526 VSS.n1991 VSS.n1946 74.5791
R16527 VSS.n2004 VSS.n1942 74.5791
R16528 VSS.n2020 VSS.n1935 74.5791
R16529 VSS.n3584 VSS.n3571 74.5791
R16530 VSS.n3619 VSS.n3568 74.5791
R16531 VSS.n3615 VSS.n3548 74.5791
R16532 VSS.n3646 VSS.n3548 74.5791
R16533 VSS.n3652 VSS.n3546 74.5791
R16534 VSS.n3678 VSS.n3515 74.5791
R16535 VSS.n3708 VSS.n3492 74.5791
R16536 VSS.n3712 VSS.n3478 74.5791
R16537 VSS.n3735 VSS.n3475 74.5791
R16538 VSS.n3735 VSS.n3476 74.5791
R16539 VSS.n3761 VSS.n3455 74.5791
R16540 VSS.n3783 VSS.n3442 74.5791
R16541 VSS.n4176 VSS.n4163 74.5791
R16542 VSS.n4211 VSS.n4160 74.5791
R16543 VSS.n4207 VSS.n4140 74.5791
R16544 VSS.n4238 VSS.n4140 74.5791
R16545 VSS.n4244 VSS.n4138 74.5791
R16546 VSS.n4270 VSS.n4107 74.5791
R16547 VSS.n4300 VSS.n4084 74.5791
R16548 VSS.n4304 VSS.n4070 74.5791
R16549 VSS.n4327 VSS.n4067 74.5791
R16550 VSS.n4327 VSS.n4068 74.5791
R16551 VSS.n4353 VSS.n4047 74.5791
R16552 VSS.n4375 VSS.n4034 74.5791
R16553 VSS.n4768 VSS.n4755 74.5791
R16554 VSS.n4803 VSS.n4752 74.5791
R16555 VSS.n4799 VSS.n4732 74.5791
R16556 VSS.n4830 VSS.n4732 74.5791
R16557 VSS.n4836 VSS.n4730 74.5791
R16558 VSS.n4862 VSS.n4699 74.5791
R16559 VSS.n4892 VSS.n4676 74.5791
R16560 VSS.n4896 VSS.n4662 74.5791
R16561 VSS.n4919 VSS.n4659 74.5791
R16562 VSS.n4919 VSS.n4660 74.5791
R16563 VSS.n4945 VSS.n4639 74.5791
R16564 VSS.n4967 VSS.n4626 74.5791
R16565 VSS.n5360 VSS.n5347 74.5791
R16566 VSS.n5395 VSS.n5344 74.5791
R16567 VSS.n5391 VSS.n5324 74.5791
R16568 VSS.n5422 VSS.n5324 74.5791
R16569 VSS.n5428 VSS.n5322 74.5791
R16570 VSS.n5454 VSS.n5291 74.5791
R16571 VSS.n5484 VSS.n5268 74.5791
R16572 VSS.n5488 VSS.n5254 74.5791
R16573 VSS.n5511 VSS.n5251 74.5791
R16574 VSS.n5511 VSS.n5252 74.5791
R16575 VSS.n5537 VSS.n5231 74.5791
R16576 VSS.n5559 VSS.n5218 74.5791
R16577 VSS.n5952 VSS.n5939 74.5791
R16578 VSS.n5987 VSS.n5936 74.5791
R16579 VSS.n5983 VSS.n5916 74.5791
R16580 VSS.n6014 VSS.n5916 74.5791
R16581 VSS.n6020 VSS.n5914 74.5791
R16582 VSS.n6046 VSS.n5883 74.5791
R16583 VSS.n6076 VSS.n5860 74.5791
R16584 VSS.n6080 VSS.n5846 74.5791
R16585 VSS.n6103 VSS.n5843 74.5791
R16586 VSS.n6103 VSS.n5844 74.5791
R16587 VSS.n6129 VSS.n5823 74.5791
R16588 VSS.n6151 VSS.n5810 74.5791
R16589 VSS.n6544 VSS.n6531 74.5791
R16590 VSS.n6579 VSS.n6528 74.5791
R16591 VSS.n6575 VSS.n6508 74.5791
R16592 VSS.n6606 VSS.n6508 74.5791
R16593 VSS.n6612 VSS.n6506 74.5791
R16594 VSS.n6638 VSS.n6475 74.5791
R16595 VSS.n6668 VSS.n6452 74.5791
R16596 VSS.n6672 VSS.n6438 74.5791
R16597 VSS.n6695 VSS.n6435 74.5791
R16598 VSS.n6695 VSS.n6436 74.5791
R16599 VSS.n6721 VSS.n6415 74.5791
R16600 VSS.n6743 VSS.n6402 74.5791
R16601 VSS.n2388 VSS.n2375 74.5791
R16602 VSS.n2423 VSS.n2372 74.5791
R16603 VSS.n2419 VSS.n2352 74.5791
R16604 VSS.n2450 VSS.n2352 74.5791
R16605 VSS.n2456 VSS.n2350 74.5791
R16606 VSS.n2482 VSS.n2319 74.5791
R16607 VSS.n2553 VSS.n2551 74.5791
R16608 VSS.n2581 VSS.n2549 74.5791
R16609 VSS.n2585 VSS.n2544 74.5791
R16610 VSS.n2589 VSS.n2544 74.5791
R16611 VSS.n2602 VSS.n2540 74.5791
R16612 VSS.n2618 VSS.n2533 74.5791
R16613 VSS.n3011 VSS.n2974 74.5791
R16614 VSS.n3015 VSS.n2962 74.5791
R16615 VSS.n3038 VSS.n2959 74.5791
R16616 VSS.n3038 VSS.n2960 74.5791
R16617 VSS.n3064 VSS.n2937 74.5791
R16618 VSS.n3087 VSS.n2924 74.5791
R16619 VSS.n3116 VSS.n2899 74.5791
R16620 VSS.n3120 VSS.n2885 74.5791
R16621 VSS.n3143 VSS.n2882 74.5791
R16622 VSS.n3143 VSS.n2883 74.5791
R16623 VSS.n3169 VSS.n2862 74.5791
R16624 VSS.n3191 VSS.n2849 74.5791
R16625 VSS.n342 VSS.n328 74.5791
R16626 VSS.n356 VSS.n325 74.5791
R16627 VSS.n360 VSS.n321 74.5791
R16628 VSS.n365 VSS.n321 74.5791
R16629 VSS.n369 VSS.n315 74.5791
R16630 VSS.n386 VSS.n313 74.5791
R16631 VSS.n9076 VSS.n166 74.5791
R16632 VSS.n9080 VSS.n152 74.5791
R16633 VSS.n9103 VSS.n149 74.5791
R16634 VSS.n9103 VSS.n150 74.5791
R16635 VSS.n9129 VSS.n129 74.5791
R16636 VSS.n9151 VSS.n116 74.5791
R16637 VSS.n547 VSS.n540 74.5791
R16638 VSS.n573 VSS.n538 74.5791
R16639 VSS.n577 VSS.n533 74.5791
R16640 VSS.n581 VSS.n533 74.5791
R16641 VSS.n594 VSS.n529 74.5791
R16642 VSS.n610 VSS.n522 74.5791
R16643 VSS.n7482 VSS.n7481 68.3621
R16644 VSS.n7583 VSS.n7582 68.3621
R16645 VSS.n7896 VSS.n7895 68.3621
R16646 VSS.n8175 VSS.n8174 68.3621
R16647 VSS.n8538 VSS.n8537 68.3621
R16648 VSS.n8632 VSS.n8631 68.3621
R16649 VSS.n1381 VSS.n1139 68.3621
R16650 VSS.n1449 VSS.n1448 68.3621
R16651 VSS.n1220 VSS.n1219 68.3621
R16652 VSS.n1314 VSS.n1313 68.3621
R16653 VSS.n1954 VSS.n1712 68.3621
R16654 VSS.n2022 VSS.n2021 68.3621
R16655 VSS.n1793 VSS.n1792 68.3621
R16656 VSS.n1887 VSS.n1886 68.3621
R16657 VSS.n3506 VSS.n3505 68.3621
R16658 VSS.n3785 VSS.n3784 68.3621
R16659 VSS.n3587 VSS.n3586 68.3621
R16660 VSS.n3681 VSS.n3680 68.3621
R16661 VSS.n4098 VSS.n4097 68.3621
R16662 VSS.n4377 VSS.n4376 68.3621
R16663 VSS.n4179 VSS.n4178 68.3621
R16664 VSS.n4273 VSS.n4272 68.3621
R16665 VSS.n4690 VSS.n4689 68.3621
R16666 VSS.n4969 VSS.n4968 68.3621
R16667 VSS.n4771 VSS.n4770 68.3621
R16668 VSS.n4865 VSS.n4864 68.3621
R16669 VSS.n5282 VSS.n5281 68.3621
R16670 VSS.n5561 VSS.n5560 68.3621
R16671 VSS.n5363 VSS.n5362 68.3621
R16672 VSS.n5457 VSS.n5456 68.3621
R16673 VSS.n5874 VSS.n5873 68.3621
R16674 VSS.n6153 VSS.n6152 68.3621
R16675 VSS.n5955 VSS.n5954 68.3621
R16676 VSS.n6049 VSS.n6048 68.3621
R16677 VSS.n6466 VSS.n6465 68.3621
R16678 VSS.n6745 VSS.n6744 68.3621
R16679 VSS.n6547 VSS.n6546 68.3621
R16680 VSS.n6641 VSS.n6640 68.3621
R16681 VSS.n2552 VSS.n2310 68.3621
R16682 VSS.n2620 VSS.n2619 68.3621
R16683 VSS.n2391 VSS.n2390 68.3621
R16684 VSS.n2485 VSS.n2484 68.3621
R16685 VSS.n2913 VSS.n2912 68.3621
R16686 VSS.n3193 VSS.n3192 68.3621
R16687 VSS.n2988 VSS.n2987 68.3621
R16688 VSS.n3089 VSS.n3088 68.3621
R16689 VSS.n185 VSS.n184 68.3621
R16690 VSS.n9153 VSS.n9152 68.3621
R16691 VSS.n343 VSS.n272 68.3621
R16692 VSS.n385 VSS.n183 68.3621
R16693 VSS.n8699 VSS.n193 68.3621
R16694 VSS.n8767 VSS.n8766 68.3621
R16695 VSS.n546 VSS.n545 68.3621
R16696 VSS.n612 VSS.n611 68.3621
R16697 VSS.n889 VSS.n438 68.3621
R16698 VSS.n956 VSS.n955 68.3621
R16699 VSS.n1070 VSS.n1005 68.3621
R16700 VSS.n1137 VSS.n1136 68.3621
R16701 VSS.n7599 VSS.n7584 63.954
R16702 VSS.n7743 VSS.n7742 63.954
R16703 VSS.n8191 VSS.n8176 63.954
R16704 VSS.n8335 VSS.n8334 63.954
R16705 VSS.n1658 VSS.n1450 63.954
R16706 VSS.n9343 VSS.n9342 63.954
R16707 VSS.n2250 VSS.n2023 63.954
R16708 VSS.n2156 VSS.n2150 63.954
R16709 VSS.n3801 VSS.n3786 63.954
R16710 VSS.n3946 VSS.n3945 63.954
R16711 VSS.n4393 VSS.n4378 63.954
R16712 VSS.n4538 VSS.n4537 63.954
R16713 VSS.n4985 VSS.n4970 63.954
R16714 VSS.n5130 VSS.n5129 63.954
R16715 VSS.n5577 VSS.n5562 63.954
R16716 VSS.n5722 VSS.n5721 63.954
R16717 VSS.n6169 VSS.n6154 63.954
R16718 VSS.n6314 VSS.n6313 63.954
R16719 VSS.n6761 VSS.n6746 63.954
R16720 VSS.n6906 VSS.n6905 63.954
R16721 VSS.n6994 VSS.n2621 63.954
R16722 VSS.n2754 VSS.n2748 63.954
R16723 VSS.n3209 VSS.n3194 63.954
R16724 VSS.n3354 VSS.n3353 63.954
R16725 VSS.n9169 VSS.n9154 63.954
R16726 VSS.n9314 VSS.n9313 63.954
R16727 VSS.n8995 VSS.n8768 63.954
R16728 VSS.n8923 VSS.n8922 63.954
R16729 VSS.n813 VSS.n613 63.954
R16730 VSS.n9335 VSS.n25 63.954
R16731 VSS.n9340 VSS.t29 55.9858
R16732 VSS.n7976 VSS.t86 53.3045
R16733 VSS.n8426 VSS.n7189 53.2877
R16734 VSS.n7322 VSS.n16 53.2877
R16735 VSS.n478 VSS.t132 46.866
R16736 VSS.n1045 VSS.t181 46.866
R16737 VSS.n7903 VSS.t213 46.866
R16738 VSS.n200 VSS.t158 46.866
R16739 VSS.n1146 VSS.t89 46.866
R16740 VSS.n1719 VSS.t137 46.866
R16741 VSS.n3513 VSS.t266 46.866
R16742 VSS.n4105 VSS.t13 46.866
R16743 VSS.n4697 VSS.t183 46.866
R16744 VSS.n5289 VSS.t11 46.866
R16745 VSS.n5881 VSS.t317 46.866
R16746 VSS.n6473 VSS.t155 46.866
R16747 VSS.n2317 VSS.t44 46.866
R16748 VSS.n2920 VSS.t46 46.866
R16749 VSS.n180 VSS.t271 46.866
R16750 VSS.n7096 VSS.t286 46.863
R16751 VSS.n7414 VSS.t72 46.863
R16752 VSS.n7828 VSS.t126 46.863
R16753 VSS.n8675 VSS.t263 46.863
R16754 VSS.n1357 VSS.t140 46.863
R16755 VSS.n1930 VSS.t173 46.863
R16756 VSS.n3438 VSS.t249 46.863
R16757 VSS.n4030 VSS.t171 46.863
R16758 VSS.n4622 VSS.t128 46.863
R16759 VSS.n5214 VSS.t97 46.863
R16760 VSS.n5806 VSS.t189 46.863
R16761 VSS.n6398 VSS.t237 46.863
R16762 VSS.n2528 VSS.t152 46.863
R16763 VSS.n2845 VSS.t25 46.863
R16764 VSS.n112 VSS.t219 46.863
R16765 VSS.n517 VSS.t28 46.863
R16766 VSS.n7067 VSS.t161 46.8459
R16767 VSS.n7464 VSS.t289 46.8459
R16768 VSS.n7878 VSS.t222 46.8459
R16769 VSS.n8646 VSS.t147 46.8459
R16770 VSS.n1328 VSS.t165 46.8459
R16771 VSS.n1901 VSS.t22 46.8459
R16772 VSS.n3488 VSS.t200 46.8459
R16773 VSS.n4080 VSS.t240 46.8459
R16774 VSS.n4672 VSS.t168 46.8459
R16775 VSS.n5264 VSS.t210 46.8459
R16776 VSS.n5856 VSS.t187 46.8459
R16777 VSS.n6448 VSS.t299 46.8459
R16778 VSS.n2499 VSS.t203 46.8459
R16779 VSS.n2895 VSS.t60 46.8459
R16780 VSS.n162 VSS.t111 46.8459
R16781 VSS.n488 VSS.t256 46.8459
R16782 VSS.n448 VSS.t269 46.8455
R16783 VSS.n1015 VSS.t20 46.8455
R16784 VSS.n7965 VSS.t87 46.8455
R16785 VSS.n262 VSS.t9 46.8455
R16786 VSS.n1208 VSS.t53 46.8455
R16787 VSS.n1781 VSS.t69 46.8455
R16788 VSS.n3575 VSS.t62 46.8455
R16789 VSS.n4167 VSS.t150 46.8455
R16790 VSS.n4759 VSS.t66 46.8455
R16791 VSS.n5351 VSS.t83 46.8455
R16792 VSS.n5943 VSS.t296 46.8455
R16793 VSS.n6535 VSS.t193 46.8455
R16794 VSS.n2379 VSS.t234 46.8455
R16795 VSS.n2971 VSS.t217 46.8455
R16796 VSS.n282 VSS.t310 46.8455
R16797 VSS.n7729 VSS.t314 46.8085
R16798 VSS.n8321 VSS.t48 46.8085
R16799 VSS.n8889 VSS.t143 46.8085
R16800 VSS.n1558 VSS.t93 46.8085
R16801 VSS.n2166 VSS.t245 46.8085
R16802 VSS.n3932 VSS.t16 46.8085
R16803 VSS.n4524 VSS.t121 46.8085
R16804 VSS.n5116 VSS.t273 46.8085
R16805 VSS.n5708 VSS.t107 46.8085
R16806 VSS.n6300 VSS.t282 46.8085
R16807 VSS.n6892 VSS.t206 46.8085
R16808 VSS.n2764 VSS.t56 46.8085
R16809 VSS.n3340 VSS.t5 46.8085
R16810 VSS.n9300 VSS.t291 46.8085
R16811 VSS.n720 VSS.t103 46.8085
R16812 VSS.n7332 VSS.t302 46.8085
R16813 VSS.n7390 VSS.t79 46.808
R16814 VSS.n7804 VSS.t226 46.808
R16815 VSS.n8970 VSS.t35 46.808
R16816 VSS.n1500 VSS.t114 46.808
R16817 VSS.n2073 VSS.t177 46.808
R16818 VSS.n3414 VSS.t252 46.808
R16819 VSS.n4006 VSS.t231 46.808
R16820 VSS.n4598 VSS.t118 46.808
R16821 VSS.n5190 VSS.t306 46.808
R16822 VSS.n5782 VSS.t278 46.808
R16823 VSS.n6374 VSS.t99 46.808
R16824 VSS.n2671 VSS.t196 46.808
R16825 VSS.n2821 VSS.t32 46.808
R16826 VSS.n88 VSS.t40 46.808
R16827 VSS.n663 VSS.t258 46.808
R16828 VSS.n7239 VSS.t76 46.808
R16829 VSS.n8474 VSS.n7057 44.8985
R16830 VSS.n8429 VSS.n7188 44.8985
R16831 VSS.n7603 VSS.n7584 44.7679
R16832 VSS.n7742 VSS.n17 44.7679
R16833 VSS.n8195 VSS.n8176 44.7679
R16834 VSS.n8334 VSS.n15 44.7679
R16835 VSS.n1662 VSS.n1450 44.7679
R16836 VSS.n9342 VSS.n9341 44.7679
R16837 VSS.n2254 VSS.n2023 44.7679
R16838 VSS.n2156 VSS.n18 44.7679
R16839 VSS.n3805 VSS.n3786 44.7679
R16840 VSS.n3945 VSS.n14 44.7679
R16841 VSS.n4397 VSS.n4378 44.7679
R16842 VSS.n4537 VSS.n19 44.7679
R16843 VSS.n4989 VSS.n4970 44.7679
R16844 VSS.n5129 VSS.n13 44.7679
R16845 VSS.n5581 VSS.n5562 44.7679
R16846 VSS.n5721 VSS.n20 44.7679
R16847 VSS.n6173 VSS.n6154 44.7679
R16848 VSS.n6313 VSS.n12 44.7679
R16849 VSS.n6765 VSS.n6746 44.7679
R16850 VSS.n6905 VSS.n21 44.7679
R16851 VSS.n6998 VSS.n2621 44.7679
R16852 VSS.n2754 VSS.n11 44.7679
R16853 VSS.n3213 VSS.n3194 44.7679
R16854 VSS.n3353 VSS.n22 44.7679
R16855 VSS.n9173 VSS.n9154 44.7679
R16856 VSS.n9313 VSS.n23 44.7679
R16857 VSS.n8999 VSS.n8768 44.7679
R16858 VSS.n8922 VSS.n10 44.7679
R16859 VSS.n817 VSS.n613 44.7679
R16860 VSS.n9339 VSS.n25 44.7679
R16861 VSS.n8421 VSS.n8420 38.0628
R16862 VSS.n8354 VSS.n8353 38.0628
R16863 VSS.n7482 VSS.n7480 37.2886
R16864 VSS.n7606 VSS.n7583 37.2886
R16865 VSS.n7896 VSS.n7894 37.2886
R16866 VSS.n8198 VSS.n8175 37.2886
R16867 VSS.n8538 VSS.n8536 37.2886
R16868 VSS.n8632 VSS.n192 37.2886
R16869 VSS.n1710 VSS.n1139 37.2886
R16870 VSS.n1665 VSS.n1449 37.2886
R16871 VSS.n1220 VSS.n1218 37.2886
R16872 VSS.n1314 VSS.n1138 37.2886
R16873 VSS.n2302 VSS.n1712 37.2886
R16874 VSS.n2257 VSS.n2022 37.2886
R16875 VSS.n1793 VSS.n1791 37.2886
R16876 VSS.n1887 VSS.n1711 37.2886
R16877 VSS.n3506 VSS.n3504 37.2886
R16878 VSS.n3808 VSS.n3785 37.2886
R16879 VSS.n3587 VSS.n3585 37.2886
R16880 VSS.n3681 VSS.n2303 37.2886
R16881 VSS.n4098 VSS.n4096 37.2886
R16882 VSS.n4400 VSS.n4377 37.2886
R16883 VSS.n4179 VSS.n4177 37.2886
R16884 VSS.n4273 VSS.n2304 37.2886
R16885 VSS.n4690 VSS.n4688 37.2886
R16886 VSS.n4992 VSS.n4969 37.2886
R16887 VSS.n4771 VSS.n4769 37.2886
R16888 VSS.n4865 VSS.n2305 37.2886
R16889 VSS.n5282 VSS.n5280 37.2886
R16890 VSS.n5584 VSS.n5561 37.2886
R16891 VSS.n5363 VSS.n5361 37.2886
R16892 VSS.n5457 VSS.n2306 37.2886
R16893 VSS.n5874 VSS.n5872 37.2886
R16894 VSS.n6176 VSS.n6153 37.2886
R16895 VSS.n5955 VSS.n5953 37.2886
R16896 VSS.n6049 VSS.n2307 37.2886
R16897 VSS.n6466 VSS.n6464 37.2886
R16898 VSS.n6768 VSS.n6745 37.2886
R16899 VSS.n6547 VSS.n6545 37.2886
R16900 VSS.n6641 VSS.n2308 37.2886
R16901 VSS.n7046 VSS.n2310 37.2886
R16902 VSS.n7001 VSS.n2620 37.2886
R16903 VSS.n2391 VSS.n2389 37.2886
R16904 VSS.n2485 VSS.n2309 37.2886
R16905 VSS.n2913 VSS.n2911 37.2886
R16906 VSS.n3216 VSS.n3193 37.2886
R16907 VSS.n2988 VSS.n2986 37.2886
R16908 VSS.n3090 VSS.n3089 37.2886
R16909 VSS.n190 VSS.n185 37.2886
R16910 VSS.n9176 VSS.n9153 37.2886
R16911 VSS.n437 VSS.n272 37.2886
R16912 VSS.n9050 VSS.n183 37.2886
R16913 VSS.n9047 VSS.n193 37.2886
R16914 VSS.n9002 VSS.n8767 37.2886
R16915 VSS.n545 VSS.n544 37.2886
R16916 VSS.n820 VSS.n612 37.2886
R16917 VSS.n1002 VSS.n438 37.2886
R16918 VSS.n957 VSS.n956 37.2886
R16919 VSS.n8523 VSS.n1005 37.2886
R16920 VSS.n8478 VSS.n1137 37.2886
R16921 VSS.n8007 VSS.n8006 36.3441
R16922 VSS.n8038 VSS.n8037 36.3441
R16923 VSS.t29 VSS.t1 34.4875
R16924 VSS.n8428 VSS.n8427 33.5883
R16925 VSS.t0 VSS.t2 32.6959
R16926 VSS.t1 VSS.t0 32.2481
R16927 VSS.n7598 VSS.n7597 31.9772
R16928 VSS.n7741 VSS.n7740 31.9772
R16929 VSS.n8190 VSS.n8189 31.9772
R16930 VSS.n8333 VSS.n8332 31.9772
R16931 VSS.n1657 VSS.n1656 31.9772
R16932 VSS.n1590 VSS.n9 31.9772
R16933 VSS.n2249 VSS.n2248 31.9772
R16934 VSS.n2182 VSS.n2181 31.9772
R16935 VSS.n3800 VSS.n3799 31.9772
R16936 VSS.n3944 VSS.n3943 31.9772
R16937 VSS.n4392 VSS.n4391 31.9772
R16938 VSS.n4536 VSS.n4535 31.9772
R16939 VSS.n4984 VSS.n4983 31.9772
R16940 VSS.n5128 VSS.n5127 31.9772
R16941 VSS.n5576 VSS.n5575 31.9772
R16942 VSS.n5720 VSS.n5719 31.9772
R16943 VSS.n6168 VSS.n6167 31.9772
R16944 VSS.n6312 VSS.n6311 31.9772
R16945 VSS.n6760 VSS.n6759 31.9772
R16946 VSS.n6904 VSS.n6903 31.9772
R16947 VSS.n6993 VSS.n6992 31.9772
R16948 VSS.n6926 VSS.n6925 31.9772
R16949 VSS.n3208 VSS.n3207 31.9772
R16950 VSS.n3352 VSS.n3351 31.9772
R16951 VSS.n9168 VSS.n9167 31.9772
R16952 VSS.n9312 VSS.n9311 31.9772
R16953 VSS.n8994 VSS.n8993 31.9772
R16954 VSS.n8921 VSS.n8920 31.9772
R16955 VSS.n812 VSS.n811 31.9772
R16956 VSS.n9334 VSS.n9333 31.9772
R16957 VSS.n8004 VSS.n8003 31.4983
R16958 VSS.n8040 VSS.n8039 31.4983
R16959 VSS.n7146 VSS.n7118 29.9325
R16960 VSS.t285 VSS.n7100 29.9325
R16961 VSS.n7977 VSS.n7976 26.6525
R16962 VSS.n8071 VSS.n8070 26.6525
R16963 VSS.n7508 VSS.n7507 24.8593
R16964 VSS.t71 VSS.n7417 24.8593
R16965 VSS.n8100 VSS.n8099 24.8593
R16966 VSS.t125 VSS.n7831 24.8593
R16967 VSS.n8564 VSS.n257 24.8593
R16968 VSS.n1407 VSS.n1379 24.8593
R16969 VSS.t139 VSS.n1361 24.8593
R16970 VSS.n1246 VSS.n1203 24.8593
R16971 VSS.n1980 VSS.n1952 24.8593
R16972 VSS.t172 VSS.n1934 24.8593
R16973 VSS.n1819 VSS.n1776 24.8593
R16974 VSS.n3710 VSS.n3709 24.8593
R16975 VSS.t248 VSS.n3441 24.8593
R16976 VSS.n3613 VSS.n3570 24.8593
R16977 VSS.n4302 VSS.n4301 24.8593
R16978 VSS.t170 VSS.n4033 24.8593
R16979 VSS.n4205 VSS.n4162 24.8593
R16980 VSS.n4894 VSS.n4893 24.8593
R16981 VSS.t127 VSS.n4625 24.8593
R16982 VSS.n4797 VSS.n4754 24.8593
R16983 VSS.n5486 VSS.n5485 24.8593
R16984 VSS.t96 VSS.n5217 24.8593
R16985 VSS.n5389 VSS.n5346 24.8593
R16986 VSS.n6078 VSS.n6077 24.8593
R16987 VSS.t188 VSS.n5809 24.8593
R16988 VSS.n5981 VSS.n5938 24.8593
R16989 VSS.n6670 VSS.n6669 24.8593
R16990 VSS.t236 VSS.n6401 24.8593
R16991 VSS.n6573 VSS.n6530 24.8593
R16992 VSS.n2578 VSS.n2550 24.8593
R16993 VSS.t151 VSS.n2532 24.8593
R16994 VSS.n2417 VSS.n2374 24.8593
R16995 VSS.n3118 VSS.n3117 24.8593
R16996 VSS.t24 VSS.n2848 24.8593
R16997 VSS.n3013 VSS.n3012 24.8593
R16998 VSS.n9078 VSS.n9077 24.8593
R16999 VSS.t218 VSS.n115 24.8593
R17000 VSS.n345 VSS.n344 24.8593
R17001 VSS.n8725 VSS.n8697 24.8593
R17002 VSS.t262 VSS.n8679 24.8593
R17003 VSS.n570 VSS.n539 24.8593
R17004 VSS.t27 VSS.n521 24.8593
R17005 VSS.n913 VSS.n887 24.8593
R17006 VSS.n1094 VSS.n1068 24.8593
R17007 VSS.n7393 VSS.n7373 24.6255
R17008 VSS.n7697 VSS.n7371 24.6255
R17009 VSS.n7807 VSS.n7787 24.6255
R17010 VSS.n8289 VSS.n7785 24.6255
R17011 VSS.n8844 VSS.n8822 24.6255
R17012 VSS.n8956 VSS.n8823 24.6255
R17013 VSS.n1627 VSS.n1502 24.6255
R17014 VSS.n1580 VSS.n1504 24.6255
R17015 VSS.n2219 VSS.n2075 24.6255
R17016 VSS.n2140 VSS.n2077 24.6255
R17017 VSS.n3417 VSS.n3397 24.6255
R17018 VSS.n3899 VSS.n3395 24.6255
R17019 VSS.n4009 VSS.n3989 24.6255
R17020 VSS.n4491 VSS.n3987 24.6255
R17021 VSS.n4601 VSS.n4581 24.6255
R17022 VSS.n5083 VSS.n4579 24.6255
R17023 VSS.n5193 VSS.n5173 24.6255
R17024 VSS.n5675 VSS.n5171 24.6255
R17025 VSS.n5785 VSS.n5765 24.6255
R17026 VSS.n6267 VSS.n5763 24.6255
R17027 VSS.n6377 VSS.n6357 24.6255
R17028 VSS.n6859 VSS.n6355 24.6255
R17029 VSS.n6963 VSS.n2673 24.6255
R17030 VSS.n2738 VSS.n2675 24.6255
R17031 VSS.n2824 VSS.n2804 24.6255
R17032 VSS.n3307 VSS.n2802 24.6255
R17033 VSS.n91 VSS.n71 24.6255
R17034 VSS.n9267 VSS.n69 24.6255
R17035 VSS.n782 VSS.n665 24.6255
R17036 VSS.n740 VSS.n667 24.6255
R17037 VSS.n8391 VSS.n7241 24.6255
R17038 VSS.n7306 VSS.n7243 24.6255
R17039 VSS.n8406 VSS.n8405 22.8379
R17040 VSS.n7315 VSS.t301 22.8379
R17041 VSS.n7642 VSS.n7392 21.5474
R17042 VSS.n7714 VSS.n7359 21.5474
R17043 VSS.n8234 VSS.n7806 21.5474
R17044 VSS.n8306 VSS.n7773 21.5474
R17045 VSS.n8835 VSS.n8825 21.5474
R17046 VSS.n8912 VSS.n8903 21.5474
R17047 VSS.n1639 VSS.n1484 21.5474
R17048 VSS.n1588 VSS.n1584 21.5474
R17049 VSS.n2231 VSS.n2057 21.5474
R17050 VSS.n2148 VSS.n2144 21.5474
R17051 VSS.n3844 VSS.n3416 21.5474
R17052 VSS.n3916 VSS.n3383 21.5474
R17053 VSS.n4436 VSS.n4008 21.5474
R17054 VSS.n4508 VSS.n3975 21.5474
R17055 VSS.n5028 VSS.n4600 21.5474
R17056 VSS.n5100 VSS.n4567 21.5474
R17057 VSS.n5620 VSS.n5192 21.5474
R17058 VSS.n5692 VSS.n5159 21.5474
R17059 VSS.n6212 VSS.n5784 21.5474
R17060 VSS.n6284 VSS.n5751 21.5474
R17061 VSS.n6804 VSS.n6376 21.5474
R17062 VSS.n6876 VSS.n6343 21.5474
R17063 VSS.n6975 VSS.n2655 21.5474
R17064 VSS.n2746 VSS.n2742 21.5474
R17065 VSS.n3252 VSS.n2823 21.5474
R17066 VSS.n3324 VSS.n2790 21.5474
R17067 VSS.n9212 VSS.n90 21.5474
R17068 VSS.n9284 VSS.n57 21.5474
R17069 VSS.n794 VSS.n647 21.5474
R17070 VSS.n742 VSS.n728 21.5474
R17071 VSS.n8403 VSS.n7223 21.5474
R17072 VSS.n7314 VSS.n7310 21.5474
R17073 VSS.n7153 VSS.n7114 21.1076
R17074 VSS.n7157 VSS.n7110 21.1076
R17075 VSS.n8005 VSS.n7959 21.1076
R17076 VSS.n8036 VSS.n7929 21.1076
R17077 VSS.n1101 VSS.n1064 21.1076
R17078 VSS.n1105 VSS.n1059 21.1076
R17079 VSS.n920 VSS.n883 21.1076
R17080 VSS.n924 VSS.n878 21.1076
R17081 VSS.n7528 VSS.n7451 21.1076
R17082 VSS.n7452 VSS.n7433 21.1076
R17083 VSS.n8120 VSS.n7865 21.1076
R17084 VSS.n7866 VSS.n7847 21.1076
R17085 VSS.n8732 VSS.n8693 21.1076
R17086 VSS.n8736 VSS.n8689 21.1076
R17087 VSS.n8566 VSS.n256 21.1076
R17088 VSS.n8597 VSS.n226 21.1076
R17089 VSS.n1248 VSS.n1202 21.1076
R17090 VSS.n1279 VSS.n1172 21.1076
R17091 VSS.n1414 VSS.n1375 21.1076
R17092 VSS.n1418 VSS.n1371 21.1076
R17093 VSS.n1821 VSS.n1775 21.1076
R17094 VSS.n1852 VSS.n1745 21.1076
R17095 VSS.n1987 VSS.n1948 21.1076
R17096 VSS.n1991 VSS.n1944 21.1076
R17097 VSS.n3615 VSS.n3569 21.1076
R17098 VSS.n3646 VSS.n3539 21.1076
R17099 VSS.n3730 VSS.n3475 21.1076
R17100 VSS.n3476 VSS.n3457 21.1076
R17101 VSS.n4207 VSS.n4161 21.1076
R17102 VSS.n4238 VSS.n4131 21.1076
R17103 VSS.n4322 VSS.n4067 21.1076
R17104 VSS.n4068 VSS.n4049 21.1076
R17105 VSS.n4799 VSS.n4753 21.1076
R17106 VSS.n4830 VSS.n4723 21.1076
R17107 VSS.n4914 VSS.n4659 21.1076
R17108 VSS.n4660 VSS.n4641 21.1076
R17109 VSS.n5391 VSS.n5345 21.1076
R17110 VSS.n5422 VSS.n5315 21.1076
R17111 VSS.n5506 VSS.n5251 21.1076
R17112 VSS.n5252 VSS.n5233 21.1076
R17113 VSS.n5983 VSS.n5937 21.1076
R17114 VSS.n6014 VSS.n5907 21.1076
R17115 VSS.n6098 VSS.n5843 21.1076
R17116 VSS.n5844 VSS.n5825 21.1076
R17117 VSS.n6575 VSS.n6529 21.1076
R17118 VSS.n6606 VSS.n6499 21.1076
R17119 VSS.n6690 VSS.n6435 21.1076
R17120 VSS.n6436 VSS.n6417 21.1076
R17121 VSS.n2419 VSS.n2373 21.1076
R17122 VSS.n2450 VSS.n2343 21.1076
R17123 VSS.n2585 VSS.n2546 21.1076
R17124 VSS.n2589 VSS.n2542 21.1076
R17125 VSS.n3033 VSS.n2959 21.1076
R17126 VSS.n2960 VSS.n2939 21.1076
R17127 VSS.n3138 VSS.n2882 21.1076
R17128 VSS.n2883 VSS.n2864 21.1076
R17129 VSS.n360 VSS.n323 21.1076
R17130 VSS.n365 VSS.n319 21.1076
R17131 VSS.n9098 VSS.n149 21.1076
R17132 VSS.n150 VSS.n131 21.1076
R17133 VSS.n577 VSS.n535 21.1076
R17134 VSS.n581 VSS.n531 21.1076
R17135 VSS.n7643 VSS.n7394 19.1865
R17136 VSS.n7716 VSS.t313 19.1865
R17137 VSS.n8235 VSS.n7808 19.1865
R17138 VSS.n8308 VSS.t47 19.1865
R17139 VSS.n1642 VSS.n1641 19.1865
R17140 VSS.n1589 VSS.t92 19.1865
R17141 VSS.n2234 VSS.n2233 19.1865
R17142 VSS.n2149 VSS.t244 19.1865
R17143 VSS.n3845 VSS.n3418 19.1865
R17144 VSS.n3918 VSS.t15 19.1865
R17145 VSS.n4437 VSS.n4010 19.1865
R17146 VSS.n4510 VSS.t120 19.1865
R17147 VSS.n5029 VSS.n4602 19.1865
R17148 VSS.n5102 VSS.t272 19.1865
R17149 VSS.n5621 VSS.n5194 19.1865
R17150 VSS.n5694 VSS.t106 19.1865
R17151 VSS.n6213 VSS.n5786 19.1865
R17152 VSS.n6286 VSS.t281 19.1865
R17153 VSS.n6805 VSS.n6378 19.1865
R17154 VSS.n6878 VSS.t205 19.1865
R17155 VSS.n6978 VSS.n6977 19.1865
R17156 VSS.n2747 VSS.t55 19.1865
R17157 VSS.n3253 VSS.n2825 19.1865
R17158 VSS.n3326 VSS.t4 19.1865
R17159 VSS.n9213 VSS.n92 19.1865
R17160 VSS.n9286 VSS.t290 19.1865
R17161 VSS.n8833 VSS.n8832 19.1865
R17162 VSS.n8914 VSS.t142 19.1865
R17163 VSS.n797 VSS.n796 19.1865
R17164 VSS.n744 VSS.t102 19.1865
R17165 VSS.n8630 VSS.t157 18.6446
R17166 VSS.n1312 VSS.t88 18.6446
R17167 VSS.n1885 VSS.t136 18.6446
R17168 VSS.n3679 VSS.t265 18.6446
R17169 VSS.n4271 VSS.t12 18.6446
R17170 VSS.n4863 VSS.t182 18.6446
R17171 VSS.n5455 VSS.t10 18.6446
R17172 VSS.n6047 VSS.t316 18.6446
R17173 VSS.n6639 VSS.t154 18.6446
R17174 VSS.n2483 VSS.t43 18.6446
R17175 VSS.t45 VSS.n2923 18.6446
R17176 VSS.n384 VSS.t270 18.6446
R17177 VSS.t131 VSS.n868 18.6446
R17178 VSS.t180 VSS.n1049 18.6446
R17179 VSS.n7596 VSS.n7592 18.4693
R17180 VSS.n7739 VSS.n7348 18.4693
R17181 VSS.n8188 VSS.n8184 18.4693
R17182 VSS.n8331 VSS.n7762 18.4693
R17183 VSS.n8992 VSS.n8774 18.4693
R17184 VSS.n8919 VSS.n8916 18.4693
R17185 VSS.n1655 VSS.n1456 18.4693
R17186 VSS.n1592 VSS.n1569 18.4693
R17187 VSS.n2247 VSS.n2029 18.4693
R17188 VSS.n2184 VSS.n2129 18.4693
R17189 VSS.n3798 VSS.n3794 18.4693
R17190 VSS.n3942 VSS.n3373 18.4693
R17191 VSS.n4390 VSS.n4386 18.4693
R17192 VSS.n4534 VSS.n3965 18.4693
R17193 VSS.n4982 VSS.n4978 18.4693
R17194 VSS.n5126 VSS.n4557 18.4693
R17195 VSS.n5574 VSS.n5570 18.4693
R17196 VSS.n5718 VSS.n5149 18.4693
R17197 VSS.n6166 VSS.n6162 18.4693
R17198 VSS.n6310 VSS.n5741 18.4693
R17199 VSS.n6758 VSS.n6754 18.4693
R17200 VSS.n6902 VSS.n6333 18.4693
R17201 VSS.n6991 VSS.n2627 18.4693
R17202 VSS.n6928 VSS.n2727 18.4693
R17203 VSS.n3206 VSS.n3202 18.4693
R17204 VSS.n3350 VSS.n2780 18.4693
R17205 VSS.n9166 VSS.n9162 18.4693
R17206 VSS.n9310 VSS.n47 18.4693
R17207 VSS.n810 VSS.n619 18.4693
R17208 VSS.n9332 VSS.n31 18.4693
R17209 VSS.n8419 VSS.n7195 18.4693
R17210 VSS.n8356 VSS.n7295 18.4693
R17211 VSS.n7145 VSS.n7117 18.2934
R17212 VSS.n7173 VSS.n7108 18.2934
R17213 VSS.n8002 VSS.n7958 18.2934
R17214 VSS.n7936 VSS.n7906 18.2934
R17215 VSS.n1093 VSS.n1067 18.2934
R17216 VSS.n1122 VSS.n1057 18.2934
R17217 VSS.n912 VSS.n886 18.2934
R17218 VSS.n941 VSS.n876 18.2934
R17219 VSS.n7510 VSS.n7467 18.2934
R17220 VSS.n7562 VSS.n7431 18.2934
R17221 VSS.n8102 VSS.n7881 18.2934
R17222 VSS.n8154 VSS.n7845 18.2934
R17223 VSS.n8724 VSS.n8696 18.2934
R17224 VSS.n8752 VSS.n8687 18.2934
R17225 VSS.n8563 VSS.n255 18.2934
R17226 VSS.n233 VSS.n203 18.2934
R17227 VSS.n1245 VSS.n1201 18.2934
R17228 VSS.n1179 VSS.n1149 18.2934
R17229 VSS.n1406 VSS.n1378 18.2934
R17230 VSS.n1434 VSS.n1369 18.2934
R17231 VSS.n1818 VSS.n1774 18.2934
R17232 VSS.n1752 VSS.n1722 18.2934
R17233 VSS.n1979 VSS.n1951 18.2934
R17234 VSS.n2007 VSS.n1942 18.2934
R17235 VSS.n3612 VSS.n3568 18.2934
R17236 VSS.n3546 VSS.n3516 18.2934
R17237 VSS.n3712 VSS.n3491 18.2934
R17238 VSS.n3764 VSS.n3455 18.2934
R17239 VSS.n4204 VSS.n4160 18.2934
R17240 VSS.n4138 VSS.n4108 18.2934
R17241 VSS.n4304 VSS.n4083 18.2934
R17242 VSS.n4356 VSS.n4047 18.2934
R17243 VSS.n4796 VSS.n4752 18.2934
R17244 VSS.n4730 VSS.n4700 18.2934
R17245 VSS.n4896 VSS.n4675 18.2934
R17246 VSS.n4948 VSS.n4639 18.2934
R17247 VSS.n5388 VSS.n5344 18.2934
R17248 VSS.n5322 VSS.n5292 18.2934
R17249 VSS.n5488 VSS.n5267 18.2934
R17250 VSS.n5540 VSS.n5231 18.2934
R17251 VSS.n5980 VSS.n5936 18.2934
R17252 VSS.n5914 VSS.n5884 18.2934
R17253 VSS.n6080 VSS.n5859 18.2934
R17254 VSS.n6132 VSS.n5823 18.2934
R17255 VSS.n6572 VSS.n6528 18.2934
R17256 VSS.n6506 VSS.n6476 18.2934
R17257 VSS.n6672 VSS.n6451 18.2934
R17258 VSS.n6724 VSS.n6415 18.2934
R17259 VSS.n2416 VSS.n2372 18.2934
R17260 VSS.n2350 VSS.n2320 18.2934
R17261 VSS.n2577 VSS.n2549 18.2934
R17262 VSS.n2605 VSS.n2540 18.2934
R17263 VSS.n3015 VSS.n2973 18.2934
R17264 VSS.n3068 VSS.n2937 18.2934
R17265 VSS.n3120 VSS.n2898 18.2934
R17266 VSS.n3172 VSS.n2862 18.2934
R17267 VSS.n346 VSS.n325 18.2934
R17268 VSS.n382 VSS.n315 18.2934
R17269 VSS.n9080 VSS.n165 18.2934
R17270 VSS.n9132 VSS.n129 18.2934
R17271 VSS.n569 VSS.n538 18.2934
R17272 VSS.n597 VSS.n529 18.2934
R17273 VSS.n7121 VSS.n7058 15.4791
R17274 VSS.n7186 VSS.n7099 15.4791
R17275 VSS.n7978 VSS.n7974 15.4791
R17276 VSS.n8072 VSS.n7905 15.4791
R17277 VSS.n1071 VSS.n1006 15.4791
R17278 VSS.n1135 VSS.n1048 15.4791
R17279 VSS.n890 VSS.n439 15.4791
R17280 VSS.n954 VSS.n867 15.4791
R17281 VSS.n7483 VSS.n7468 15.4791
R17282 VSS.n7581 VSS.n7416 15.4791
R17283 VSS.n7897 VSS.n7882 15.4791
R17284 VSS.n8173 VSS.n7830 15.4791
R17285 VSS.n8700 VSS.n194 15.4791
R17286 VSS.n8765 VSS.n8678 15.4791
R17287 VSS.n8539 VSS.n271 15.4791
R17288 VSS.n8633 VSS.n202 15.4791
R17289 VSS.n1221 VSS.n1217 15.4791
R17290 VSS.n1315 VSS.n1148 15.4791
R17291 VSS.n1382 VSS.n1140 15.4791
R17292 VSS.n1447 VSS.n1360 15.4791
R17293 VSS.n1794 VSS.n1790 15.4791
R17294 VSS.n1888 VSS.n1721 15.4791
R17295 VSS.n1955 VSS.n1713 15.4791
R17296 VSS.n2020 VSS.n1933 15.4791
R17297 VSS.n3588 VSS.n3584 15.4791
R17298 VSS.n3682 VSS.n3515 15.4791
R17299 VSS.n3507 VSS.n3492 15.4791
R17300 VSS.n3783 VSS.n3440 15.4791
R17301 VSS.n4180 VSS.n4176 15.4791
R17302 VSS.n4274 VSS.n4107 15.4791
R17303 VSS.n4099 VSS.n4084 15.4791
R17304 VSS.n4375 VSS.n4032 15.4791
R17305 VSS.n4772 VSS.n4768 15.4791
R17306 VSS.n4866 VSS.n4699 15.4791
R17307 VSS.n4691 VSS.n4676 15.4791
R17308 VSS.n4967 VSS.n4624 15.4791
R17309 VSS.n5364 VSS.n5360 15.4791
R17310 VSS.n5458 VSS.n5291 15.4791
R17311 VSS.n5283 VSS.n5268 15.4791
R17312 VSS.n5559 VSS.n5216 15.4791
R17313 VSS.n5956 VSS.n5952 15.4791
R17314 VSS.n6050 VSS.n5883 15.4791
R17315 VSS.n5875 VSS.n5860 15.4791
R17316 VSS.n6151 VSS.n5808 15.4791
R17317 VSS.n6548 VSS.n6544 15.4791
R17318 VSS.n6642 VSS.n6475 15.4791
R17319 VSS.n6467 VSS.n6452 15.4791
R17320 VSS.n6743 VSS.n6400 15.4791
R17321 VSS.n2392 VSS.n2388 15.4791
R17322 VSS.n2486 VSS.n2319 15.4791
R17323 VSS.n2553 VSS.n2311 15.4791
R17324 VSS.n2618 VSS.n2531 15.4791
R17325 VSS.n2989 VSS.n2974 15.4791
R17326 VSS.n3087 VSS.n2922 15.4791
R17327 VSS.n2914 VSS.n2899 15.4791
R17328 VSS.n3191 VSS.n2847 15.4791
R17329 VSS.n342 VSS.n273 15.4791
R17330 VSS.n386 VSS.n182 15.4791
R17331 VSS.n188 VSS.n166 15.4791
R17332 VSS.n9151 VSS.n114 15.4791
R17333 VSS.n547 VSS.n542 15.4791
R17334 VSS.n610 VSS.n520 15.4791
R17335 VSS.n7600 VSS.n7585 15.3911
R17336 VSS.n7744 VSS.n7346 15.3911
R17337 VSS.n8192 VSS.n8177 15.3911
R17338 VSS.n8336 VSS.n7760 15.3911
R17339 VSS.n8996 VSS.n8769 15.3911
R17340 VSS.n8924 VSS.n8901 15.3911
R17341 VSS.n1659 VSS.n1451 15.3911
R17342 VSS.n9344 VSS.n8 15.3911
R17343 VSS.n2251 VSS.n2024 15.3911
R17344 VSS.n2157 VSS.n2151 15.3911
R17345 VSS.n3802 VSS.n3787 15.3911
R17346 VSS.n3947 VSS.n3371 15.3911
R17347 VSS.n4394 VSS.n4379 15.3911
R17348 VSS.n4539 VSS.n3963 15.3911
R17349 VSS.n4986 VSS.n4971 15.3911
R17350 VSS.n5131 VSS.n4555 15.3911
R17351 VSS.n5578 VSS.n5563 15.3911
R17352 VSS.n5723 VSS.n5147 15.3911
R17353 VSS.n6170 VSS.n6155 15.3911
R17354 VSS.n6315 VSS.n5739 15.3911
R17355 VSS.n6762 VSS.n6747 15.3911
R17356 VSS.n6907 VSS.n6331 15.3911
R17357 VSS.n6995 VSS.n2622 15.3911
R17358 VSS.n2755 VSS.n2749 15.3911
R17359 VSS.n3210 VSS.n3195 15.3911
R17360 VSS.n3355 VSS.n2778 15.3911
R17361 VSS.n9170 VSS.n9155 15.3911
R17362 VSS.n9315 VSS.n45 15.3911
R17363 VSS.n814 VSS.n614 15.3911
R17364 VSS.n9336 VSS.n26 15.3911
R17365 VSS.n8423 VSS.n7190 15.3911
R17366 VSS.n7323 VSS.n7317 15.3911
R17367 VSS.n7148 VSS.n7113 14.9665
R17368 VSS.n7171 VSS.n7109 14.9665
R17369 VSS.n7977 VSS.n7975 14.5379
R17370 VSS.n8071 VSS.n7056 14.5379
R17371 VSS.n7529 VSS.n7453 12.4299
R17372 VSS.n7560 VSS.n7432 12.4299
R17373 VSS.n8121 VSS.n7867 12.4299
R17374 VSS.n8152 VSS.n7846 12.4299
R17375 VSS.n8569 VSS.n8568 12.4299
R17376 VSS.n8602 VSS.n8599 12.4299
R17377 VSS.n1409 VSS.n1374 12.4299
R17378 VSS.n1432 VSS.n1370 12.4299
R17379 VSS.n1251 VSS.n1250 12.4299
R17380 VSS.n1284 VSS.n1281 12.4299
R17381 VSS.n1982 VSS.n1947 12.4299
R17382 VSS.n2005 VSS.n1943 12.4299
R17383 VSS.n1824 VSS.n1823 12.4299
R17384 VSS.n1857 VSS.n1854 12.4299
R17385 VSS.n3731 VSS.n3477 12.4299
R17386 VSS.n3762 VSS.n3456 12.4299
R17387 VSS.n3618 VSS.n3617 12.4299
R17388 VSS.n3651 VSS.n3648 12.4299
R17389 VSS.n4323 VSS.n4069 12.4299
R17390 VSS.n4354 VSS.n4048 12.4299
R17391 VSS.n4210 VSS.n4209 12.4299
R17392 VSS.n4243 VSS.n4240 12.4299
R17393 VSS.n4915 VSS.n4661 12.4299
R17394 VSS.n4946 VSS.n4640 12.4299
R17395 VSS.n4802 VSS.n4801 12.4299
R17396 VSS.n4835 VSS.n4832 12.4299
R17397 VSS.n5507 VSS.n5253 12.4299
R17398 VSS.n5538 VSS.n5232 12.4299
R17399 VSS.n5394 VSS.n5393 12.4299
R17400 VSS.n5427 VSS.n5424 12.4299
R17401 VSS.n6099 VSS.n5845 12.4299
R17402 VSS.n6130 VSS.n5824 12.4299
R17403 VSS.n5986 VSS.n5985 12.4299
R17404 VSS.n6019 VSS.n6016 12.4299
R17405 VSS.n6691 VSS.n6437 12.4299
R17406 VSS.n6722 VSS.n6416 12.4299
R17407 VSS.n6578 VSS.n6577 12.4299
R17408 VSS.n6611 VSS.n6608 12.4299
R17409 VSS.n2580 VSS.n2545 12.4299
R17410 VSS.n2603 VSS.n2541 12.4299
R17411 VSS.n2422 VSS.n2421 12.4299
R17412 VSS.n2455 VSS.n2452 12.4299
R17413 VSS.n3139 VSS.n2884 12.4299
R17414 VSS.n3170 VSS.n2863 12.4299
R17415 VSS.n3034 VSS.n2961 12.4299
R17416 VSS.n3065 VSS.n2938 12.4299
R17417 VSS.n9099 VSS.n151 12.4299
R17418 VSS.n9130 VSS.n130 12.4299
R17419 VSS.n358 VSS.n357 12.4299
R17420 VSS.n368 VSS.n367 12.4299
R17421 VSS.n8727 VSS.n8692 12.4299
R17422 VSS.n8750 VSS.n8688 12.4299
R17423 VSS.n572 VSS.n534 12.4299
R17424 VSS.n595 VSS.n530 12.4299
R17425 VSS.n915 VSS.n882 12.4299
R17426 VSS.n938 VSS.n877 12.4299
R17427 VSS.n1096 VSS.n1063 12.4299
R17428 VSS.n1119 VSS.n1058 12.4299
R17429 VSS.n8003 VSS.n7960 9.69213
R17430 VSS.n8473 VSS.n8472 9.38145
R17431 VSS.n8522 VSS.n8521 9.38145
R17432 VSS.n7485 VSS.n7478 9.38145
R17433 VSS.n7980 VSS.n7972 9.38145
R17434 VSS.n7899 VSS.n7892 9.38145
R17435 VSS.n9046 VSS.n9045 9.38145
R17436 VSS.n8541 VSS.n269 9.38145
R17437 VSS.n1709 VSS.n1708 9.38145
R17438 VSS.n1223 VSS.n1215 9.38145
R17439 VSS.n2301 VSS.n2300 9.38145
R17440 VSS.n1796 VSS.n1788 9.38145
R17441 VSS.n3509 VSS.n3502 9.38145
R17442 VSS.n3590 VSS.n3582 9.38145
R17443 VSS.n4101 VSS.n4094 9.38145
R17444 VSS.n4182 VSS.n4174 9.38145
R17445 VSS.n4693 VSS.n4686 9.38145
R17446 VSS.n4774 VSS.n4766 9.38145
R17447 VSS.n5285 VSS.n5278 9.38145
R17448 VSS.n5366 VSS.n5358 9.38145
R17449 VSS.n5877 VSS.n5870 9.38145
R17450 VSS.n5958 VSS.n5950 9.38145
R17451 VSS.n6469 VSS.n6462 9.38145
R17452 VSS.n6550 VSS.n6542 9.38145
R17453 VSS.n7045 VSS.n7044 9.38145
R17454 VSS.n2394 VSS.n2386 9.38145
R17455 VSS.n2916 VSS.n2909 9.38145
R17456 VSS.n2991 VSS.n2984 9.38145
R17457 VSS.n189 VSS.n176 9.38145
R17458 VSS.n436 VSS.n435 9.38145
R17459 VSS.n543 VSS.n481 9.38145
R17460 VSS.n1001 VSS.n1000 9.38145
R17461 VSS.n7745 VSS.n7341 9.30555
R17462 VSS.n7601 VSS.n7589 9.30555
R17463 VSS.n8337 VSS.n7755 9.30555
R17464 VSS.n8193 VSS.n8181 9.30555
R17465 VSS.n8925 VSS.n8895 9.30555
R17466 VSS.n8997 VSS.n8771 9.30555
R17467 VSS.n9345 VSS.n3 9.30555
R17468 VSS.n1660 VSS.n1453 9.30555
R17469 VSS.n2160 VSS.n2159 9.30555
R17470 VSS.n2252 VSS.n2026 9.30555
R17471 VSS.n3948 VSS.n3366 9.30555
R17472 VSS.n3803 VSS.n3791 9.30555
R17473 VSS.n4540 VSS.n3958 9.30555
R17474 VSS.n4395 VSS.n4383 9.30555
R17475 VSS.n5132 VSS.n4550 9.30555
R17476 VSS.n4987 VSS.n4975 9.30555
R17477 VSS.n5724 VSS.n5142 9.30555
R17478 VSS.n5579 VSS.n5567 9.30555
R17479 VSS.n6316 VSS.n5734 9.30555
R17480 VSS.n6171 VSS.n6159 9.30555
R17481 VSS.n6908 VSS.n6326 9.30555
R17482 VSS.n6763 VSS.n6751 9.30555
R17483 VSS.n2758 VSS.n2757 9.30555
R17484 VSS.n6996 VSS.n2624 9.30555
R17485 VSS.n3356 VSS.n2773 9.30555
R17486 VSS.n3211 VSS.n3199 9.30555
R17487 VSS.n9316 VSS.n40 9.30555
R17488 VSS.n9171 VSS.n9159 9.30555
R17489 VSS.n9337 VSS.n28 9.30555
R17490 VSS.n815 VSS.n616 9.30555
R17491 VSS.n7326 VSS.n7325 9.30555
R17492 VSS.n8424 VSS.n7192 9.30555
R17493 VSS.n7142 VSS.n7141 9.3005
R17494 VSS.n7163 VSS.n7162 9.3005
R17495 VSS.n7103 VSS.n7102 9.3005
R17496 VSS.n7184 VSS.n7183 9.3005
R17497 VSS.n1090 VSS.n1089 9.3005
R17498 VSS.n1111 VSS.n1110 9.3005
R17499 VSS.n1052 VSS.n1051 9.3005
R17500 VSS.n1133 VSS.n1132 9.3005
R17501 VSS.n7650 VSS.n7649 9.3005
R17502 VSS.n7343 VSS.n7342 9.3005
R17503 VSS.n7700 VSS.n7369 9.3005
R17504 VSS.n7377 VSS.n7375 9.3005
R17505 VSS.n7665 VSS.n7664 9.3005
R17506 VSS.n7719 VSS.n7357 9.3005
R17507 VSS.n7721 VSS.n7720 9.3005
R17508 VSS.n7703 VSS.n7701 9.3005
R17509 VSS.n7651 VSS.n7389 9.3005
R17510 VSS.n7663 VSS.n7382 9.3005
R17511 VSS.n7678 VSS.n7677 9.3005
R17512 VSS.n7593 VSS.n7409 9.3005
R17513 VSS.n7630 VSS.n7400 9.3005
R17514 VSS.n7632 VSS.n7631 9.3005
R17515 VSS.n7513 VSS.n7512 9.3005
R17516 VSS.n7551 VSS.n7550 9.3005
R17517 VSS.n7420 VSS.n7419 9.3005
R17518 VSS.n7579 VSS.n7578 9.3005
R17519 VSS.n7558 VSS.n7557 9.3005
R17520 VSS.n7559 VSS.n7558 9.3005
R17521 VSS.n7560 VSS.n7559 9.3005
R17522 VSS.n7526 VSS.n7525 9.3005
R17523 VSS.n7526 VSS.n7454 9.3005
R17524 VSS.n7454 VSS.n7453 9.3005
R17525 VSS.n7506 VSS.n7505 9.3005
R17526 VSS.n7507 VSS.n7506 9.3005
R17527 VSS.n7566 VSS.n7565 9.3005
R17528 VSS.n7565 VSS.n7418 9.3005
R17529 VSS.n7418 VSS.n7417 9.3005
R17530 VSS.n7608 VSS.n7607 9.3005
R17531 VSS.n7607 VSS.n7606 9.3005
R17532 VSS.n7480 VSS.n7478 9.3005
R17533 VSS.n7736 VSS.n7735 9.3005
R17534 VSS.n7736 VSS.n7348 9.3005
R17535 VSS.n7348 VSS.n7347 9.3005
R17536 VSS.n7713 VSS.n7712 9.3005
R17537 VSS.n7714 VSS.n7713 9.3005
R17538 VSS.n7715 VSS.n7714 9.3005
R17539 VSS.n7681 VSS.n7370 9.3005
R17540 VSS.n7371 VSS.n7370 9.3005
R17541 VSS.n7695 VSS.n7371 9.3005
R17542 VSS.n7640 VSS.n7639 9.3005
R17543 VSS.n7640 VSS.n7392 9.3005
R17544 VSS.n7644 VSS.n7392 9.3005
R17545 VSS.n7660 VSS.n7383 9.3005
R17546 VSS.n7383 VSS.n7373 9.3005
R17547 VSS.n7373 VSS.n7372 9.3005
R17548 VSS.n7745 VSS.n7744 9.3005
R17549 VSS.n7744 VSS.n7743 9.3005
R17550 VSS.n7601 VSS.n7600 9.3005
R17551 VSS.n7600 VSS.n7599 9.3005
R17552 VSS.n7402 VSS.n7401 9.3005
R17553 VSS.n7592 VSS.n7401 9.3005
R17554 VSS.n7592 VSS.n7591 9.3005
R17555 VSS.n7956 VSS.n7952 9.3005
R17556 VSS.n7934 VSS.n7933 9.3005
R17557 VSS.n7914 VSS.n7913 9.3005
R17558 VSS.n7917 VSS.n7916 9.3005
R17559 VSS.n8242 VSS.n8241 9.3005
R17560 VSS.n7757 VSS.n7756 9.3005
R17561 VSS.n8292 VSS.n7783 9.3005
R17562 VSS.n7791 VSS.n7789 9.3005
R17563 VSS.n8257 VSS.n8256 9.3005
R17564 VSS.n8311 VSS.n7771 9.3005
R17565 VSS.n8313 VSS.n8312 9.3005
R17566 VSS.n8295 VSS.n8293 9.3005
R17567 VSS.n8243 VSS.n7803 9.3005
R17568 VSS.n8255 VSS.n7796 9.3005
R17569 VSS.n8270 VSS.n8269 9.3005
R17570 VSS.n8185 VSS.n7823 9.3005
R17571 VSS.n8222 VSS.n7814 9.3005
R17572 VSS.n8224 VSS.n8223 9.3005
R17573 VSS.n8105 VSS.n8104 9.3005
R17574 VSS.n8143 VSS.n8142 9.3005
R17575 VSS.n7834 VSS.n7833 9.3005
R17576 VSS.n8171 VSS.n8170 9.3005
R17577 VSS.n8150 VSS.n8149 9.3005
R17578 VSS.n8151 VSS.n8150 9.3005
R17579 VSS.n8152 VSS.n8151 9.3005
R17580 VSS.n8118 VSS.n8117 9.3005
R17581 VSS.n8118 VSS.n7868 9.3005
R17582 VSS.n7868 VSS.n7867 9.3005
R17583 VSS.n8098 VSS.n8097 9.3005
R17584 VSS.n8099 VSS.n8098 9.3005
R17585 VSS.n8158 VSS.n8157 9.3005
R17586 VSS.n8157 VSS.n7832 9.3005
R17587 VSS.n7832 VSS.n7831 9.3005
R17588 VSS.n8200 VSS.n8199 9.3005
R17589 VSS.n8199 VSS.n8198 9.3005
R17590 VSS.n7894 VSS.n7892 9.3005
R17591 VSS.n8328 VSS.n8327 9.3005
R17592 VSS.n8328 VSS.n7762 9.3005
R17593 VSS.n7762 VSS.n7761 9.3005
R17594 VSS.n8305 VSS.n8304 9.3005
R17595 VSS.n8306 VSS.n8305 9.3005
R17596 VSS.n8307 VSS.n8306 9.3005
R17597 VSS.n8273 VSS.n7784 9.3005
R17598 VSS.n7785 VSS.n7784 9.3005
R17599 VSS.n8287 VSS.n7785 9.3005
R17600 VSS.n8232 VSS.n8231 9.3005
R17601 VSS.n8232 VSS.n7806 9.3005
R17602 VSS.n8236 VSS.n7806 9.3005
R17603 VSS.n8252 VSS.n7797 9.3005
R17604 VSS.n7797 VSS.n7787 9.3005
R17605 VSS.n7787 VSS.n7786 9.3005
R17606 VSS.n8337 VSS.n8336 9.3005
R17607 VSS.n8336 VSS.n8335 9.3005
R17608 VSS.n8193 VSS.n8192 9.3005
R17609 VSS.n8192 VSS.n8191 9.3005
R17610 VSS.n7816 VSS.n7815 9.3005
R17611 VSS.n8184 VSS.n7815 9.3005
R17612 VSS.n8184 VSS.n8183 9.3005
R17613 VSS.n8721 VSS.n8720 9.3005
R17614 VSS.n8742 VSS.n8741 9.3005
R17615 VSS.n8682 VSS.n8681 9.3005
R17616 VSS.n8763 VSS.n8762 9.3005
R17617 VSS.n8972 VSS.n8971 9.3005
R17618 VSS.n8898 VSS.n8897 9.3005
R17619 VSS.n8953 VSS.n8952 9.3005
R17620 VSS.n8865 VSS.n8859 9.3005
R17621 VSS.n8820 VSS.n8818 9.3005
R17622 VSS.n8945 VSS.n8944 9.3005
R17623 VSS.n8943 VSS.n8882 9.3005
R17624 VSS.n8951 VSS.n8850 9.3005
R17625 VSS.n8973 VSS.n8805 9.3005
R17626 VSS.n8839 VSS.n8838 9.3005
R17627 VSS.n8867 VSS.n8866 9.3005
R17628 VSS.n8786 VSS.n8785 9.3005
R17629 VSS.n8827 VSS.n8826 9.3005
R17630 VSS.n8828 VSS.n8802 9.3005
R17631 VSS.n253 VSS.n249 9.3005
R17632 VSS.n231 VSS.n230 9.3005
R17633 VSS.n211 VSS.n210 9.3005
R17634 VSS.n214 VSS.n213 9.3005
R17635 VSS.n8605 VSS.n8604 9.3005
R17636 VSS.n8604 VSS.n8603 9.3005
R17637 VSS.n8603 VSS.n8602 9.3005
R17638 VSS.n8571 VSS.n252 9.3005
R17639 VSS.n8571 VSS.n8570 9.3005
R17640 VSS.n8570 VSS.n8569 9.3005
R17641 VSS.n8560 VSS.n258 9.3005
R17642 VSS.n258 VSS.n257 9.3005
R17643 VSS.n8628 VSS.n8627 9.3005
R17644 VSS.n8629 VSS.n8628 9.3005
R17645 VSS.n8630 VSS.n8629 9.3005
R17646 VSS.n8635 VSS.n8634 9.3005
R17647 VSS.n8634 VSS.n192 9.3005
R17648 VSS.n8536 VSS.n269 9.3005
R17649 VSS.n1403 VSS.n1402 9.3005
R17650 VSS.n1424 VSS.n1423 9.3005
R17651 VSS.n1364 VSS.n1363 9.3005
R17652 VSS.n1445 VSS.n1444 9.3005
R17653 VSS.n1430 VSS.n1429 9.3005
R17654 VSS.n1431 VSS.n1430 9.3005
R17655 VSS.n1432 VSS.n1431 9.3005
R17656 VSS.n1411 VSS.n1377 9.3005
R17657 VSS.n1411 VSS.n1410 9.3005
R17658 VSS.n1410 VSS.n1409 9.3005
R17659 VSS.n1396 VSS.n1380 9.3005
R17660 VSS.n1380 VSS.n1379 9.3005
R17661 VSS.n1436 VSS.n1367 9.3005
R17662 VSS.n1436 VSS.n1362 9.3005
R17663 VSS.n1362 VSS.n1361 9.3005
R17664 VSS.n1667 VSS.n1666 9.3005
R17665 VSS.n1666 VSS.n1665 9.3005
R17666 VSS.n1710 VSS.n1709 9.3005
R17667 VSS.n1631 VSS.n1630 9.3005
R17668 VSS.n5 VSS.n4 9.3005
R17669 VSS.n1612 VSS.n1611 9.3005
R17670 VSS.n1508 VSS.n1506 9.3005
R17671 VSS.n1526 VSS.n1525 9.3005
R17672 VSS.n1593 VSS.n1564 9.3005
R17673 VSS.n1593 VSS.n1592 9.3005
R17674 VSS.n1592 VSS.n1591 9.3005
R17675 VSS.n1585 VSS.n1543 9.3005
R17676 VSS.n1565 VSS.n1551 9.3005
R17677 VSS.n1542 VSS.n1538 9.3005
R17678 VSS.n1584 VSS.n1538 9.3005
R17679 VSS.n1584 VSS.n1570 9.3005
R17680 VSS.n1610 VSS.n1536 9.3005
R17681 VSS.n1578 VSS.n1577 9.3005
R17682 VSS.n1578 VSS.n1504 9.3005
R17683 VSS.n1504 VSS.n1503 9.3005
R17684 VSS.n1638 VSS.n1637 9.3005
R17685 VSS.n1639 VSS.n1638 9.3005
R17686 VSS.n1640 VSS.n1639 9.3005
R17687 VSS.n1632 VSS.n1499 9.3005
R17688 VSS.n1521 VSS.n1501 9.3005
R17689 VSS.n1502 VSS.n1501 9.3005
R17690 VSS.n1625 VSS.n1502 9.3005
R17691 VSS.n1524 VSS.n1513 9.3005
R17692 VSS.n1573 VSS.n1572 9.3005
R17693 VSS.n9345 VSS.n9344 9.3005
R17694 VSS.n9344 VSS.n9343 9.3005
R17695 VSS.n1467 VSS.n1466 9.3005
R17696 VSS.n1660 VSS.n1659 9.3005
R17697 VSS.n1659 VSS.n1658 9.3005
R17698 VSS.n1653 VSS.n1652 9.3005
R17699 VSS.n1653 VSS.n1456 9.3005
R17700 VSS.n1456 VSS.n1455 9.3005
R17701 VSS.n1647 VSS.n1646 9.3005
R17702 VSS.n1645 VSS.n1482 9.3005
R17703 VSS.n1199 VSS.n1195 9.3005
R17704 VSS.n1177 VSS.n1176 9.3005
R17705 VSS.n1157 VSS.n1156 9.3005
R17706 VSS.n1160 VSS.n1159 9.3005
R17707 VSS.n1287 VSS.n1286 9.3005
R17708 VSS.n1286 VSS.n1285 9.3005
R17709 VSS.n1285 VSS.n1284 9.3005
R17710 VSS.n1253 VSS.n1198 9.3005
R17711 VSS.n1253 VSS.n1252 9.3005
R17712 VSS.n1252 VSS.n1251 9.3005
R17713 VSS.n1242 VSS.n1204 9.3005
R17714 VSS.n1204 VSS.n1203 9.3005
R17715 VSS.n1310 VSS.n1309 9.3005
R17716 VSS.n1311 VSS.n1310 9.3005
R17717 VSS.n1312 VSS.n1311 9.3005
R17718 VSS.n1317 VSS.n1316 9.3005
R17719 VSS.n1316 VSS.n1138 9.3005
R17720 VSS.n1218 VSS.n1215 9.3005
R17721 VSS.n1976 VSS.n1975 9.3005
R17722 VSS.n1997 VSS.n1996 9.3005
R17723 VSS.n1937 VSS.n1936 9.3005
R17724 VSS.n2018 VSS.n2017 9.3005
R17725 VSS.n2003 VSS.n2002 9.3005
R17726 VSS.n2004 VSS.n2003 9.3005
R17727 VSS.n2005 VSS.n2004 9.3005
R17728 VSS.n1984 VSS.n1950 9.3005
R17729 VSS.n1984 VSS.n1983 9.3005
R17730 VSS.n1983 VSS.n1982 9.3005
R17731 VSS.n1969 VSS.n1953 9.3005
R17732 VSS.n1953 VSS.n1952 9.3005
R17733 VSS.n2009 VSS.n1940 9.3005
R17734 VSS.n2009 VSS.n1935 9.3005
R17735 VSS.n1935 VSS.n1934 9.3005
R17736 VSS.n2259 VSS.n2258 9.3005
R17737 VSS.n2258 VSS.n2257 9.3005
R17738 VSS.n2302 VSS.n2301 9.3005
R17739 VSS.n2223 VSS.n2222 9.3005
R17740 VSS.n2178 VSS.n2177 9.3005
R17741 VSS.n2204 VSS.n2203 9.3005
R17742 VSS.n2081 VSS.n2079 9.3005
R17743 VSS.n2099 VSS.n2098 9.3005
R17744 VSS.n2185 VSS.n2125 9.3005
R17745 VSS.n2185 VSS.n2184 9.3005
R17746 VSS.n2184 VSS.n2183 9.3005
R17747 VSS.n2145 VSS.n2116 9.3005
R17748 VSS.n2126 VSS.n2124 9.3005
R17749 VSS.n2115 VSS.n2111 9.3005
R17750 VSS.n2144 VSS.n2111 9.3005
R17751 VSS.n2144 VSS.n2130 9.3005
R17752 VSS.n2202 VSS.n2109 9.3005
R17753 VSS.n2138 VSS.n2137 9.3005
R17754 VSS.n2138 VSS.n2077 9.3005
R17755 VSS.n2077 VSS.n2076 9.3005
R17756 VSS.n2230 VSS.n2229 9.3005
R17757 VSS.n2231 VSS.n2230 9.3005
R17758 VSS.n2232 VSS.n2231 9.3005
R17759 VSS.n2224 VSS.n2072 9.3005
R17760 VSS.n2094 VSS.n2074 9.3005
R17761 VSS.n2075 VSS.n2074 9.3005
R17762 VSS.n2217 VSS.n2075 9.3005
R17763 VSS.n2097 VSS.n2086 9.3005
R17764 VSS.n2133 VSS.n2132 9.3005
R17765 VSS.n2159 VSS.n2151 9.3005
R17766 VSS.n2151 VSS.n2150 9.3005
R17767 VSS.n2040 VSS.n2039 9.3005
R17768 VSS.n2252 VSS.n2251 9.3005
R17769 VSS.n2251 VSS.n2250 9.3005
R17770 VSS.n2245 VSS.n2244 9.3005
R17771 VSS.n2245 VSS.n2029 9.3005
R17772 VSS.n2029 VSS.n2028 9.3005
R17773 VSS.n2239 VSS.n2238 9.3005
R17774 VSS.n2237 VSS.n2055 9.3005
R17775 VSS.n1772 VSS.n1768 9.3005
R17776 VSS.n1750 VSS.n1749 9.3005
R17777 VSS.n1730 VSS.n1729 9.3005
R17778 VSS.n1733 VSS.n1732 9.3005
R17779 VSS.n1860 VSS.n1859 9.3005
R17780 VSS.n1859 VSS.n1858 9.3005
R17781 VSS.n1858 VSS.n1857 9.3005
R17782 VSS.n1826 VSS.n1771 9.3005
R17783 VSS.n1826 VSS.n1825 9.3005
R17784 VSS.n1825 VSS.n1824 9.3005
R17785 VSS.n1815 VSS.n1777 9.3005
R17786 VSS.n1777 VSS.n1776 9.3005
R17787 VSS.n1883 VSS.n1882 9.3005
R17788 VSS.n1884 VSS.n1883 9.3005
R17789 VSS.n1885 VSS.n1884 9.3005
R17790 VSS.n1890 VSS.n1889 9.3005
R17791 VSS.n1889 VSS.n1711 9.3005
R17792 VSS.n1791 VSS.n1788 9.3005
R17793 VSS.n3715 VSS.n3714 9.3005
R17794 VSS.n3753 VSS.n3752 9.3005
R17795 VSS.n3444 VSS.n3443 9.3005
R17796 VSS.n3781 VSS.n3780 9.3005
R17797 VSS.n3760 VSS.n3759 9.3005
R17798 VSS.n3761 VSS.n3760 9.3005
R17799 VSS.n3762 VSS.n3761 9.3005
R17800 VSS.n3728 VSS.n3727 9.3005
R17801 VSS.n3728 VSS.n3478 9.3005
R17802 VSS.n3478 VSS.n3477 9.3005
R17803 VSS.n3708 VSS.n3707 9.3005
R17804 VSS.n3709 VSS.n3708 9.3005
R17805 VSS.n3768 VSS.n3767 9.3005
R17806 VSS.n3767 VSS.n3442 9.3005
R17807 VSS.n3442 VSS.n3441 9.3005
R17808 VSS.n3810 VSS.n3809 9.3005
R17809 VSS.n3809 VSS.n3808 9.3005
R17810 VSS.n3504 VSS.n3502 9.3005
R17811 VSS.n3852 VSS.n3851 9.3005
R17812 VSS.n3368 VSS.n3367 9.3005
R17813 VSS.n3902 VSS.n3393 9.3005
R17814 VSS.n3401 VSS.n3399 9.3005
R17815 VSS.n3867 VSS.n3866 9.3005
R17816 VSS.n3939 VSS.n3938 9.3005
R17817 VSS.n3939 VSS.n3373 9.3005
R17818 VSS.n3373 VSS.n3372 9.3005
R17819 VSS.n3921 VSS.n3381 9.3005
R17820 VSS.n3923 VSS.n3922 9.3005
R17821 VSS.n3915 VSS.n3914 9.3005
R17822 VSS.n3916 VSS.n3915 9.3005
R17823 VSS.n3917 VSS.n3916 9.3005
R17824 VSS.n3905 VSS.n3903 9.3005
R17825 VSS.n3883 VSS.n3394 9.3005
R17826 VSS.n3395 VSS.n3394 9.3005
R17827 VSS.n3897 VSS.n3395 9.3005
R17828 VSS.n3842 VSS.n3841 9.3005
R17829 VSS.n3842 VSS.n3416 9.3005
R17830 VSS.n3846 VSS.n3416 9.3005
R17831 VSS.n3853 VSS.n3413 9.3005
R17832 VSS.n3862 VSS.n3407 9.3005
R17833 VSS.n3407 VSS.n3397 9.3005
R17834 VSS.n3397 VSS.n3396 9.3005
R17835 VSS.n3865 VSS.n3406 9.3005
R17836 VSS.n3880 VSS.n3879 9.3005
R17837 VSS.n3948 VSS.n3947 9.3005
R17838 VSS.n3947 VSS.n3946 9.3005
R17839 VSS.n3795 VSS.n3433 9.3005
R17840 VSS.n3803 VSS.n3802 9.3005
R17841 VSS.n3802 VSS.n3801 9.3005
R17842 VSS.n3426 VSS.n3425 9.3005
R17843 VSS.n3794 VSS.n3425 9.3005
R17844 VSS.n3794 VSS.n3793 9.3005
R17845 VSS.n3832 VSS.n3424 9.3005
R17846 VSS.n3834 VSS.n3833 9.3005
R17847 VSS.n3566 VSS.n3562 9.3005
R17848 VSS.n3544 VSS.n3543 9.3005
R17849 VSS.n3524 VSS.n3523 9.3005
R17850 VSS.n3527 VSS.n3526 9.3005
R17851 VSS.n3654 VSS.n3653 9.3005
R17852 VSS.n3653 VSS.n3652 9.3005
R17853 VSS.n3652 VSS.n3651 9.3005
R17854 VSS.n3620 VSS.n3565 9.3005
R17855 VSS.n3620 VSS.n3619 9.3005
R17856 VSS.n3619 VSS.n3618 9.3005
R17857 VSS.n3609 VSS.n3571 9.3005
R17858 VSS.n3571 VSS.n3570 9.3005
R17859 VSS.n3677 VSS.n3676 9.3005
R17860 VSS.n3678 VSS.n3677 9.3005
R17861 VSS.n3679 VSS.n3678 9.3005
R17862 VSS.n3684 VSS.n3683 9.3005
R17863 VSS.n3683 VSS.n2303 9.3005
R17864 VSS.n3585 VSS.n3582 9.3005
R17865 VSS.n4307 VSS.n4306 9.3005
R17866 VSS.n4345 VSS.n4344 9.3005
R17867 VSS.n4036 VSS.n4035 9.3005
R17868 VSS.n4373 VSS.n4372 9.3005
R17869 VSS.n4352 VSS.n4351 9.3005
R17870 VSS.n4353 VSS.n4352 9.3005
R17871 VSS.n4354 VSS.n4353 9.3005
R17872 VSS.n4320 VSS.n4319 9.3005
R17873 VSS.n4320 VSS.n4070 9.3005
R17874 VSS.n4070 VSS.n4069 9.3005
R17875 VSS.n4300 VSS.n4299 9.3005
R17876 VSS.n4301 VSS.n4300 9.3005
R17877 VSS.n4360 VSS.n4359 9.3005
R17878 VSS.n4359 VSS.n4034 9.3005
R17879 VSS.n4034 VSS.n4033 9.3005
R17880 VSS.n4402 VSS.n4401 9.3005
R17881 VSS.n4401 VSS.n4400 9.3005
R17882 VSS.n4096 VSS.n4094 9.3005
R17883 VSS.n4444 VSS.n4443 9.3005
R17884 VSS.n3960 VSS.n3959 9.3005
R17885 VSS.n4494 VSS.n3985 9.3005
R17886 VSS.n3993 VSS.n3991 9.3005
R17887 VSS.n4459 VSS.n4458 9.3005
R17888 VSS.n4531 VSS.n4530 9.3005
R17889 VSS.n4531 VSS.n3965 9.3005
R17890 VSS.n3965 VSS.n3964 9.3005
R17891 VSS.n4513 VSS.n3973 9.3005
R17892 VSS.n4515 VSS.n4514 9.3005
R17893 VSS.n4507 VSS.n4506 9.3005
R17894 VSS.n4508 VSS.n4507 9.3005
R17895 VSS.n4509 VSS.n4508 9.3005
R17896 VSS.n4497 VSS.n4495 9.3005
R17897 VSS.n4475 VSS.n3986 9.3005
R17898 VSS.n3987 VSS.n3986 9.3005
R17899 VSS.n4489 VSS.n3987 9.3005
R17900 VSS.n4434 VSS.n4433 9.3005
R17901 VSS.n4434 VSS.n4008 9.3005
R17902 VSS.n4438 VSS.n4008 9.3005
R17903 VSS.n4445 VSS.n4005 9.3005
R17904 VSS.n4454 VSS.n3999 9.3005
R17905 VSS.n3999 VSS.n3989 9.3005
R17906 VSS.n3989 VSS.n3988 9.3005
R17907 VSS.n4457 VSS.n3998 9.3005
R17908 VSS.n4472 VSS.n4471 9.3005
R17909 VSS.n4540 VSS.n4539 9.3005
R17910 VSS.n4539 VSS.n4538 9.3005
R17911 VSS.n4387 VSS.n4025 9.3005
R17912 VSS.n4395 VSS.n4394 9.3005
R17913 VSS.n4394 VSS.n4393 9.3005
R17914 VSS.n4018 VSS.n4017 9.3005
R17915 VSS.n4386 VSS.n4017 9.3005
R17916 VSS.n4386 VSS.n4385 9.3005
R17917 VSS.n4424 VSS.n4016 9.3005
R17918 VSS.n4426 VSS.n4425 9.3005
R17919 VSS.n4158 VSS.n4154 9.3005
R17920 VSS.n4136 VSS.n4135 9.3005
R17921 VSS.n4116 VSS.n4115 9.3005
R17922 VSS.n4119 VSS.n4118 9.3005
R17923 VSS.n4246 VSS.n4245 9.3005
R17924 VSS.n4245 VSS.n4244 9.3005
R17925 VSS.n4244 VSS.n4243 9.3005
R17926 VSS.n4212 VSS.n4157 9.3005
R17927 VSS.n4212 VSS.n4211 9.3005
R17928 VSS.n4211 VSS.n4210 9.3005
R17929 VSS.n4201 VSS.n4163 9.3005
R17930 VSS.n4163 VSS.n4162 9.3005
R17931 VSS.n4269 VSS.n4268 9.3005
R17932 VSS.n4270 VSS.n4269 9.3005
R17933 VSS.n4271 VSS.n4270 9.3005
R17934 VSS.n4276 VSS.n4275 9.3005
R17935 VSS.n4275 VSS.n2304 9.3005
R17936 VSS.n4177 VSS.n4174 9.3005
R17937 VSS.n4899 VSS.n4898 9.3005
R17938 VSS.n4937 VSS.n4936 9.3005
R17939 VSS.n4628 VSS.n4627 9.3005
R17940 VSS.n4965 VSS.n4964 9.3005
R17941 VSS.n4944 VSS.n4943 9.3005
R17942 VSS.n4945 VSS.n4944 9.3005
R17943 VSS.n4946 VSS.n4945 9.3005
R17944 VSS.n4912 VSS.n4911 9.3005
R17945 VSS.n4912 VSS.n4662 9.3005
R17946 VSS.n4662 VSS.n4661 9.3005
R17947 VSS.n4892 VSS.n4891 9.3005
R17948 VSS.n4893 VSS.n4892 9.3005
R17949 VSS.n4952 VSS.n4951 9.3005
R17950 VSS.n4951 VSS.n4626 9.3005
R17951 VSS.n4626 VSS.n4625 9.3005
R17952 VSS.n4994 VSS.n4993 9.3005
R17953 VSS.n4993 VSS.n4992 9.3005
R17954 VSS.n4688 VSS.n4686 9.3005
R17955 VSS.n5036 VSS.n5035 9.3005
R17956 VSS.n4552 VSS.n4551 9.3005
R17957 VSS.n5086 VSS.n4577 9.3005
R17958 VSS.n4585 VSS.n4583 9.3005
R17959 VSS.n5051 VSS.n5050 9.3005
R17960 VSS.n5123 VSS.n5122 9.3005
R17961 VSS.n5123 VSS.n4557 9.3005
R17962 VSS.n4557 VSS.n4556 9.3005
R17963 VSS.n5105 VSS.n4565 9.3005
R17964 VSS.n5107 VSS.n5106 9.3005
R17965 VSS.n5099 VSS.n5098 9.3005
R17966 VSS.n5100 VSS.n5099 9.3005
R17967 VSS.n5101 VSS.n5100 9.3005
R17968 VSS.n5089 VSS.n5087 9.3005
R17969 VSS.n5067 VSS.n4578 9.3005
R17970 VSS.n4579 VSS.n4578 9.3005
R17971 VSS.n5081 VSS.n4579 9.3005
R17972 VSS.n5026 VSS.n5025 9.3005
R17973 VSS.n5026 VSS.n4600 9.3005
R17974 VSS.n5030 VSS.n4600 9.3005
R17975 VSS.n5037 VSS.n4597 9.3005
R17976 VSS.n5046 VSS.n4591 9.3005
R17977 VSS.n4591 VSS.n4581 9.3005
R17978 VSS.n4581 VSS.n4580 9.3005
R17979 VSS.n5049 VSS.n4590 9.3005
R17980 VSS.n5064 VSS.n5063 9.3005
R17981 VSS.n5132 VSS.n5131 9.3005
R17982 VSS.n5131 VSS.n5130 9.3005
R17983 VSS.n4979 VSS.n4617 9.3005
R17984 VSS.n4987 VSS.n4986 9.3005
R17985 VSS.n4986 VSS.n4985 9.3005
R17986 VSS.n4610 VSS.n4609 9.3005
R17987 VSS.n4978 VSS.n4609 9.3005
R17988 VSS.n4978 VSS.n4977 9.3005
R17989 VSS.n5016 VSS.n4608 9.3005
R17990 VSS.n5018 VSS.n5017 9.3005
R17991 VSS.n4750 VSS.n4746 9.3005
R17992 VSS.n4728 VSS.n4727 9.3005
R17993 VSS.n4708 VSS.n4707 9.3005
R17994 VSS.n4711 VSS.n4710 9.3005
R17995 VSS.n4838 VSS.n4837 9.3005
R17996 VSS.n4837 VSS.n4836 9.3005
R17997 VSS.n4836 VSS.n4835 9.3005
R17998 VSS.n4804 VSS.n4749 9.3005
R17999 VSS.n4804 VSS.n4803 9.3005
R18000 VSS.n4803 VSS.n4802 9.3005
R18001 VSS.n4793 VSS.n4755 9.3005
R18002 VSS.n4755 VSS.n4754 9.3005
R18003 VSS.n4861 VSS.n4860 9.3005
R18004 VSS.n4862 VSS.n4861 9.3005
R18005 VSS.n4863 VSS.n4862 9.3005
R18006 VSS.n4868 VSS.n4867 9.3005
R18007 VSS.n4867 VSS.n2305 9.3005
R18008 VSS.n4769 VSS.n4766 9.3005
R18009 VSS.n5491 VSS.n5490 9.3005
R18010 VSS.n5529 VSS.n5528 9.3005
R18011 VSS.n5220 VSS.n5219 9.3005
R18012 VSS.n5557 VSS.n5556 9.3005
R18013 VSS.n5536 VSS.n5535 9.3005
R18014 VSS.n5537 VSS.n5536 9.3005
R18015 VSS.n5538 VSS.n5537 9.3005
R18016 VSS.n5504 VSS.n5503 9.3005
R18017 VSS.n5504 VSS.n5254 9.3005
R18018 VSS.n5254 VSS.n5253 9.3005
R18019 VSS.n5484 VSS.n5483 9.3005
R18020 VSS.n5485 VSS.n5484 9.3005
R18021 VSS.n5544 VSS.n5543 9.3005
R18022 VSS.n5543 VSS.n5218 9.3005
R18023 VSS.n5218 VSS.n5217 9.3005
R18024 VSS.n5586 VSS.n5585 9.3005
R18025 VSS.n5585 VSS.n5584 9.3005
R18026 VSS.n5280 VSS.n5278 9.3005
R18027 VSS.n5628 VSS.n5627 9.3005
R18028 VSS.n5144 VSS.n5143 9.3005
R18029 VSS.n5678 VSS.n5169 9.3005
R18030 VSS.n5177 VSS.n5175 9.3005
R18031 VSS.n5643 VSS.n5642 9.3005
R18032 VSS.n5715 VSS.n5714 9.3005
R18033 VSS.n5715 VSS.n5149 9.3005
R18034 VSS.n5149 VSS.n5148 9.3005
R18035 VSS.n5697 VSS.n5157 9.3005
R18036 VSS.n5699 VSS.n5698 9.3005
R18037 VSS.n5691 VSS.n5690 9.3005
R18038 VSS.n5692 VSS.n5691 9.3005
R18039 VSS.n5693 VSS.n5692 9.3005
R18040 VSS.n5681 VSS.n5679 9.3005
R18041 VSS.n5659 VSS.n5170 9.3005
R18042 VSS.n5171 VSS.n5170 9.3005
R18043 VSS.n5673 VSS.n5171 9.3005
R18044 VSS.n5618 VSS.n5617 9.3005
R18045 VSS.n5618 VSS.n5192 9.3005
R18046 VSS.n5622 VSS.n5192 9.3005
R18047 VSS.n5629 VSS.n5189 9.3005
R18048 VSS.n5638 VSS.n5183 9.3005
R18049 VSS.n5183 VSS.n5173 9.3005
R18050 VSS.n5173 VSS.n5172 9.3005
R18051 VSS.n5641 VSS.n5182 9.3005
R18052 VSS.n5656 VSS.n5655 9.3005
R18053 VSS.n5724 VSS.n5723 9.3005
R18054 VSS.n5723 VSS.n5722 9.3005
R18055 VSS.n5571 VSS.n5209 9.3005
R18056 VSS.n5579 VSS.n5578 9.3005
R18057 VSS.n5578 VSS.n5577 9.3005
R18058 VSS.n5202 VSS.n5201 9.3005
R18059 VSS.n5570 VSS.n5201 9.3005
R18060 VSS.n5570 VSS.n5569 9.3005
R18061 VSS.n5608 VSS.n5200 9.3005
R18062 VSS.n5610 VSS.n5609 9.3005
R18063 VSS.n5342 VSS.n5338 9.3005
R18064 VSS.n5320 VSS.n5319 9.3005
R18065 VSS.n5300 VSS.n5299 9.3005
R18066 VSS.n5303 VSS.n5302 9.3005
R18067 VSS.n5430 VSS.n5429 9.3005
R18068 VSS.n5429 VSS.n5428 9.3005
R18069 VSS.n5428 VSS.n5427 9.3005
R18070 VSS.n5396 VSS.n5341 9.3005
R18071 VSS.n5396 VSS.n5395 9.3005
R18072 VSS.n5395 VSS.n5394 9.3005
R18073 VSS.n5385 VSS.n5347 9.3005
R18074 VSS.n5347 VSS.n5346 9.3005
R18075 VSS.n5453 VSS.n5452 9.3005
R18076 VSS.n5454 VSS.n5453 9.3005
R18077 VSS.n5455 VSS.n5454 9.3005
R18078 VSS.n5460 VSS.n5459 9.3005
R18079 VSS.n5459 VSS.n2306 9.3005
R18080 VSS.n5361 VSS.n5358 9.3005
R18081 VSS.n6083 VSS.n6082 9.3005
R18082 VSS.n6121 VSS.n6120 9.3005
R18083 VSS.n5812 VSS.n5811 9.3005
R18084 VSS.n6149 VSS.n6148 9.3005
R18085 VSS.n6128 VSS.n6127 9.3005
R18086 VSS.n6129 VSS.n6128 9.3005
R18087 VSS.n6130 VSS.n6129 9.3005
R18088 VSS.n6096 VSS.n6095 9.3005
R18089 VSS.n6096 VSS.n5846 9.3005
R18090 VSS.n5846 VSS.n5845 9.3005
R18091 VSS.n6076 VSS.n6075 9.3005
R18092 VSS.n6077 VSS.n6076 9.3005
R18093 VSS.n6136 VSS.n6135 9.3005
R18094 VSS.n6135 VSS.n5810 9.3005
R18095 VSS.n5810 VSS.n5809 9.3005
R18096 VSS.n6178 VSS.n6177 9.3005
R18097 VSS.n6177 VSS.n6176 9.3005
R18098 VSS.n5872 VSS.n5870 9.3005
R18099 VSS.n6220 VSS.n6219 9.3005
R18100 VSS.n5736 VSS.n5735 9.3005
R18101 VSS.n6270 VSS.n5761 9.3005
R18102 VSS.n5769 VSS.n5767 9.3005
R18103 VSS.n6235 VSS.n6234 9.3005
R18104 VSS.n6307 VSS.n6306 9.3005
R18105 VSS.n6307 VSS.n5741 9.3005
R18106 VSS.n5741 VSS.n5740 9.3005
R18107 VSS.n6289 VSS.n5749 9.3005
R18108 VSS.n6291 VSS.n6290 9.3005
R18109 VSS.n6283 VSS.n6282 9.3005
R18110 VSS.n6284 VSS.n6283 9.3005
R18111 VSS.n6285 VSS.n6284 9.3005
R18112 VSS.n6273 VSS.n6271 9.3005
R18113 VSS.n6251 VSS.n5762 9.3005
R18114 VSS.n5763 VSS.n5762 9.3005
R18115 VSS.n6265 VSS.n5763 9.3005
R18116 VSS.n6210 VSS.n6209 9.3005
R18117 VSS.n6210 VSS.n5784 9.3005
R18118 VSS.n6214 VSS.n5784 9.3005
R18119 VSS.n6221 VSS.n5781 9.3005
R18120 VSS.n6230 VSS.n5775 9.3005
R18121 VSS.n5775 VSS.n5765 9.3005
R18122 VSS.n5765 VSS.n5764 9.3005
R18123 VSS.n6233 VSS.n5774 9.3005
R18124 VSS.n6248 VSS.n6247 9.3005
R18125 VSS.n6316 VSS.n6315 9.3005
R18126 VSS.n6315 VSS.n6314 9.3005
R18127 VSS.n6163 VSS.n5801 9.3005
R18128 VSS.n6171 VSS.n6170 9.3005
R18129 VSS.n6170 VSS.n6169 9.3005
R18130 VSS.n5794 VSS.n5793 9.3005
R18131 VSS.n6162 VSS.n5793 9.3005
R18132 VSS.n6162 VSS.n6161 9.3005
R18133 VSS.n6200 VSS.n5792 9.3005
R18134 VSS.n6202 VSS.n6201 9.3005
R18135 VSS.n5934 VSS.n5930 9.3005
R18136 VSS.n5912 VSS.n5911 9.3005
R18137 VSS.n5892 VSS.n5891 9.3005
R18138 VSS.n5895 VSS.n5894 9.3005
R18139 VSS.n6022 VSS.n6021 9.3005
R18140 VSS.n6021 VSS.n6020 9.3005
R18141 VSS.n6020 VSS.n6019 9.3005
R18142 VSS.n5988 VSS.n5933 9.3005
R18143 VSS.n5988 VSS.n5987 9.3005
R18144 VSS.n5987 VSS.n5986 9.3005
R18145 VSS.n5977 VSS.n5939 9.3005
R18146 VSS.n5939 VSS.n5938 9.3005
R18147 VSS.n6045 VSS.n6044 9.3005
R18148 VSS.n6046 VSS.n6045 9.3005
R18149 VSS.n6047 VSS.n6046 9.3005
R18150 VSS.n6052 VSS.n6051 9.3005
R18151 VSS.n6051 VSS.n2307 9.3005
R18152 VSS.n5953 VSS.n5950 9.3005
R18153 VSS.n6675 VSS.n6674 9.3005
R18154 VSS.n6713 VSS.n6712 9.3005
R18155 VSS.n6404 VSS.n6403 9.3005
R18156 VSS.n6741 VSS.n6740 9.3005
R18157 VSS.n6720 VSS.n6719 9.3005
R18158 VSS.n6721 VSS.n6720 9.3005
R18159 VSS.n6722 VSS.n6721 9.3005
R18160 VSS.n6688 VSS.n6687 9.3005
R18161 VSS.n6688 VSS.n6438 9.3005
R18162 VSS.n6438 VSS.n6437 9.3005
R18163 VSS.n6668 VSS.n6667 9.3005
R18164 VSS.n6669 VSS.n6668 9.3005
R18165 VSS.n6728 VSS.n6727 9.3005
R18166 VSS.n6727 VSS.n6402 9.3005
R18167 VSS.n6402 VSS.n6401 9.3005
R18168 VSS.n6770 VSS.n6769 9.3005
R18169 VSS.n6769 VSS.n6768 9.3005
R18170 VSS.n6464 VSS.n6462 9.3005
R18171 VSS.n6812 VSS.n6811 9.3005
R18172 VSS.n6328 VSS.n6327 9.3005
R18173 VSS.n6862 VSS.n6353 9.3005
R18174 VSS.n6361 VSS.n6359 9.3005
R18175 VSS.n6827 VSS.n6826 9.3005
R18176 VSS.n6899 VSS.n6898 9.3005
R18177 VSS.n6899 VSS.n6333 9.3005
R18178 VSS.n6333 VSS.n6332 9.3005
R18179 VSS.n6881 VSS.n6341 9.3005
R18180 VSS.n6883 VSS.n6882 9.3005
R18181 VSS.n6875 VSS.n6874 9.3005
R18182 VSS.n6876 VSS.n6875 9.3005
R18183 VSS.n6877 VSS.n6876 9.3005
R18184 VSS.n6865 VSS.n6863 9.3005
R18185 VSS.n6843 VSS.n6354 9.3005
R18186 VSS.n6355 VSS.n6354 9.3005
R18187 VSS.n6857 VSS.n6355 9.3005
R18188 VSS.n6802 VSS.n6801 9.3005
R18189 VSS.n6802 VSS.n6376 9.3005
R18190 VSS.n6806 VSS.n6376 9.3005
R18191 VSS.n6813 VSS.n6373 9.3005
R18192 VSS.n6822 VSS.n6367 9.3005
R18193 VSS.n6367 VSS.n6357 9.3005
R18194 VSS.n6357 VSS.n6356 9.3005
R18195 VSS.n6825 VSS.n6366 9.3005
R18196 VSS.n6840 VSS.n6839 9.3005
R18197 VSS.n6908 VSS.n6907 9.3005
R18198 VSS.n6907 VSS.n6906 9.3005
R18199 VSS.n6755 VSS.n6393 9.3005
R18200 VSS.n6763 VSS.n6762 9.3005
R18201 VSS.n6762 VSS.n6761 9.3005
R18202 VSS.n6386 VSS.n6385 9.3005
R18203 VSS.n6754 VSS.n6385 9.3005
R18204 VSS.n6754 VSS.n6753 9.3005
R18205 VSS.n6792 VSS.n6384 9.3005
R18206 VSS.n6794 VSS.n6793 9.3005
R18207 VSS.n6526 VSS.n6522 9.3005
R18208 VSS.n6504 VSS.n6503 9.3005
R18209 VSS.n6484 VSS.n6483 9.3005
R18210 VSS.n6487 VSS.n6486 9.3005
R18211 VSS.n6614 VSS.n6613 9.3005
R18212 VSS.n6613 VSS.n6612 9.3005
R18213 VSS.n6612 VSS.n6611 9.3005
R18214 VSS.n6580 VSS.n6525 9.3005
R18215 VSS.n6580 VSS.n6579 9.3005
R18216 VSS.n6579 VSS.n6578 9.3005
R18217 VSS.n6569 VSS.n6531 9.3005
R18218 VSS.n6531 VSS.n6530 9.3005
R18219 VSS.n6637 VSS.n6636 9.3005
R18220 VSS.n6638 VSS.n6637 9.3005
R18221 VSS.n6639 VSS.n6638 9.3005
R18222 VSS.n6644 VSS.n6643 9.3005
R18223 VSS.n6643 VSS.n2308 9.3005
R18224 VSS.n6545 VSS.n6542 9.3005
R18225 VSS.n2574 VSS.n2573 9.3005
R18226 VSS.n2595 VSS.n2594 9.3005
R18227 VSS.n2535 VSS.n2534 9.3005
R18228 VSS.n2616 VSS.n2615 9.3005
R18229 VSS.n2601 VSS.n2600 9.3005
R18230 VSS.n2602 VSS.n2601 9.3005
R18231 VSS.n2603 VSS.n2602 9.3005
R18232 VSS.n2582 VSS.n2548 9.3005
R18233 VSS.n2582 VSS.n2581 9.3005
R18234 VSS.n2581 VSS.n2580 9.3005
R18235 VSS.n2567 VSS.n2551 9.3005
R18236 VSS.n2551 VSS.n2550 9.3005
R18237 VSS.n2607 VSS.n2538 9.3005
R18238 VSS.n2607 VSS.n2533 9.3005
R18239 VSS.n2533 VSS.n2532 9.3005
R18240 VSS.n7003 VSS.n7002 9.3005
R18241 VSS.n7002 VSS.n7001 9.3005
R18242 VSS.n7046 VSS.n7045 9.3005
R18243 VSS.n6967 VSS.n6966 9.3005
R18244 VSS.n6922 VSS.n6921 9.3005
R18245 VSS.n6948 VSS.n6947 9.3005
R18246 VSS.n2679 VSS.n2677 9.3005
R18247 VSS.n2697 VSS.n2696 9.3005
R18248 VSS.n6929 VSS.n2723 9.3005
R18249 VSS.n6929 VSS.n6928 9.3005
R18250 VSS.n6928 VSS.n6927 9.3005
R18251 VSS.n2743 VSS.n2714 9.3005
R18252 VSS.n2724 VSS.n2722 9.3005
R18253 VSS.n2713 VSS.n2709 9.3005
R18254 VSS.n2742 VSS.n2709 9.3005
R18255 VSS.n2742 VSS.n2728 9.3005
R18256 VSS.n6946 VSS.n2707 9.3005
R18257 VSS.n2736 VSS.n2735 9.3005
R18258 VSS.n2736 VSS.n2675 9.3005
R18259 VSS.n2675 VSS.n2674 9.3005
R18260 VSS.n6974 VSS.n6973 9.3005
R18261 VSS.n6975 VSS.n6974 9.3005
R18262 VSS.n6976 VSS.n6975 9.3005
R18263 VSS.n6968 VSS.n2670 9.3005
R18264 VSS.n2692 VSS.n2672 9.3005
R18265 VSS.n2673 VSS.n2672 9.3005
R18266 VSS.n6961 VSS.n2673 9.3005
R18267 VSS.n2695 VSS.n2684 9.3005
R18268 VSS.n2731 VSS.n2730 9.3005
R18269 VSS.n2757 VSS.n2749 9.3005
R18270 VSS.n2749 VSS.n2748 9.3005
R18271 VSS.n2638 VSS.n2637 9.3005
R18272 VSS.n6996 VSS.n6995 9.3005
R18273 VSS.n6995 VSS.n6994 9.3005
R18274 VSS.n6989 VSS.n6988 9.3005
R18275 VSS.n6989 VSS.n2627 9.3005
R18276 VSS.n2627 VSS.n2626 9.3005
R18277 VSS.n6983 VSS.n6982 9.3005
R18278 VSS.n6981 VSS.n2653 9.3005
R18279 VSS.n2370 VSS.n2366 9.3005
R18280 VSS.n2348 VSS.n2347 9.3005
R18281 VSS.n2328 VSS.n2327 9.3005
R18282 VSS.n2331 VSS.n2330 9.3005
R18283 VSS.n2458 VSS.n2457 9.3005
R18284 VSS.n2457 VSS.n2456 9.3005
R18285 VSS.n2456 VSS.n2455 9.3005
R18286 VSS.n2424 VSS.n2369 9.3005
R18287 VSS.n2424 VSS.n2423 9.3005
R18288 VSS.n2423 VSS.n2422 9.3005
R18289 VSS.n2413 VSS.n2375 9.3005
R18290 VSS.n2375 VSS.n2374 9.3005
R18291 VSS.n2481 VSS.n2480 9.3005
R18292 VSS.n2482 VSS.n2481 9.3005
R18293 VSS.n2483 VSS.n2482 9.3005
R18294 VSS.n2488 VSS.n2487 9.3005
R18295 VSS.n2487 VSS.n2309 9.3005
R18296 VSS.n2389 VSS.n2386 9.3005
R18297 VSS.n3123 VSS.n3122 9.3005
R18298 VSS.n3161 VSS.n3160 9.3005
R18299 VSS.n2851 VSS.n2850 9.3005
R18300 VSS.n3189 VSS.n3188 9.3005
R18301 VSS.n3168 VSS.n3167 9.3005
R18302 VSS.n3169 VSS.n3168 9.3005
R18303 VSS.n3170 VSS.n3169 9.3005
R18304 VSS.n3136 VSS.n3135 9.3005
R18305 VSS.n3136 VSS.n2885 9.3005
R18306 VSS.n2885 VSS.n2884 9.3005
R18307 VSS.n3116 VSS.n3115 9.3005
R18308 VSS.n3117 VSS.n3116 9.3005
R18309 VSS.n3176 VSS.n3175 9.3005
R18310 VSS.n3175 VSS.n2849 9.3005
R18311 VSS.n2849 VSS.n2848 9.3005
R18312 VSS.n3218 VSS.n3217 9.3005
R18313 VSS.n3217 VSS.n3216 9.3005
R18314 VSS.n2911 VSS.n2909 9.3005
R18315 VSS.n3260 VSS.n3259 9.3005
R18316 VSS.n2775 VSS.n2774 9.3005
R18317 VSS.n3310 VSS.n2800 9.3005
R18318 VSS.n2808 VSS.n2806 9.3005
R18319 VSS.n3275 VSS.n3274 9.3005
R18320 VSS.n3347 VSS.n3346 9.3005
R18321 VSS.n3347 VSS.n2780 9.3005
R18322 VSS.n2780 VSS.n2779 9.3005
R18323 VSS.n3329 VSS.n2788 9.3005
R18324 VSS.n3331 VSS.n3330 9.3005
R18325 VSS.n3323 VSS.n3322 9.3005
R18326 VSS.n3324 VSS.n3323 9.3005
R18327 VSS.n3325 VSS.n3324 9.3005
R18328 VSS.n3313 VSS.n3311 9.3005
R18329 VSS.n3291 VSS.n2801 9.3005
R18330 VSS.n2802 VSS.n2801 9.3005
R18331 VSS.n3305 VSS.n2802 9.3005
R18332 VSS.n3250 VSS.n3249 9.3005
R18333 VSS.n3250 VSS.n2823 9.3005
R18334 VSS.n3254 VSS.n2823 9.3005
R18335 VSS.n3261 VSS.n2820 9.3005
R18336 VSS.n3270 VSS.n2814 9.3005
R18337 VSS.n2814 VSS.n2804 9.3005
R18338 VSS.n2804 VSS.n2803 9.3005
R18339 VSS.n3273 VSS.n2813 9.3005
R18340 VSS.n3288 VSS.n3287 9.3005
R18341 VSS.n3356 VSS.n3355 9.3005
R18342 VSS.n3355 VSS.n3354 9.3005
R18343 VSS.n3203 VSS.n2840 9.3005
R18344 VSS.n3211 VSS.n3210 9.3005
R18345 VSS.n3210 VSS.n3209 9.3005
R18346 VSS.n2833 VSS.n2832 9.3005
R18347 VSS.n3202 VSS.n2832 9.3005
R18348 VSS.n3202 VSS.n3201 9.3005
R18349 VSS.n3240 VSS.n2831 9.3005
R18350 VSS.n3242 VSS.n3241 9.3005
R18351 VSS.n3018 VSS.n3017 9.3005
R18352 VSS.n3056 VSS.n3055 9.3005
R18353 VSS.n2926 VSS.n2925 9.3005
R18354 VSS.n3085 VSS.n3084 9.3005
R18355 VSS.n3063 VSS.n3062 9.3005
R18356 VSS.n3064 VSS.n3063 9.3005
R18357 VSS.n3065 VSS.n3064 9.3005
R18358 VSS.n3031 VSS.n3030 9.3005
R18359 VSS.n3031 VSS.n2962 9.3005
R18360 VSS.n2962 VSS.n2961 9.3005
R18361 VSS.n3011 VSS.n3010 9.3005
R18362 VSS.n3012 VSS.n3011 9.3005
R18363 VSS.n3072 VSS.n3071 9.3005
R18364 VSS.n3071 VSS.n2924 9.3005
R18365 VSS.n2924 VSS.n2923 9.3005
R18366 VSS.n3092 VSS.n3091 9.3005
R18367 VSS.n3091 VSS.n3090 9.3005
R18368 VSS.n2986 VSS.n2984 9.3005
R18369 VSS.n9083 VSS.n9082 9.3005
R18370 VSS.n9121 VSS.n9120 9.3005
R18371 VSS.n118 VSS.n117 9.3005
R18372 VSS.n9149 VSS.n9148 9.3005
R18373 VSS.n9128 VSS.n9127 9.3005
R18374 VSS.n9129 VSS.n9128 9.3005
R18375 VSS.n9130 VSS.n9129 9.3005
R18376 VSS.n9096 VSS.n9095 9.3005
R18377 VSS.n9096 VSS.n152 9.3005
R18378 VSS.n152 VSS.n151 9.3005
R18379 VSS.n9076 VSS.n9075 9.3005
R18380 VSS.n9077 VSS.n9076 9.3005
R18381 VSS.n9136 VSS.n9135 9.3005
R18382 VSS.n9135 VSS.n116 9.3005
R18383 VSS.n116 VSS.n115 9.3005
R18384 VSS.n9178 VSS.n9177 9.3005
R18385 VSS.n9177 VSS.n9176 9.3005
R18386 VSS.n190 VSS.n189 9.3005
R18387 VSS.n9220 VSS.n9219 9.3005
R18388 VSS.n42 VSS.n41 9.3005
R18389 VSS.n9270 VSS.n67 9.3005
R18390 VSS.n75 VSS.n73 9.3005
R18391 VSS.n9235 VSS.n9234 9.3005
R18392 VSS.n9307 VSS.n9306 9.3005
R18393 VSS.n9307 VSS.n47 9.3005
R18394 VSS.n47 VSS.n46 9.3005
R18395 VSS.n9289 VSS.n55 9.3005
R18396 VSS.n9291 VSS.n9290 9.3005
R18397 VSS.n9283 VSS.n9282 9.3005
R18398 VSS.n9284 VSS.n9283 9.3005
R18399 VSS.n9285 VSS.n9284 9.3005
R18400 VSS.n9273 VSS.n9271 9.3005
R18401 VSS.n9251 VSS.n68 9.3005
R18402 VSS.n69 VSS.n68 9.3005
R18403 VSS.n9265 VSS.n69 9.3005
R18404 VSS.n9210 VSS.n9209 9.3005
R18405 VSS.n9210 VSS.n90 9.3005
R18406 VSS.n9214 VSS.n90 9.3005
R18407 VSS.n9221 VSS.n87 9.3005
R18408 VSS.n9230 VSS.n81 9.3005
R18409 VSS.n81 VSS.n71 9.3005
R18410 VSS.n71 VSS.n70 9.3005
R18411 VSS.n9233 VSS.n80 9.3005
R18412 VSS.n9248 VSS.n9247 9.3005
R18413 VSS.n9316 VSS.n9315 9.3005
R18414 VSS.n9315 VSS.n9314 9.3005
R18415 VSS.n9163 VSS.n107 9.3005
R18416 VSS.n9171 VSS.n9170 9.3005
R18417 VSS.n9170 VSS.n9169 9.3005
R18418 VSS.n100 VSS.n99 9.3005
R18419 VSS.n9162 VSS.n99 9.3005
R18420 VSS.n9162 VSS.n9161 9.3005
R18421 VSS.n9200 VSS.n98 9.3005
R18422 VSS.n9202 VSS.n9201 9.3005
R18423 VSS.n350 VSS.n349 9.3005
R18424 VSS.n377 VSS.n376 9.3005
R18425 VSS.n390 VSS.n389 9.3005
R18426 VSS.n388 VSS.n309 9.3005
R18427 VSS.n371 VSS.n370 9.3005
R18428 VSS.n370 VSS.n369 9.3005
R18429 VSS.n369 VSS.n368 9.3005
R18430 VSS.n355 VSS.n354 9.3005
R18431 VSS.n356 VSS.n355 9.3005
R18432 VSS.n357 VSS.n356 9.3005
R18433 VSS.n328 VSS.n327 9.3005
R18434 VSS.n344 VSS.n328 9.3005
R18435 VSS.n380 VSS.n379 9.3005
R18436 VSS.n380 VSS.n313 9.3005
R18437 VSS.n384 VSS.n313 9.3005
R18438 VSS.n9052 VSS.n9051 9.3005
R18439 VSS.n9051 VSS.n9050 9.3005
R18440 VSS.n437 VSS.n436 9.3005
R18441 VSS.n8748 VSS.n8747 9.3005
R18442 VSS.n8749 VSS.n8748 9.3005
R18443 VSS.n8750 VSS.n8749 9.3005
R18444 VSS.n8729 VSS.n8695 9.3005
R18445 VSS.n8729 VSS.n8728 9.3005
R18446 VSS.n8728 VSS.n8727 9.3005
R18447 VSS.n8714 VSS.n8698 9.3005
R18448 VSS.n8698 VSS.n8697 9.3005
R18449 VSS.n8754 VSS.n8685 9.3005
R18450 VSS.n8754 VSS.n8680 9.3005
R18451 VSS.n8680 VSS.n8679 9.3005
R18452 VSS.n9004 VSS.n9003 9.3005
R18453 VSS.n9003 VSS.n9002 9.3005
R18454 VSS.n9047 VSS.n9046 9.3005
R18455 VSS.n8886 VSS.n8884 9.3005
R18456 VSS.n8916 VSS.n8884 9.3005
R18457 VSS.n8916 VSS.n8902 9.3005
R18458 VSS.n8911 VSS.n8910 9.3005
R18459 VSS.n8912 VSS.n8911 9.3005
R18460 VSS.n8913 VSS.n8912 9.3005
R18461 VSS.n8870 VSS.n8849 9.3005
R18462 VSS.n8849 VSS.n8823 9.3005
R18463 VSS.n8958 VSS.n8823 9.3005
R18464 VSS.n8806 VSS.n8803 9.3005
R18465 VSS.n8835 VSS.n8806 9.3005
R18466 VSS.n8835 VSS.n8834 9.3005
R18467 VSS.n8842 VSS.n8841 9.3005
R18468 VSS.n8842 VSS.n8822 9.3005
R18469 VSS.n8846 VSS.n8822 9.3005
R18470 VSS.n8925 VSS.n8924 9.3005
R18471 VSS.n8924 VSS.n8923 9.3005
R18472 VSS.n8997 VSS.n8996 9.3005
R18473 VSS.n8996 VSS.n8995 9.3005
R18474 VSS.n8990 VSS.n8989 9.3005
R18475 VSS.n8990 VSS.n8774 9.3005
R18476 VSS.n8774 VSS.n8773 9.3005
R18477 VSS.n566 VSS.n565 9.3005
R18478 VSS.n587 VSS.n586 9.3005
R18479 VSS.n524 VSS.n523 9.3005
R18480 VSS.n608 VSS.n607 9.3005
R18481 VSS.n593 VSS.n592 9.3005
R18482 VSS.n594 VSS.n593 9.3005
R18483 VSS.n595 VSS.n594 9.3005
R18484 VSS.n574 VSS.n537 9.3005
R18485 VSS.n574 VSS.n573 9.3005
R18486 VSS.n573 VSS.n572 9.3005
R18487 VSS.n559 VSS.n540 9.3005
R18488 VSS.n540 VSS.n539 9.3005
R18489 VSS.n599 VSS.n527 9.3005
R18490 VSS.n599 VSS.n522 9.3005
R18491 VSS.n522 VSS.n521 9.3005
R18492 VSS.n822 VSS.n821 9.3005
R18493 VSS.n821 VSS.n820 9.3005
R18494 VSS.n544 VSS.n543 9.3005
R18495 VSS.n9329 VSS.n9328 9.3005
R18496 VSS.n748 VSS.n714 9.3005
R18497 VSS.n767 VSS.n766 9.3005
R18498 VSS.n765 VSS.n699 9.3005
R18499 VSS.n732 VSS.n731 9.3005
R18500 VSS.n689 VSS.n688 9.3005
R18501 VSS.n802 VSS.n801 9.3005
R18502 VSS.n815 VSS.n814 9.3005
R18503 VSS.n814 VSS.n813 9.3005
R18504 VSS.n630 VSS.n629 9.3005
R18505 VSS.n800 VSS.n645 9.3005
R18506 VSS.n808 VSS.n807 9.3005
R18507 VSS.n808 VSS.n619 9.3005
R18508 VSS.n619 VSS.n618 9.3005
R18509 VSS.n793 VSS.n792 9.3005
R18510 VSS.n794 VSS.n793 9.3005
R18511 VSS.n795 VSS.n794 9.3005
R18512 VSS.n787 VSS.n662 9.3005
R18513 VSS.n786 VSS.n785 9.3005
R18514 VSS.n684 VSS.n664 9.3005
R18515 VSS.n665 VSS.n664 9.3005
R18516 VSS.n780 VSS.n665 9.3005
R18517 VSS.n687 VSS.n676 9.3005
R18518 VSS.n671 VSS.n669 9.3005
R18519 VSS.n737 VSS.n736 9.3005
R18520 VSS.n737 VSS.n667 9.3005
R18521 VSS.n667 VSS.n666 9.3005
R18522 VSS.n705 VSS.n701 9.3005
R18523 VSS.n742 VSS.n701 9.3005
R18524 VSS.n743 VSS.n742 9.3005
R18525 VSS.n747 VSS.n706 9.3005
R18526 VSS.n726 VSS.n32 9.3005
R18527 VSS.n32 VSS.n31 9.3005
R18528 VSS.n31 VSS.n30 9.3005
R18529 VSS.n9337 VSS.n9336 9.3005
R18530 VSS.n9336 VSS.n9335 9.3005
R18531 VSS.n909 VSS.n908 9.3005
R18532 VSS.n930 VSS.n929 9.3005
R18533 VSS.n871 VSS.n870 9.3005
R18534 VSS.n952 VSS.n951 9.3005
R18535 VSS.n936 VSS.n935 9.3005
R18536 VSS.n937 VSS.n936 9.3005
R18537 VSS.n938 VSS.n937 9.3005
R18538 VSS.n917 VSS.n885 9.3005
R18539 VSS.n917 VSS.n916 9.3005
R18540 VSS.n916 VSS.n915 9.3005
R18541 VSS.n904 VSS.n888 9.3005
R18542 VSS.n888 VSS.n887 9.3005
R18543 VSS.n943 VSS.n874 9.3005
R18544 VSS.n943 VSS.n869 9.3005
R18545 VSS.n869 VSS.n868 9.3005
R18546 VSS.n959 VSS.n958 9.3005
R18547 VSS.n958 VSS.n957 9.3005
R18548 VSS.n1002 VSS.n1001 9.3005
R18549 VSS.n1117 VSS.n1116 9.3005
R18550 VSS.n1118 VSS.n1117 9.3005
R18551 VSS.n1119 VSS.n1118 9.3005
R18552 VSS.n1098 VSS.n1066 9.3005
R18553 VSS.n1098 VSS.n1097 9.3005
R18554 VSS.n1097 VSS.n1096 9.3005
R18555 VSS.n1085 VSS.n1069 9.3005
R18556 VSS.n1069 VSS.n1068 9.3005
R18557 VSS.n1124 VSS.n1055 9.3005
R18558 VSS.n1124 VSS.n1050 9.3005
R18559 VSS.n1050 VSS.n1049 9.3005
R18560 VSS.n8480 VSS.n8479 9.3005
R18561 VSS.n8479 VSS.n8478 9.3005
R18562 VSS.n8523 VSS.n8522 9.3005
R18563 VSS.n8044 VSS.n8043 9.3005
R18564 VSS.n8043 VSS.n8042 9.3005
R18565 VSS.n8042 VSS.n8041 9.3005
R18566 VSS.n8010 VSS.n7955 9.3005
R18567 VSS.n8010 VSS.n8009 9.3005
R18568 VSS.n8009 VSS.n8008 9.3005
R18569 VSS.n7999 VSS.n7961 9.3005
R18570 VSS.n7961 VSS.n7960 9.3005
R18571 VSS.n8067 VSS.n8066 9.3005
R18572 VSS.n8068 VSS.n8067 9.3005
R18573 VSS.n8069 VSS.n8068 9.3005
R18574 VSS.n8074 VSS.n8073 9.3005
R18575 VSS.n8073 VSS.n7056 9.3005
R18576 VSS.n7975 VSS.n7972 9.3005
R18577 VSS.n7169 VSS.n7168 9.3005
R18578 VSS.n7170 VSS.n7169 9.3005
R18579 VSS.n7171 VSS.n7170 9.3005
R18580 VSS.n7150 VSS.n7116 9.3005
R18581 VSS.n7150 VSS.n7149 9.3005
R18582 VSS.n7149 VSS.n7148 9.3005
R18583 VSS.n7135 VSS.n7119 9.3005
R18584 VSS.n7119 VSS.n7118 9.3005
R18585 VSS.n7175 VSS.n7106 9.3005
R18586 VSS.n7175 VSS.n7101 9.3005
R18587 VSS.n7101 VSS.n7100 9.3005
R18588 VSS.n8431 VSS.n8430 9.3005
R18589 VSS.n8430 VSS.n8429 9.3005
R18590 VSS.n8474 VSS.n8473 9.3005
R18591 VSS.n8395 VSS.n8394 9.3005
R18592 VSS.n8350 VSS.n8349 9.3005
R18593 VSS.n8376 VSS.n8375 9.3005
R18594 VSS.n7247 VSS.n7245 9.3005
R18595 VSS.n7265 VSS.n7264 9.3005
R18596 VSS.n8357 VSS.n7291 9.3005
R18597 VSS.n8357 VSS.n8356 9.3005
R18598 VSS.n8356 VSS.n8355 9.3005
R18599 VSS.n7311 VSS.n7282 9.3005
R18600 VSS.n7292 VSS.n7290 9.3005
R18601 VSS.n7281 VSS.n7277 9.3005
R18602 VSS.n7310 VSS.n7277 9.3005
R18603 VSS.n7310 VSS.n7296 9.3005
R18604 VSS.n8374 VSS.n7275 9.3005
R18605 VSS.n7304 VSS.n7303 9.3005
R18606 VSS.n7304 VSS.n7243 9.3005
R18607 VSS.n7243 VSS.n7242 9.3005
R18608 VSS.n8402 VSS.n8401 9.3005
R18609 VSS.n8403 VSS.n8402 9.3005
R18610 VSS.n8404 VSS.n8403 9.3005
R18611 VSS.n8396 VSS.n7238 9.3005
R18612 VSS.n7260 VSS.n7240 9.3005
R18613 VSS.n7241 VSS.n7240 9.3005
R18614 VSS.n8389 VSS.n7241 9.3005
R18615 VSS.n7263 VSS.n7252 9.3005
R18616 VSS.n7299 VSS.n7298 9.3005
R18617 VSS.n7325 VSS.n7317 9.3005
R18618 VSS.n7317 VSS.n7316 9.3005
R18619 VSS.n7206 VSS.n7205 9.3005
R18620 VSS.n8424 VSS.n8423 9.3005
R18621 VSS.n8423 VSS.n8422 9.3005
R18622 VSS.n8417 VSS.n8416 9.3005
R18623 VSS.n8417 VSS.n7195 9.3005
R18624 VSS.n7195 VSS.n7194 9.3005
R18625 VSS.n8411 VSS.n8410 9.3005
R18626 VSS.n8409 VSS.n7221 9.3005
R18627 VSS.n7534 VSS.n7533 9.15497
R18628 VSS.n7533 VSS.n7532 9.15497
R18629 VSS.n8126 VSS.n8125 9.15497
R18630 VSS.n8125 VSS.n8124 9.15497
R18631 VSS.n8595 VSS.n235 9.15497
R18632 VSS.n235 VSS.n234 9.15497
R18633 VSS.n1373 VSS.n1372 9.15497
R18634 VSS.n1416 VSS.n1373 9.15497
R18635 VSS.n1277 VSS.n1181 9.15497
R18636 VSS.n1181 VSS.n1180 9.15497
R18637 VSS.n1946 VSS.n1945 9.15497
R18638 VSS.n1989 VSS.n1946 9.15497
R18639 VSS.n1850 VSS.n1754 9.15497
R18640 VSS.n1754 VSS.n1753 9.15497
R18641 VSS.n3736 VSS.n3735 9.15497
R18642 VSS.n3735 VSS.n3734 9.15497
R18643 VSS.n3644 VSS.n3548 9.15497
R18644 VSS.n3548 VSS.n3547 9.15497
R18645 VSS.n4328 VSS.n4327 9.15497
R18646 VSS.n4327 VSS.n4326 9.15497
R18647 VSS.n4236 VSS.n4140 9.15497
R18648 VSS.n4140 VSS.n4139 9.15497
R18649 VSS.n4920 VSS.n4919 9.15497
R18650 VSS.n4919 VSS.n4918 9.15497
R18651 VSS.n4828 VSS.n4732 9.15497
R18652 VSS.n4732 VSS.n4731 9.15497
R18653 VSS.n5512 VSS.n5511 9.15497
R18654 VSS.n5511 VSS.n5510 9.15497
R18655 VSS.n5420 VSS.n5324 9.15497
R18656 VSS.n5324 VSS.n5323 9.15497
R18657 VSS.n6104 VSS.n6103 9.15497
R18658 VSS.n6103 VSS.n6102 9.15497
R18659 VSS.n6012 VSS.n5916 9.15497
R18660 VSS.n5916 VSS.n5915 9.15497
R18661 VSS.n6696 VSS.n6695 9.15497
R18662 VSS.n6695 VSS.n6694 9.15497
R18663 VSS.n6604 VSS.n6508 9.15497
R18664 VSS.n6508 VSS.n6507 9.15497
R18665 VSS.n2544 VSS.n2543 9.15497
R18666 VSS.n2587 VSS.n2544 9.15497
R18667 VSS.n2448 VSS.n2352 9.15497
R18668 VSS.n2352 VSS.n2351 9.15497
R18669 VSS.n3144 VSS.n3143 9.15497
R18670 VSS.n3143 VSS.n3142 9.15497
R18671 VSS.n3039 VSS.n3038 9.15497
R18672 VSS.n3038 VSS.n3037 9.15497
R18673 VSS.n9104 VSS.n9103 9.15497
R18674 VSS.n9103 VSS.n9102 9.15497
R18675 VSS.n363 VSS.n321 9.15497
R18676 VSS.n321 VSS.n320 9.15497
R18677 VSS.n8691 VSS.n8690 9.15497
R18678 VSS.n8734 VSS.n8691 9.15497
R18679 VSS.n533 VSS.n532 9.15497
R18680 VSS.n579 VSS.n533 9.15497
R18681 VSS.n881 VSS.n880 9.15497
R18682 VSS.n922 VSS.n881 9.15497
R18683 VSS.n1062 VSS.n1061 9.15497
R18684 VSS.n1103 VSS.n1062 9.15497
R18685 VSS.n8034 VSS.n7938 9.15497
R18686 VSS.n7938 VSS.n7937 9.15497
R18687 VSS.n7112 VSS.n7111 9.15497
R18688 VSS.n7155 VSS.n7112 9.15497
R18689 VSS.n8473 VSS.n7058 8.44336
R18690 VSS.n8430 VSS.n7099 8.44336
R18691 VSS.n7978 VSS.n7972 8.44336
R18692 VSS.n8073 VSS.n8072 8.44336
R18693 VSS.n8522 VSS.n1006 8.44336
R18694 VSS.n8479 VSS.n1048 8.44336
R18695 VSS.n1001 VSS.n439 8.44336
R18696 VSS.n958 VSS.n867 8.44336
R18697 VSS.n7483 VSS.n7478 8.44336
R18698 VSS.n7607 VSS.n7416 8.44336
R18699 VSS.n7897 VSS.n7892 8.44336
R18700 VSS.n8199 VSS.n7830 8.44336
R18701 VSS.n9046 VSS.n194 8.44336
R18702 VSS.n9003 VSS.n8678 8.44336
R18703 VSS.n8539 VSS.n269 8.44336
R18704 VSS.n8634 VSS.n8633 8.44336
R18705 VSS.n1221 VSS.n1215 8.44336
R18706 VSS.n1316 VSS.n1315 8.44336
R18707 VSS.n1709 VSS.n1140 8.44336
R18708 VSS.n1666 VSS.n1360 8.44336
R18709 VSS.n1794 VSS.n1788 8.44336
R18710 VSS.n1889 VSS.n1888 8.44336
R18711 VSS.n2301 VSS.n1713 8.44336
R18712 VSS.n2258 VSS.n1933 8.44336
R18713 VSS.n3588 VSS.n3582 8.44336
R18714 VSS.n3683 VSS.n3682 8.44336
R18715 VSS.n3507 VSS.n3502 8.44336
R18716 VSS.n3809 VSS.n3440 8.44336
R18717 VSS.n4180 VSS.n4174 8.44336
R18718 VSS.n4275 VSS.n4274 8.44336
R18719 VSS.n4099 VSS.n4094 8.44336
R18720 VSS.n4401 VSS.n4032 8.44336
R18721 VSS.n4772 VSS.n4766 8.44336
R18722 VSS.n4867 VSS.n4866 8.44336
R18723 VSS.n4691 VSS.n4686 8.44336
R18724 VSS.n4993 VSS.n4624 8.44336
R18725 VSS.n5364 VSS.n5358 8.44336
R18726 VSS.n5459 VSS.n5458 8.44336
R18727 VSS.n5283 VSS.n5278 8.44336
R18728 VSS.n5585 VSS.n5216 8.44336
R18729 VSS.n5956 VSS.n5950 8.44336
R18730 VSS.n6051 VSS.n6050 8.44336
R18731 VSS.n5875 VSS.n5870 8.44336
R18732 VSS.n6177 VSS.n5808 8.44336
R18733 VSS.n6548 VSS.n6542 8.44336
R18734 VSS.n6643 VSS.n6642 8.44336
R18735 VSS.n6467 VSS.n6462 8.44336
R18736 VSS.n6769 VSS.n6400 8.44336
R18737 VSS.n2392 VSS.n2386 8.44336
R18738 VSS.n2487 VSS.n2486 8.44336
R18739 VSS.n7045 VSS.n2311 8.44336
R18740 VSS.n7002 VSS.n2531 8.44336
R18741 VSS.n2989 VSS.n2984 8.44336
R18742 VSS.n3091 VSS.n2922 8.44336
R18743 VSS.n2914 VSS.n2909 8.44336
R18744 VSS.n3217 VSS.n2847 8.44336
R18745 VSS.n436 VSS.n273 8.44336
R18746 VSS.n9051 VSS.n182 8.44336
R18747 VSS.n189 VSS.n188 8.44336
R18748 VSS.n9177 VSS.n114 8.44336
R18749 VSS.n543 VSS.n542 8.44336
R18750 VSS.n821 VSS.n520 8.44336
R18751 VSS.n7596 VSS.n7590 7.69581
R18752 VSS.n7739 VSS.n7345 7.69581
R18753 VSS.n8188 VSS.n8182 7.69581
R18754 VSS.n8331 VSS.n7759 7.69581
R18755 VSS.n8992 VSS.n8772 7.69581
R18756 VSS.n8919 VSS.n8900 7.69581
R18757 VSS.n1655 VSS.n1454 7.69581
R18758 VSS.n1569 VSS.n7 7.69581
R18759 VSS.n2247 VSS.n2027 7.69581
R18760 VSS.n2180 VSS.n2129 7.69581
R18761 VSS.n3798 VSS.n3792 7.69581
R18762 VSS.n3942 VSS.n3370 7.69581
R18763 VSS.n4390 VSS.n4384 7.69581
R18764 VSS.n4534 VSS.n3962 7.69581
R18765 VSS.n4982 VSS.n4976 7.69581
R18766 VSS.n5126 VSS.n4554 7.69581
R18767 VSS.n5574 VSS.n5568 7.69581
R18768 VSS.n5718 VSS.n5146 7.69581
R18769 VSS.n6166 VSS.n6160 7.69581
R18770 VSS.n6310 VSS.n5738 7.69581
R18771 VSS.n6758 VSS.n6752 7.69581
R18772 VSS.n6902 VSS.n6330 7.69581
R18773 VSS.n6991 VSS.n2625 7.69581
R18774 VSS.n6924 VSS.n2727 7.69581
R18775 VSS.n3206 VSS.n3200 7.69581
R18776 VSS.n3350 VSS.n2777 7.69581
R18777 VSS.n9166 VSS.n9160 7.69581
R18778 VSS.n9310 VSS.n44 7.69581
R18779 VSS.n810 VSS.n617 7.69581
R18780 VSS.n9332 VSS.n29 7.69581
R18781 VSS.n8419 VSS.n7193 7.69581
R18782 VSS.n8352 VSS.n7295 7.69581
R18783 VSS.n8390 VSS.n7224 7.61296
R18784 VSS.n7308 VSS.n7307 7.61296
R18785 VSS.n8069 VSS.t212 7.26922
R18786 VSS.n7646 VSS.n7645 6.39585
R18787 VSS.n7696 VSS.n7360 6.39585
R18788 VSS.n8238 VSS.n8237 6.39585
R18789 VSS.n8288 VSS.n7774 6.39585
R18790 VSS.n1626 VSS.n1485 6.39585
R18791 VSS.n1582 VSS.n1581 6.39585
R18792 VSS.n2218 VSS.n2058 6.39585
R18793 VSS.n2142 VSS.n2141 6.39585
R18794 VSS.n3848 VSS.n3847 6.39585
R18795 VSS.n3898 VSS.n3384 6.39585
R18796 VSS.n4440 VSS.n4439 6.39585
R18797 VSS.n4490 VSS.n3976 6.39585
R18798 VSS.n5032 VSS.n5031 6.39585
R18799 VSS.n5082 VSS.n4568 6.39585
R18800 VSS.n5624 VSS.n5623 6.39585
R18801 VSS.n5674 VSS.n5160 6.39585
R18802 VSS.n6216 VSS.n6215 6.39585
R18803 VSS.n6266 VSS.n5752 6.39585
R18804 VSS.n6808 VSS.n6807 6.39585
R18805 VSS.n6858 VSS.n6344 6.39585
R18806 VSS.n6962 VSS.n2656 6.39585
R18807 VSS.n2740 VSS.n2739 6.39585
R18808 VSS.n3256 VSS.n3255 6.39585
R18809 VSS.n3306 VSS.n2791 6.39585
R18810 VSS.n9216 VSS.n9215 6.39585
R18811 VSS.n9266 VSS.n58 6.39585
R18812 VSS.n8845 VSS.n8824 6.39585
R18813 VSS.n8957 VSS.n8847 6.39585
R18814 VSS.n781 VSS.n648 6.39585
R18815 VSS.n739 VSS.n729 6.39585
R18816 VSS.n8600 VSS.t157 6.21519
R18817 VSS.n1282 VSS.t88 6.21519
R18818 VSS.n1855 VSS.t136 6.21519
R18819 VSS.n3649 VSS.t265 6.21519
R18820 VSS.n4241 VSS.t12 6.21519
R18821 VSS.n4833 VSS.t182 6.21519
R18822 VSS.n5425 VSS.t10 6.21519
R18823 VSS.n6017 VSS.t316 6.21519
R18824 VSS.n6609 VSS.t154 6.21519
R18825 VSS.n2453 VSS.t43 6.21519
R18826 VSS.n3067 VSS.t45 6.21519
R18827 VSS.t270 VSS.n383 6.21519
R18828 VSS.n940 VSS.t131 6.21519
R18829 VSS.n1121 VSS.t180 6.21519
R18830 VSS.n7145 VSS.n7119 5.62907
R18831 VSS.n7173 VSS.n7101 5.62907
R18832 VSS.n8002 VSS.n7961 5.62907
R18833 VSS.n8068 VSS.n7906 5.62907
R18834 VSS.n1093 VSS.n1069 5.62907
R18835 VSS.n1122 VSS.n1050 5.62907
R18836 VSS.n912 VSS.n888 5.62907
R18837 VSS.n941 VSS.n869 5.62907
R18838 VSS.n7506 VSS.n7467 5.62907
R18839 VSS.n7562 VSS.n7418 5.62907
R18840 VSS.n8098 VSS.n7881 5.62907
R18841 VSS.n8154 VSS.n7832 5.62907
R18842 VSS.n8724 VSS.n8698 5.62907
R18843 VSS.n8752 VSS.n8680 5.62907
R18844 VSS.n8563 VSS.n258 5.62907
R18845 VSS.n8629 VSS.n203 5.62907
R18846 VSS.n1245 VSS.n1204 5.62907
R18847 VSS.n1311 VSS.n1149 5.62907
R18848 VSS.n1406 VSS.n1380 5.62907
R18849 VSS.n1434 VSS.n1362 5.62907
R18850 VSS.n1818 VSS.n1777 5.62907
R18851 VSS.n1884 VSS.n1722 5.62907
R18852 VSS.n1979 VSS.n1953 5.62907
R18853 VSS.n2007 VSS.n1935 5.62907
R18854 VSS.n3612 VSS.n3571 5.62907
R18855 VSS.n3678 VSS.n3516 5.62907
R18856 VSS.n3708 VSS.n3491 5.62907
R18857 VSS.n3764 VSS.n3442 5.62907
R18858 VSS.n4204 VSS.n4163 5.62907
R18859 VSS.n4270 VSS.n4108 5.62907
R18860 VSS.n4300 VSS.n4083 5.62907
R18861 VSS.n4356 VSS.n4034 5.62907
R18862 VSS.n4796 VSS.n4755 5.62907
R18863 VSS.n4862 VSS.n4700 5.62907
R18864 VSS.n4892 VSS.n4675 5.62907
R18865 VSS.n4948 VSS.n4626 5.62907
R18866 VSS.n5388 VSS.n5347 5.62907
R18867 VSS.n5454 VSS.n5292 5.62907
R18868 VSS.n5484 VSS.n5267 5.62907
R18869 VSS.n5540 VSS.n5218 5.62907
R18870 VSS.n5980 VSS.n5939 5.62907
R18871 VSS.n6046 VSS.n5884 5.62907
R18872 VSS.n6076 VSS.n5859 5.62907
R18873 VSS.n6132 VSS.n5810 5.62907
R18874 VSS.n6572 VSS.n6531 5.62907
R18875 VSS.n6638 VSS.n6476 5.62907
R18876 VSS.n6668 VSS.n6451 5.62907
R18877 VSS.n6724 VSS.n6402 5.62907
R18878 VSS.n2416 VSS.n2375 5.62907
R18879 VSS.n2482 VSS.n2320 5.62907
R18880 VSS.n2577 VSS.n2551 5.62907
R18881 VSS.n2605 VSS.n2533 5.62907
R18882 VSS.n3011 VSS.n2973 5.62907
R18883 VSS.n3068 VSS.n2924 5.62907
R18884 VSS.n3116 VSS.n2898 5.62907
R18885 VSS.n3172 VSS.n2849 5.62907
R18886 VSS.n346 VSS.n328 5.62907
R18887 VSS.n382 VSS.n313 5.62907
R18888 VSS.n9076 VSS.n165 5.62907
R18889 VSS.n9132 VSS.n116 5.62907
R18890 VSS.n569 VSS.n540 5.62907
R18891 VSS.n597 VSS.n522 5.62907
R18892 VSS.n7346 VSS.n7344 5.33568
R18893 VSS.n7602 VSS.n7585 5.33568
R18894 VSS.n7760 VSS.n7758 5.33568
R18895 VSS.n8194 VSS.n8177 5.33568
R18896 VSS.n8 VSS.n6 5.33568
R18897 VSS.n1661 VSS.n1451 5.33568
R18898 VSS.n2158 VSS.n2157 5.33568
R18899 VSS.n2253 VSS.n2024 5.33568
R18900 VSS.n3371 VSS.n3369 5.33568
R18901 VSS.n3804 VSS.n3787 5.33568
R18902 VSS.n3963 VSS.n3961 5.33568
R18903 VSS.n4396 VSS.n4379 5.33568
R18904 VSS.n4555 VSS.n4553 5.33568
R18905 VSS.n4988 VSS.n4971 5.33568
R18906 VSS.n5147 VSS.n5145 5.33568
R18907 VSS.n5580 VSS.n5563 5.33568
R18908 VSS.n5739 VSS.n5737 5.33568
R18909 VSS.n6172 VSS.n6155 5.33568
R18910 VSS.n6331 VSS.n6329 5.33568
R18911 VSS.n6764 VSS.n6747 5.33568
R18912 VSS.n2756 VSS.n2755 5.33568
R18913 VSS.n6997 VSS.n2622 5.33568
R18914 VSS.n2778 VSS.n2776 5.33568
R18915 VSS.n3212 VSS.n3195 5.33568
R18916 VSS.n45 VSS.n43 5.33568
R18917 VSS.n9172 VSS.n9155 5.33568
R18918 VSS.n8901 VSS.n8899 5.33568
R18919 VSS.n8998 VSS.n8769 5.33568
R18920 VSS.n816 VSS.n614 5.33568
R18921 VSS.n9338 VSS.n26 5.33568
R18922 VSS.n7324 VSS.n7323 5.33568
R18923 VSS.n8425 VSS.n7190 5.33568
R18924 VSS.n8008 VSS.n8007 4.84631
R18925 VSS.n8041 VSS.n8038 4.84631
R18926 VSS.n7152 VSS.n7111 4.84621
R18927 VSS.n7158 VSS.n7111 4.84621
R18928 VSS.n1100 VSS.n1061 4.84621
R18929 VSS.n1106 VSS.n1061 4.84621
R18930 VSS.n7534 VSS.n7449 4.84621
R18931 VSS.n7534 VSS.n7450 4.84621
R18932 VSS.n8034 VSS.n7939 4.84621
R18933 VSS.n8035 VSS.n8034 4.84621
R18934 VSS.n8126 VSS.n7863 4.84621
R18935 VSS.n8126 VSS.n7864 4.84621
R18936 VSS.n8731 VSS.n8690 4.84621
R18937 VSS.n8737 VSS.n8690 4.84621
R18938 VSS.n8595 VSS.n236 4.84621
R18939 VSS.n8596 VSS.n8595 4.84621
R18940 VSS.n1413 VSS.n1372 4.84621
R18941 VSS.n1419 VSS.n1372 4.84621
R18942 VSS.n1277 VSS.n1182 4.84621
R18943 VSS.n1278 VSS.n1277 4.84621
R18944 VSS.n1986 VSS.n1945 4.84621
R18945 VSS.n1992 VSS.n1945 4.84621
R18946 VSS.n1850 VSS.n1755 4.84621
R18947 VSS.n1851 VSS.n1850 4.84621
R18948 VSS.n3736 VSS.n3473 4.84621
R18949 VSS.n3736 VSS.n3474 4.84621
R18950 VSS.n3644 VSS.n3549 4.84621
R18951 VSS.n3645 VSS.n3644 4.84621
R18952 VSS.n4328 VSS.n4065 4.84621
R18953 VSS.n4328 VSS.n4066 4.84621
R18954 VSS.n4236 VSS.n4141 4.84621
R18955 VSS.n4237 VSS.n4236 4.84621
R18956 VSS.n4920 VSS.n4657 4.84621
R18957 VSS.n4920 VSS.n4658 4.84621
R18958 VSS.n4828 VSS.n4733 4.84621
R18959 VSS.n4829 VSS.n4828 4.84621
R18960 VSS.n5512 VSS.n5249 4.84621
R18961 VSS.n5512 VSS.n5250 4.84621
R18962 VSS.n5420 VSS.n5325 4.84621
R18963 VSS.n5421 VSS.n5420 4.84621
R18964 VSS.n6104 VSS.n5841 4.84621
R18965 VSS.n6104 VSS.n5842 4.84621
R18966 VSS.n6012 VSS.n5917 4.84621
R18967 VSS.n6013 VSS.n6012 4.84621
R18968 VSS.n6696 VSS.n6433 4.84621
R18969 VSS.n6696 VSS.n6434 4.84621
R18970 VSS.n6604 VSS.n6509 4.84621
R18971 VSS.n6605 VSS.n6604 4.84621
R18972 VSS.n2584 VSS.n2543 4.84621
R18973 VSS.n2590 VSS.n2543 4.84621
R18974 VSS.n2448 VSS.n2353 4.84621
R18975 VSS.n2449 VSS.n2448 4.84621
R18976 VSS.n3144 VSS.n2880 4.84621
R18977 VSS.n3144 VSS.n2881 4.84621
R18978 VSS.n3039 VSS.n2957 4.84621
R18979 VSS.n3039 VSS.n2958 4.84621
R18980 VSS.n9104 VSS.n147 4.84621
R18981 VSS.n9104 VSS.n148 4.84621
R18982 VSS.n363 VSS.n361 4.84621
R18983 VSS.n364 VSS.n363 4.84621
R18984 VSS.n576 VSS.n532 4.84621
R18985 VSS.n582 VSS.n532 4.84621
R18986 VSS.n919 VSS.n880 4.84621
R18987 VSS.n925 VSS.n880 4.84621
R18988 VSS.n7129 VSS.n7123 4.6505
R18989 VSS.n1079 VSS.n1073 4.6505
R18990 VSS.n7490 VSS.n7469 4.6505
R18991 VSS.n7984 VSS.n7962 4.6505
R18992 VSS.n8082 VSS.n7883 4.6505
R18993 VSS.n8708 VSS.n8702 4.6505
R18994 VSS.n8545 VSS.n259 4.6505
R18995 VSS.n1390 VSS.n1384 4.6505
R18996 VSS.n1227 VSS.n1205 4.6505
R18997 VSS.n1963 VSS.n1957 4.6505
R18998 VSS.n1800 VSS.n1778 4.6505
R18999 VSS.n3692 VSS.n3493 4.6505
R19000 VSS.n3594 VSS.n3572 4.6505
R19001 VSS.n4284 VSS.n4085 4.6505
R19002 VSS.n4186 VSS.n4164 4.6505
R19003 VSS.n4876 VSS.n4677 4.6505
R19004 VSS.n4778 VSS.n4756 4.6505
R19005 VSS.n5468 VSS.n5269 4.6505
R19006 VSS.n5370 VSS.n5348 4.6505
R19007 VSS.n6060 VSS.n5861 4.6505
R19008 VSS.n5962 VSS.n5940 4.6505
R19009 VSS.n6652 VSS.n6453 4.6505
R19010 VSS.n6554 VSS.n6532 4.6505
R19011 VSS.n2561 VSS.n2555 4.6505
R19012 VSS.n2398 VSS.n2376 4.6505
R19013 VSS.n3100 VSS.n2900 4.6505
R19014 VSS.n2995 VSS.n2975 4.6505
R19015 VSS.n9060 VSS.n167 4.6505
R19016 VSS.n340 VSS.n339 4.6505
R19017 VSS.n553 VSS.n549 4.6505
R19018 VSS.n898 VSS.n892 4.6505
R19019 VSS.n7642 VSS.n7395 4.61769
R19020 VSS.n7717 VSS.n7359 4.61769
R19021 VSS.n8234 VSS.n7809 4.61769
R19022 VSS.n8309 VSS.n7773 4.61769
R19023 VSS.n8831 VSS.n8825 4.61769
R19024 VSS.n8915 VSS.n8903 4.61769
R19025 VSS.n1643 VSS.n1484 4.61769
R19026 VSS.n1588 VSS.n1568 4.61769
R19027 VSS.n2235 VSS.n2057 4.61769
R19028 VSS.n2148 VSS.n2128 4.61769
R19029 VSS.n3844 VSS.n3419 4.61769
R19030 VSS.n3919 VSS.n3383 4.61769
R19031 VSS.n4436 VSS.n4011 4.61769
R19032 VSS.n4511 VSS.n3975 4.61769
R19033 VSS.n5028 VSS.n4603 4.61769
R19034 VSS.n5103 VSS.n4567 4.61769
R19035 VSS.n5620 VSS.n5195 4.61769
R19036 VSS.n5695 VSS.n5159 4.61769
R19037 VSS.n6212 VSS.n5787 4.61769
R19038 VSS.n6287 VSS.n5751 4.61769
R19039 VSS.n6804 VSS.n6379 4.61769
R19040 VSS.n6879 VSS.n6343 4.61769
R19041 VSS.n6979 VSS.n2655 4.61769
R19042 VSS.n2746 VSS.n2726 4.61769
R19043 VSS.n3252 VSS.n2826 4.61769
R19044 VSS.n3327 VSS.n2790 4.61769
R19045 VSS.n9212 VSS.n93 4.61769
R19046 VSS.n9287 VSS.n57 4.61769
R19047 VSS.n798 VSS.n647 4.61769
R19048 VSS.n745 VSS.n728 4.61769
R19049 VSS.n8407 VSS.n7223 4.61769
R19050 VSS.n7314 VSS.n7294 4.61769
R19051 VSS.n7179 VSS.n7178 4.5005
R19052 VSS.n7182 VSS.n7181 4.5005
R19053 VSS.n7165 VSS.n7164 4.5005
R19054 VSS.n7140 VSS.n7139 4.5005
R19055 VSS.n7131 VSS.n7130 4.5005
R19056 VSS.n7132 VSS.n7124 4.5005
R19057 VSS.n7128 VSS.n7125 4.5005
R19058 VSS.n7089 VSS.n7087 4.5005
R19059 VSS.n8441 VSS.n8440 4.5005
R19060 VSS.n8448 VSS.n7079 4.5005
R19061 VSS.n8455 VSS.n8454 4.5005
R19062 VSS.n8456 VSS.n7071 4.5005
R19063 VSS.n7136 VSS.n7068 4.5005
R19064 VSS.n8463 VSS.n8462 4.5005
R19065 VSS.n8447 VSS.n8446 4.5005
R19066 VSS.n7180 VSS.n7104 4.5005
R19067 VSS.n8471 VSS.n8470 4.5005
R19068 VSS.n7177 VSS.n7105 4.5005
R19069 VSS.n7177 VSS.n7176 4.5005
R19070 VSS.n7138 VSS.n7137 4.5005
R19071 VSS.n7137 VSS.n7115 4.5005
R19072 VSS.n7134 VSS.n7133 4.5005
R19073 VSS.n7167 VSS.n7166 4.5005
R19074 VSS.n7167 VSS.n7160 4.5005
R19075 VSS.n8433 VSS.n7097 4.5005
R19076 VSS.n8433 VSS.n8432 4.5005
R19077 VSS.n1128 VSS.n1127 4.5005
R19078 VSS.n1131 VSS.n1130 4.5005
R19079 VSS.n1113 VSS.n1112 4.5005
R19080 VSS.n1088 VSS.n1016 4.5005
R19081 VSS.n1081 VSS.n1080 4.5005
R19082 VSS.n1082 VSS.n1074 4.5005
R19083 VSS.n8520 VSS.n8519 4.5005
R19084 VSS.n1078 VSS.n1075 4.5005
R19085 VSS.n1126 VSS.n1054 4.5005
R19086 VSS.n1126 VSS.n1125 4.5005
R19087 VSS.n1038 VSS.n1036 4.5005
R19088 VSS.n8490 VSS.n8489 4.5005
R19089 VSS.n8497 VSS.n1028 4.5005
R19090 VSS.n8504 VSS.n8503 4.5005
R19091 VSS.n1060 VSS.n1024 4.5005
R19092 VSS.n8505 VSS.n1019 4.5005
R19093 VSS.n1087 VSS.n1086 4.5005
R19094 VSS.n1087 VSS.n1065 4.5005
R19095 VSS.n8512 VSS.n8511 4.5005
R19096 VSS.n1084 VSS.n1083 4.5005
R19097 VSS.n8496 VSS.n8495 4.5005
R19098 VSS.n1115 VSS.n1114 4.5005
R19099 VSS.n1115 VSS.n1108 4.5005
R19100 VSS.n1129 VSS.n1053 4.5005
R19101 VSS.n8482 VSS.n1046 4.5005
R19102 VSS.n8482 VSS.n8481 4.5005
R19103 VSS.n7734 VSS.n7733 4.5005
R19104 VSS.n7675 VSS.n7379 4.5005
R19105 VSS.n7638 VSS.n7637 4.5005
R19106 VSS.n7588 VSS.n7586 4.5005
R19107 VSS.n7617 VSS.n7616 4.5005
R19108 VSS.n7628 VSS.n7627 4.5005
R19109 VSS.n7629 VSS.n7628 4.5005
R19110 VSS.n7662 VSS.n7661 4.5005
R19111 VSS.n7635 VSS.n7634 4.5005
R19112 VSS.n7388 VSS.n7387 4.5005
R19113 VSS.n7397 VSS.n7388 4.5005
R19114 VSS.n7728 VSS.n7727 4.5005
R19115 VSS.n7702 VSS.n7368 4.5005
R19116 VSS.n7702 VSS.n7362 4.5005
R19117 VSS.n7709 VSS.n7364 4.5005
R19118 VSS.n7680 VSS.n7676 4.5005
R19119 VSS.n7680 VSS.n7679 4.5005
R19120 VSS.n7683 VSS.n7674 4.5005
R19121 VSS.n7667 VSS.n7666 4.5005
R19122 VSS.n7666 VSS.n7374 4.5005
R19123 VSS.n7732 VSS.n7352 4.5005
R19124 VSS.n7356 VSS.n7350 4.5005
R19125 VSS.n7350 VSS.n7349 4.5005
R19126 VSS.n7690 VSS.n7689 4.5005
R19127 VSS.n7691 VSS.n7690 4.5005
R19128 VSS.n7365 VSS.n7363 4.5005
R19129 VSS.n7747 VSS.n7746 4.5005
R19130 VSS.n7619 VSS.n7618 4.5005
R19131 VSS.n7620 VSS.n7408 4.5005
R19132 VSS.n7427 VSS.n7422 4.5005
R19133 VSS.n7577 VSS.n7576 4.5005
R19134 VSS.n7554 VSS.n7437 4.5005
R19135 VSS.n7465 VSS.n7463 4.5005
R19136 VSS.n7493 VSS.n7491 4.5005
R19137 VSS.n7492 VSS.n7470 4.5005
R19138 VSS.n7495 VSS.n7494 4.5005
R19139 VSS.n7553 VSS.n7552 4.5005
R19140 VSS.n7439 VSS.n7426 4.5005
R19141 VSS.n7543 VSS.n7542 4.5005
R19142 VSS.n7448 VSS.n7446 4.5005
R19143 VSS.n7460 VSS.n7459 4.5005
R19144 VSS.n7515 VSS.n7514 4.5005
R19145 VSS.n7472 VSS.n7462 4.5005
R19146 VSS.n7544 VSS.n7441 4.5005
R19147 VSS.n7575 VSS.n7421 4.5005
R19148 VSS.n7489 VSS.n7488 4.5005
R19149 VSS.n7429 VSS.n7428 4.5005
R19150 VSS.n7564 VSS.n7429 4.5005
R19151 VSS.n7458 VSS.n7456 4.5005
R19152 VSS.n7456 VSS.n7455 4.5005
R19153 VSS.n7504 VSS.n7471 4.5005
R19154 VSS.n7556 VSS.n7555 4.5005
R19155 VSS.n7556 VSS.n7435 4.5005
R19156 VSS.n7611 VSS.n7610 4.5005
R19157 VSS.n7610 VSS.n7609 4.5005
R19158 VSS.n8063 VSS.n7910 4.5005
R19159 VSS.n8062 VSS.n8061 4.5005
R19160 VSS.n7932 VSS.n7931 4.5005
R19161 VSS.n8014 VSS.n8013 4.5005
R19162 VSS.n7987 VSS.n7985 4.5005
R19163 VSS.n7986 VSS.n7963 4.5005
R19164 VSS.n7983 VSS.n7982 4.5005
R19165 VSS.n7989 VSS.n7988 4.5005
R19166 VSS.n8065 VSS.n8064 4.5005
R19167 VSS.n8065 VSS.n7908 4.5005
R19168 VSS.n7921 VSS.n7920 4.5005
R19169 VSS.n8052 VSS.n8051 4.5005
R19170 VSS.n7944 VSS.n7943 4.5005
R19171 VSS.n8023 VSS.n8022 4.5005
R19172 VSS.n8033 VSS.n7941 4.5005
R19173 VSS.n8021 VSS.n8020 4.5005
R19174 VSS.n8012 VSS.n7951 4.5005
R19175 VSS.n8012 VSS.n8011 4.5005
R19176 VSS.n7966 VSS.n7950 4.5005
R19177 VSS.n7998 VSS.n7964 4.5005
R19178 VSS.n7925 VSS.n7923 4.5005
R19179 VSS.n7930 VSS.n7926 4.5005
R19180 VSS.n7928 VSS.n7926 4.5005
R19181 VSS.n8060 VSS.n7912 4.5005
R19182 VSS.n8077 VSS.n8076 4.5005
R19183 VSS.n8076 VSS.n8075 4.5005
R19184 VSS.n8326 VSS.n8325 4.5005
R19185 VSS.n8267 VSS.n7793 4.5005
R19186 VSS.n8230 VSS.n8229 4.5005
R19187 VSS.n8180 VSS.n8178 4.5005
R19188 VSS.n8209 VSS.n8208 4.5005
R19189 VSS.n8220 VSS.n8219 4.5005
R19190 VSS.n8221 VSS.n8220 4.5005
R19191 VSS.n8254 VSS.n8253 4.5005
R19192 VSS.n8227 VSS.n8226 4.5005
R19193 VSS.n7802 VSS.n7801 4.5005
R19194 VSS.n7811 VSS.n7802 4.5005
R19195 VSS.n8320 VSS.n8319 4.5005
R19196 VSS.n8294 VSS.n7782 4.5005
R19197 VSS.n8294 VSS.n7776 4.5005
R19198 VSS.n8301 VSS.n7778 4.5005
R19199 VSS.n8272 VSS.n8268 4.5005
R19200 VSS.n8272 VSS.n8271 4.5005
R19201 VSS.n8275 VSS.n8266 4.5005
R19202 VSS.n8259 VSS.n8258 4.5005
R19203 VSS.n8258 VSS.n7788 4.5005
R19204 VSS.n8324 VSS.n7766 4.5005
R19205 VSS.n7770 VSS.n7764 4.5005
R19206 VSS.n7764 VSS.n7763 4.5005
R19207 VSS.n8282 VSS.n8281 4.5005
R19208 VSS.n8283 VSS.n8282 4.5005
R19209 VSS.n7779 VSS.n7777 4.5005
R19210 VSS.n8339 VSS.n8338 4.5005
R19211 VSS.n8211 VSS.n8210 4.5005
R19212 VSS.n8212 VSS.n7822 4.5005
R19213 VSS.n7841 VSS.n7836 4.5005
R19214 VSS.n8169 VSS.n8168 4.5005
R19215 VSS.n8146 VSS.n7851 4.5005
R19216 VSS.n7879 VSS.n7877 4.5005
R19217 VSS.n8085 VSS.n8083 4.5005
R19218 VSS.n8084 VSS.n7884 4.5005
R19219 VSS.n8087 VSS.n8086 4.5005
R19220 VSS.n8145 VSS.n8144 4.5005
R19221 VSS.n7853 VSS.n7840 4.5005
R19222 VSS.n8135 VSS.n8134 4.5005
R19223 VSS.n7862 VSS.n7860 4.5005
R19224 VSS.n7874 VSS.n7873 4.5005
R19225 VSS.n8107 VSS.n8106 4.5005
R19226 VSS.n7886 VSS.n7876 4.5005
R19227 VSS.n8136 VSS.n7855 4.5005
R19228 VSS.n8167 VSS.n7835 4.5005
R19229 VSS.n8081 VSS.n8080 4.5005
R19230 VSS.n7843 VSS.n7842 4.5005
R19231 VSS.n8156 VSS.n7843 4.5005
R19232 VSS.n7872 VSS.n7870 4.5005
R19233 VSS.n7870 VSS.n7869 4.5005
R19234 VSS.n8096 VSS.n7885 4.5005
R19235 VSS.n8148 VSS.n8147 4.5005
R19236 VSS.n8148 VSS.n7849 4.5005
R19237 VSS.n8203 VSS.n8202 4.5005
R19238 VSS.n8202 VSS.n8201 4.5005
R19239 VSS.n8758 VSS.n8757 4.5005
R19240 VSS.n8761 VSS.n8760 4.5005
R19241 VSS.n8744 VSS.n8743 4.5005
R19242 VSS.n8719 VSS.n8718 4.5005
R19243 VSS.n8710 VSS.n8709 4.5005
R19244 VSS.n8711 VSS.n8703 4.5005
R19245 VSS.n9044 VSS.n9043 4.5005
R19246 VSS.n8707 VSS.n8704 4.5005
R19247 VSS.n8756 VSS.n8684 4.5005
R19248 VSS.n8756 VSS.n8755 4.5005
R19249 VSS.n8668 VSS.n8666 4.5005
R19250 VSS.n9014 VSS.n9013 4.5005
R19251 VSS.n9021 VSS.n8658 4.5005
R19252 VSS.n9028 VSS.n9027 4.5005
R19253 VSS.n9029 VSS.n8650 4.5005
R19254 VSS.n8715 VSS.n8647 4.5005
R19255 VSS.n8717 VSS.n8716 4.5005
R19256 VSS.n8716 VSS.n8694 4.5005
R19257 VSS.n9036 VSS.n9035 4.5005
R19258 VSS.n8713 VSS.n8712 4.5005
R19259 VSS.n9020 VSS.n9019 4.5005
R19260 VSS.n8746 VSS.n8745 4.5005
R19261 VSS.n8746 VSS.n8739 4.5005
R19262 VSS.n8759 VSS.n8683 4.5005
R19263 VSS.n9006 VSS.n8676 4.5005
R19264 VSS.n9006 VSS.n9005 4.5005
R19265 VSS.n8938 VSS.n8937 4.5005
R19266 VSS.n8860 VSS.n8857 4.5005
R19267 VSS.n8977 VSS.n8976 4.5005
R19268 VSS.n8787 VSS.n8770 4.5005
R19269 VSS.n8795 VSS.n8794 4.5005
R19270 VSS.n8988 VSS.n8987 4.5005
R19271 VSS.n8988 VSS.n8776 4.5005
R19272 VSS.n8840 VSS.n8837 4.5005
R19273 VSS.n8980 VSS.n8801 4.5005
R19274 VSS.n8975 VSS.n8804 4.5005
R19275 VSS.n8975 VSS.n8974 4.5005
R19276 VSS.n8896 VSS.n8894 4.5005
R19277 VSS.n8854 VSS.n8852 4.5005
R19278 VSS.n8904 VSS.n8852 4.5005
R19279 VSS.n8881 VSS.n8879 4.5005
R19280 VSS.n8869 VSS.n8858 4.5005
R19281 VSS.n8869 VSS.n8868 4.5005
R19282 VSS.n8874 VSS.n8851 4.5005
R19283 VSS.n8964 VSS.n8963 4.5005
R19284 VSS.n8963 VSS.n8962 4.5005
R19285 VSS.n8936 VSS.n8888 4.5005
R19286 VSS.n8941 VSS.n8940 4.5005
R19287 VSS.n8942 VSS.n8941 4.5005
R19288 VSS.n8864 VSS.n8863 4.5005
R19289 VSS.n8864 VSS.n8821 4.5005
R19290 VSS.n8907 VSS.n8906 4.5005
R19291 VSS.n8927 VSS.n8926 4.5005
R19292 VSS.n8783 VSS.n8777 4.5005
R19293 VSS.n8796 VSS.n8784 4.5005
R19294 VSS.n8624 VSS.n207 4.5005
R19295 VSS.n8623 VSS.n8622 4.5005
R19296 VSS.n229 VSS.n228 4.5005
R19297 VSS.n8575 VSS.n8574 4.5005
R19298 VSS.n8548 VSS.n8546 4.5005
R19299 VSS.n8547 VSS.n260 4.5005
R19300 VSS.n8550 VSS.n8549 4.5005
R19301 VSS.n218 VSS.n217 4.5005
R19302 VSS.n8613 VSS.n8612 4.5005
R19303 VSS.n241 VSS.n240 4.5005
R19304 VSS.n8584 VSS.n8583 4.5005
R19305 VSS.n8582 VSS.n8581 4.5005
R19306 VSS.n263 VSS.n247 4.5005
R19307 VSS.n222 VSS.n220 4.5005
R19308 VSS.n8621 VSS.n209 4.5005
R19309 VSS.n8544 VSS.n8543 4.5005
R19310 VSS.n8626 VSS.n8625 4.5005
R19311 VSS.n8626 VSS.n205 4.5005
R19312 VSS.n8594 VSS.n238 4.5005
R19313 VSS.n8573 VSS.n248 4.5005
R19314 VSS.n8573 VSS.n8572 4.5005
R19315 VSS.n8559 VSS.n261 4.5005
R19316 VSS.n227 VSS.n223 4.5005
R19317 VSS.n225 VSS.n223 4.5005
R19318 VSS.n8638 VSS.n8637 4.5005
R19319 VSS.n8637 VSS.n8636 4.5005
R19320 VSS.n1440 VSS.n1439 4.5005
R19321 VSS.n1443 VSS.n1442 4.5005
R19322 VSS.n1426 VSS.n1425 4.5005
R19323 VSS.n1401 VSS.n1400 4.5005
R19324 VSS.n1392 VSS.n1391 4.5005
R19325 VSS.n1393 VSS.n1385 4.5005
R19326 VSS.n1389 VSS.n1386 4.5005
R19327 VSS.n1350 VSS.n1348 4.5005
R19328 VSS.n1677 VSS.n1676 4.5005
R19329 VSS.n1684 VSS.n1340 4.5005
R19330 VSS.n1691 VSS.n1690 4.5005
R19331 VSS.n1692 VSS.n1332 4.5005
R19332 VSS.n1397 VSS.n1329 4.5005
R19333 VSS.n1699 VSS.n1698 4.5005
R19334 VSS.n1683 VSS.n1682 4.5005
R19335 VSS.n1441 VSS.n1365 4.5005
R19336 VSS.n1707 VSS.n1706 4.5005
R19337 VSS.n1438 VSS.n1366 4.5005
R19338 VSS.n1438 VSS.n1437 4.5005
R19339 VSS.n1399 VSS.n1398 4.5005
R19340 VSS.n1398 VSS.n1376 4.5005
R19341 VSS.n1395 VSS.n1394 4.5005
R19342 VSS.n1428 VSS.n1427 4.5005
R19343 VSS.n1428 VSS.n1421 4.5005
R19344 VSS.n1669 VSS.n1358 4.5005
R19345 VSS.n1669 VSS.n1668 4.5005
R19346 VSS.n1562 VSS.n1552 4.5005
R19347 VSS.n1574 VSS.n1510 4.5005
R19348 VSS.n1636 VSS.n1635 4.5005
R19349 VSS.n1468 VSS.n1452 4.5005
R19350 VSS.n1476 VSS.n1475 4.5005
R19351 VSS.n1650 VSS.n1460 4.5005
R19352 VSS.n1460 VSS.n1458 4.5005
R19353 VSS.n1523 VSS.n1522 4.5005
R19354 VSS.n1494 VSS.n1493 4.5005
R19355 VSS.n1634 VSS.n1489 4.5005
R19356 VSS.n1489 VSS.n1487 4.5005
R19357 VSS.n1557 VSS.n1556 4.5005
R19358 VSS.n1608 VSS.n1607 4.5005
R19359 VSS.n1609 VSS.n1608 4.5005
R19360 VSS.n1603 VSS.n1541 4.5005
R19361 VSS.n1576 VSS.n1575 4.5005
R19362 VSS.n1576 VSS.n1571 4.5005
R19363 VSS.n1613 VSS.n1534 4.5005
R19364 VSS.n1528 VSS.n1527 4.5005
R19365 VSS.n1527 VSS.n1505 4.5005
R19366 VSS.n1561 VSS.n1560 4.5005
R19367 VSS.n1595 VSS.n1550 4.5005
R19368 VSS.n1595 VSS.n1594 4.5005
R19369 VSS.n1620 VSS.n1619 4.5005
R19370 VSS.n1621 VSS.n1620 4.5005
R19371 VSS.n1606 VSS.n1539 4.5005
R19372 VSS.n9347 VSS.n9346 4.5005
R19373 VSS.n1461 VSS.n1459 4.5005
R19374 VSS.n1477 VSS.n1465 4.5005
R19375 VSS.n1306 VSS.n1153 4.5005
R19376 VSS.n1305 VSS.n1304 4.5005
R19377 VSS.n1175 VSS.n1174 4.5005
R19378 VSS.n1257 VSS.n1256 4.5005
R19379 VSS.n1230 VSS.n1228 4.5005
R19380 VSS.n1229 VSS.n1206 4.5005
R19381 VSS.n1232 VSS.n1231 4.5005
R19382 VSS.n1164 VSS.n1163 4.5005
R19383 VSS.n1295 VSS.n1294 4.5005
R19384 VSS.n1187 VSS.n1186 4.5005
R19385 VSS.n1266 VSS.n1265 4.5005
R19386 VSS.n1264 VSS.n1263 4.5005
R19387 VSS.n1209 VSS.n1193 4.5005
R19388 VSS.n1168 VSS.n1166 4.5005
R19389 VSS.n1303 VSS.n1155 4.5005
R19390 VSS.n1226 VSS.n1225 4.5005
R19391 VSS.n1308 VSS.n1307 4.5005
R19392 VSS.n1308 VSS.n1151 4.5005
R19393 VSS.n1276 VSS.n1184 4.5005
R19394 VSS.n1255 VSS.n1194 4.5005
R19395 VSS.n1255 VSS.n1254 4.5005
R19396 VSS.n1241 VSS.n1207 4.5005
R19397 VSS.n1173 VSS.n1169 4.5005
R19398 VSS.n1171 VSS.n1169 4.5005
R19399 VSS.n1320 VSS.n1319 4.5005
R19400 VSS.n1319 VSS.n1318 4.5005
R19401 VSS.n2013 VSS.n2012 4.5005
R19402 VSS.n2016 VSS.n2015 4.5005
R19403 VSS.n1999 VSS.n1998 4.5005
R19404 VSS.n1974 VSS.n1973 4.5005
R19405 VSS.n1965 VSS.n1964 4.5005
R19406 VSS.n1966 VSS.n1958 4.5005
R19407 VSS.n1962 VSS.n1959 4.5005
R19408 VSS.n1923 VSS.n1921 4.5005
R19409 VSS.n2269 VSS.n2268 4.5005
R19410 VSS.n2276 VSS.n1913 4.5005
R19411 VSS.n2283 VSS.n2282 4.5005
R19412 VSS.n2284 VSS.n1905 4.5005
R19413 VSS.n1970 VSS.n1902 4.5005
R19414 VSS.n2291 VSS.n2290 4.5005
R19415 VSS.n2275 VSS.n2274 4.5005
R19416 VSS.n2014 VSS.n1938 4.5005
R19417 VSS.n2299 VSS.n2298 4.5005
R19418 VSS.n2011 VSS.n1939 4.5005
R19419 VSS.n2011 VSS.n2010 4.5005
R19420 VSS.n1972 VSS.n1971 4.5005
R19421 VSS.n1971 VSS.n1949 4.5005
R19422 VSS.n1968 VSS.n1967 4.5005
R19423 VSS.n2001 VSS.n2000 4.5005
R19424 VSS.n2001 VSS.n1994 4.5005
R19425 VSS.n2261 VSS.n1931 4.5005
R19426 VSS.n2261 VSS.n2260 4.5005
R19427 VSS.n2164 VSS.n2163 4.5005
R19428 VSS.n2134 VSS.n2083 4.5005
R19429 VSS.n2228 VSS.n2227 4.5005
R19430 VSS.n2041 VSS.n2025 4.5005
R19431 VSS.n2049 VSS.n2048 4.5005
R19432 VSS.n2242 VSS.n2033 4.5005
R19433 VSS.n2033 VSS.n2031 4.5005
R19434 VSS.n2096 VSS.n2095 4.5005
R19435 VSS.n2067 VSS.n2066 4.5005
R19436 VSS.n2226 VSS.n2062 4.5005
R19437 VSS.n2062 VSS.n2060 4.5005
R19438 VSS.n2169 VSS.n2153 4.5005
R19439 VSS.n2200 VSS.n2199 4.5005
R19440 VSS.n2201 VSS.n2200 4.5005
R19441 VSS.n2195 VSS.n2114 4.5005
R19442 VSS.n2136 VSS.n2135 4.5005
R19443 VSS.n2136 VSS.n2131 4.5005
R19444 VSS.n2205 VSS.n2107 4.5005
R19445 VSS.n2101 VSS.n2100 4.5005
R19446 VSS.n2100 VSS.n2078 4.5005
R19447 VSS.n2165 VSS.n2161 4.5005
R19448 VSS.n2187 VSS.n2123 4.5005
R19449 VSS.n2187 VSS.n2186 4.5005
R19450 VSS.n2212 VSS.n2211 4.5005
R19451 VSS.n2213 VSS.n2212 4.5005
R19452 VSS.n2198 VSS.n2112 4.5005
R19453 VSS.n2154 VSS.n2152 4.5005
R19454 VSS.n2034 VSS.n2032 4.5005
R19455 VSS.n2050 VSS.n2038 4.5005
R19456 VSS.n1879 VSS.n1726 4.5005
R19457 VSS.n1878 VSS.n1877 4.5005
R19458 VSS.n1748 VSS.n1747 4.5005
R19459 VSS.n1830 VSS.n1829 4.5005
R19460 VSS.n1803 VSS.n1801 4.5005
R19461 VSS.n1802 VSS.n1779 4.5005
R19462 VSS.n1805 VSS.n1804 4.5005
R19463 VSS.n1737 VSS.n1736 4.5005
R19464 VSS.n1868 VSS.n1867 4.5005
R19465 VSS.n1760 VSS.n1759 4.5005
R19466 VSS.n1839 VSS.n1838 4.5005
R19467 VSS.n1837 VSS.n1836 4.5005
R19468 VSS.n1782 VSS.n1766 4.5005
R19469 VSS.n1741 VSS.n1739 4.5005
R19470 VSS.n1876 VSS.n1728 4.5005
R19471 VSS.n1799 VSS.n1798 4.5005
R19472 VSS.n1881 VSS.n1880 4.5005
R19473 VSS.n1881 VSS.n1724 4.5005
R19474 VSS.n1849 VSS.n1757 4.5005
R19475 VSS.n1828 VSS.n1767 4.5005
R19476 VSS.n1828 VSS.n1827 4.5005
R19477 VSS.n1814 VSS.n1780 4.5005
R19478 VSS.n1746 VSS.n1742 4.5005
R19479 VSS.n1744 VSS.n1742 4.5005
R19480 VSS.n1893 VSS.n1892 4.5005
R19481 VSS.n1892 VSS.n1891 4.5005
R19482 VSS.n3451 VSS.n3446 4.5005
R19483 VSS.n3779 VSS.n3778 4.5005
R19484 VSS.n3756 VSS.n3461 4.5005
R19485 VSS.n3489 VSS.n3487 4.5005
R19486 VSS.n3695 VSS.n3693 4.5005
R19487 VSS.n3694 VSS.n3494 4.5005
R19488 VSS.n3697 VSS.n3696 4.5005
R19489 VSS.n3755 VSS.n3754 4.5005
R19490 VSS.n3463 VSS.n3450 4.5005
R19491 VSS.n3745 VSS.n3744 4.5005
R19492 VSS.n3472 VSS.n3470 4.5005
R19493 VSS.n3484 VSS.n3483 4.5005
R19494 VSS.n3717 VSS.n3716 4.5005
R19495 VSS.n3496 VSS.n3486 4.5005
R19496 VSS.n3746 VSS.n3465 4.5005
R19497 VSS.n3777 VSS.n3445 4.5005
R19498 VSS.n3691 VSS.n3690 4.5005
R19499 VSS.n3453 VSS.n3452 4.5005
R19500 VSS.n3766 VSS.n3453 4.5005
R19501 VSS.n3482 VSS.n3480 4.5005
R19502 VSS.n3480 VSS.n3479 4.5005
R19503 VSS.n3706 VSS.n3495 4.5005
R19504 VSS.n3758 VSS.n3757 4.5005
R19505 VSS.n3758 VSS.n3459 4.5005
R19506 VSS.n3813 VSS.n3812 4.5005
R19507 VSS.n3812 VSS.n3811 4.5005
R19508 VSS.n3936 VSS.n3376 4.5005
R19509 VSS.n3877 VSS.n3403 4.5005
R19510 VSS.n3840 VSS.n3839 4.5005
R19511 VSS.n3790 VSS.n3788 4.5005
R19512 VSS.n3819 VSS.n3818 4.5005
R19513 VSS.n3830 VSS.n3829 4.5005
R19514 VSS.n3831 VSS.n3830 4.5005
R19515 VSS.n3864 VSS.n3863 4.5005
R19516 VSS.n3837 VSS.n3836 4.5005
R19517 VSS.n3412 VSS.n3411 4.5005
R19518 VSS.n3421 VSS.n3412 4.5005
R19519 VSS.n3931 VSS.n3930 4.5005
R19520 VSS.n3904 VSS.n3392 4.5005
R19521 VSS.n3904 VSS.n3386 4.5005
R19522 VSS.n3911 VSS.n3388 4.5005
R19523 VSS.n3882 VSS.n3878 4.5005
R19524 VSS.n3882 VSS.n3881 4.5005
R19525 VSS.n3885 VSS.n3876 4.5005
R19526 VSS.n3869 VSS.n3868 4.5005
R19527 VSS.n3868 VSS.n3398 4.5005
R19528 VSS.n3935 VSS.n3934 4.5005
R19529 VSS.n3377 VSS.n3375 4.5005
R19530 VSS.n3375 VSS.n3374 4.5005
R19531 VSS.n3892 VSS.n3891 4.5005
R19532 VSS.n3893 VSS.n3892 4.5005
R19533 VSS.n3389 VSS.n3387 4.5005
R19534 VSS.n3950 VSS.n3949 4.5005
R19535 VSS.n3821 VSS.n3820 4.5005
R19536 VSS.n3822 VSS.n3432 4.5005
R19537 VSS.n3673 VSS.n3520 4.5005
R19538 VSS.n3672 VSS.n3671 4.5005
R19539 VSS.n3542 VSS.n3541 4.5005
R19540 VSS.n3624 VSS.n3623 4.5005
R19541 VSS.n3597 VSS.n3595 4.5005
R19542 VSS.n3596 VSS.n3573 4.5005
R19543 VSS.n3599 VSS.n3598 4.5005
R19544 VSS.n3531 VSS.n3530 4.5005
R19545 VSS.n3662 VSS.n3661 4.5005
R19546 VSS.n3554 VSS.n3553 4.5005
R19547 VSS.n3633 VSS.n3632 4.5005
R19548 VSS.n3631 VSS.n3630 4.5005
R19549 VSS.n3576 VSS.n3560 4.5005
R19550 VSS.n3535 VSS.n3533 4.5005
R19551 VSS.n3670 VSS.n3522 4.5005
R19552 VSS.n3593 VSS.n3592 4.5005
R19553 VSS.n3675 VSS.n3674 4.5005
R19554 VSS.n3675 VSS.n3518 4.5005
R19555 VSS.n3643 VSS.n3551 4.5005
R19556 VSS.n3622 VSS.n3561 4.5005
R19557 VSS.n3622 VSS.n3621 4.5005
R19558 VSS.n3608 VSS.n3574 4.5005
R19559 VSS.n3540 VSS.n3536 4.5005
R19560 VSS.n3538 VSS.n3536 4.5005
R19561 VSS.n3687 VSS.n3686 4.5005
R19562 VSS.n3686 VSS.n3685 4.5005
R19563 VSS.n4043 VSS.n4038 4.5005
R19564 VSS.n4371 VSS.n4370 4.5005
R19565 VSS.n4348 VSS.n4053 4.5005
R19566 VSS.n4081 VSS.n4079 4.5005
R19567 VSS.n4287 VSS.n4285 4.5005
R19568 VSS.n4286 VSS.n4086 4.5005
R19569 VSS.n4289 VSS.n4288 4.5005
R19570 VSS.n4347 VSS.n4346 4.5005
R19571 VSS.n4055 VSS.n4042 4.5005
R19572 VSS.n4337 VSS.n4336 4.5005
R19573 VSS.n4064 VSS.n4062 4.5005
R19574 VSS.n4076 VSS.n4075 4.5005
R19575 VSS.n4309 VSS.n4308 4.5005
R19576 VSS.n4088 VSS.n4078 4.5005
R19577 VSS.n4338 VSS.n4057 4.5005
R19578 VSS.n4369 VSS.n4037 4.5005
R19579 VSS.n4283 VSS.n4282 4.5005
R19580 VSS.n4045 VSS.n4044 4.5005
R19581 VSS.n4358 VSS.n4045 4.5005
R19582 VSS.n4074 VSS.n4072 4.5005
R19583 VSS.n4072 VSS.n4071 4.5005
R19584 VSS.n4298 VSS.n4087 4.5005
R19585 VSS.n4350 VSS.n4349 4.5005
R19586 VSS.n4350 VSS.n4051 4.5005
R19587 VSS.n4405 VSS.n4404 4.5005
R19588 VSS.n4404 VSS.n4403 4.5005
R19589 VSS.n4528 VSS.n3968 4.5005
R19590 VSS.n4469 VSS.n3995 4.5005
R19591 VSS.n4432 VSS.n4431 4.5005
R19592 VSS.n4382 VSS.n4380 4.5005
R19593 VSS.n4411 VSS.n4410 4.5005
R19594 VSS.n4422 VSS.n4421 4.5005
R19595 VSS.n4423 VSS.n4422 4.5005
R19596 VSS.n4456 VSS.n4455 4.5005
R19597 VSS.n4429 VSS.n4428 4.5005
R19598 VSS.n4004 VSS.n4003 4.5005
R19599 VSS.n4013 VSS.n4004 4.5005
R19600 VSS.n4523 VSS.n4522 4.5005
R19601 VSS.n4496 VSS.n3984 4.5005
R19602 VSS.n4496 VSS.n3978 4.5005
R19603 VSS.n4503 VSS.n3980 4.5005
R19604 VSS.n4474 VSS.n4470 4.5005
R19605 VSS.n4474 VSS.n4473 4.5005
R19606 VSS.n4477 VSS.n4468 4.5005
R19607 VSS.n4461 VSS.n4460 4.5005
R19608 VSS.n4460 VSS.n3990 4.5005
R19609 VSS.n4527 VSS.n4526 4.5005
R19610 VSS.n3969 VSS.n3967 4.5005
R19611 VSS.n3967 VSS.n3966 4.5005
R19612 VSS.n4484 VSS.n4483 4.5005
R19613 VSS.n4485 VSS.n4484 4.5005
R19614 VSS.n3981 VSS.n3979 4.5005
R19615 VSS.n4542 VSS.n4541 4.5005
R19616 VSS.n4413 VSS.n4412 4.5005
R19617 VSS.n4414 VSS.n4024 4.5005
R19618 VSS.n4265 VSS.n4112 4.5005
R19619 VSS.n4264 VSS.n4263 4.5005
R19620 VSS.n4134 VSS.n4133 4.5005
R19621 VSS.n4216 VSS.n4215 4.5005
R19622 VSS.n4189 VSS.n4187 4.5005
R19623 VSS.n4188 VSS.n4165 4.5005
R19624 VSS.n4191 VSS.n4190 4.5005
R19625 VSS.n4123 VSS.n4122 4.5005
R19626 VSS.n4254 VSS.n4253 4.5005
R19627 VSS.n4146 VSS.n4145 4.5005
R19628 VSS.n4225 VSS.n4224 4.5005
R19629 VSS.n4223 VSS.n4222 4.5005
R19630 VSS.n4168 VSS.n4152 4.5005
R19631 VSS.n4127 VSS.n4125 4.5005
R19632 VSS.n4262 VSS.n4114 4.5005
R19633 VSS.n4185 VSS.n4184 4.5005
R19634 VSS.n4267 VSS.n4266 4.5005
R19635 VSS.n4267 VSS.n4110 4.5005
R19636 VSS.n4235 VSS.n4143 4.5005
R19637 VSS.n4214 VSS.n4153 4.5005
R19638 VSS.n4214 VSS.n4213 4.5005
R19639 VSS.n4200 VSS.n4166 4.5005
R19640 VSS.n4132 VSS.n4128 4.5005
R19641 VSS.n4130 VSS.n4128 4.5005
R19642 VSS.n4279 VSS.n4278 4.5005
R19643 VSS.n4278 VSS.n4277 4.5005
R19644 VSS.n4635 VSS.n4630 4.5005
R19645 VSS.n4963 VSS.n4962 4.5005
R19646 VSS.n4940 VSS.n4645 4.5005
R19647 VSS.n4673 VSS.n4671 4.5005
R19648 VSS.n4879 VSS.n4877 4.5005
R19649 VSS.n4878 VSS.n4678 4.5005
R19650 VSS.n4881 VSS.n4880 4.5005
R19651 VSS.n4939 VSS.n4938 4.5005
R19652 VSS.n4647 VSS.n4634 4.5005
R19653 VSS.n4929 VSS.n4928 4.5005
R19654 VSS.n4656 VSS.n4654 4.5005
R19655 VSS.n4668 VSS.n4667 4.5005
R19656 VSS.n4901 VSS.n4900 4.5005
R19657 VSS.n4680 VSS.n4670 4.5005
R19658 VSS.n4930 VSS.n4649 4.5005
R19659 VSS.n4961 VSS.n4629 4.5005
R19660 VSS.n4875 VSS.n4874 4.5005
R19661 VSS.n4637 VSS.n4636 4.5005
R19662 VSS.n4950 VSS.n4637 4.5005
R19663 VSS.n4666 VSS.n4664 4.5005
R19664 VSS.n4664 VSS.n4663 4.5005
R19665 VSS.n4890 VSS.n4679 4.5005
R19666 VSS.n4942 VSS.n4941 4.5005
R19667 VSS.n4942 VSS.n4643 4.5005
R19668 VSS.n4997 VSS.n4996 4.5005
R19669 VSS.n4996 VSS.n4995 4.5005
R19670 VSS.n5120 VSS.n4560 4.5005
R19671 VSS.n5061 VSS.n4587 4.5005
R19672 VSS.n5024 VSS.n5023 4.5005
R19673 VSS.n4974 VSS.n4972 4.5005
R19674 VSS.n5003 VSS.n5002 4.5005
R19675 VSS.n5014 VSS.n5013 4.5005
R19676 VSS.n5015 VSS.n5014 4.5005
R19677 VSS.n5048 VSS.n5047 4.5005
R19678 VSS.n5021 VSS.n5020 4.5005
R19679 VSS.n4596 VSS.n4595 4.5005
R19680 VSS.n4605 VSS.n4596 4.5005
R19681 VSS.n5115 VSS.n5114 4.5005
R19682 VSS.n5088 VSS.n4576 4.5005
R19683 VSS.n5088 VSS.n4570 4.5005
R19684 VSS.n5095 VSS.n4572 4.5005
R19685 VSS.n5066 VSS.n5062 4.5005
R19686 VSS.n5066 VSS.n5065 4.5005
R19687 VSS.n5069 VSS.n5060 4.5005
R19688 VSS.n5053 VSS.n5052 4.5005
R19689 VSS.n5052 VSS.n4582 4.5005
R19690 VSS.n5119 VSS.n5118 4.5005
R19691 VSS.n4561 VSS.n4559 4.5005
R19692 VSS.n4559 VSS.n4558 4.5005
R19693 VSS.n5076 VSS.n5075 4.5005
R19694 VSS.n5077 VSS.n5076 4.5005
R19695 VSS.n4573 VSS.n4571 4.5005
R19696 VSS.n5134 VSS.n5133 4.5005
R19697 VSS.n5005 VSS.n5004 4.5005
R19698 VSS.n5006 VSS.n4616 4.5005
R19699 VSS.n4857 VSS.n4704 4.5005
R19700 VSS.n4856 VSS.n4855 4.5005
R19701 VSS.n4726 VSS.n4725 4.5005
R19702 VSS.n4808 VSS.n4807 4.5005
R19703 VSS.n4781 VSS.n4779 4.5005
R19704 VSS.n4780 VSS.n4757 4.5005
R19705 VSS.n4783 VSS.n4782 4.5005
R19706 VSS.n4715 VSS.n4714 4.5005
R19707 VSS.n4846 VSS.n4845 4.5005
R19708 VSS.n4738 VSS.n4737 4.5005
R19709 VSS.n4817 VSS.n4816 4.5005
R19710 VSS.n4815 VSS.n4814 4.5005
R19711 VSS.n4760 VSS.n4744 4.5005
R19712 VSS.n4719 VSS.n4717 4.5005
R19713 VSS.n4854 VSS.n4706 4.5005
R19714 VSS.n4777 VSS.n4776 4.5005
R19715 VSS.n4859 VSS.n4858 4.5005
R19716 VSS.n4859 VSS.n4702 4.5005
R19717 VSS.n4827 VSS.n4735 4.5005
R19718 VSS.n4806 VSS.n4745 4.5005
R19719 VSS.n4806 VSS.n4805 4.5005
R19720 VSS.n4792 VSS.n4758 4.5005
R19721 VSS.n4724 VSS.n4720 4.5005
R19722 VSS.n4722 VSS.n4720 4.5005
R19723 VSS.n4871 VSS.n4870 4.5005
R19724 VSS.n4870 VSS.n4869 4.5005
R19725 VSS.n5227 VSS.n5222 4.5005
R19726 VSS.n5555 VSS.n5554 4.5005
R19727 VSS.n5532 VSS.n5237 4.5005
R19728 VSS.n5265 VSS.n5263 4.5005
R19729 VSS.n5471 VSS.n5469 4.5005
R19730 VSS.n5470 VSS.n5270 4.5005
R19731 VSS.n5473 VSS.n5472 4.5005
R19732 VSS.n5531 VSS.n5530 4.5005
R19733 VSS.n5239 VSS.n5226 4.5005
R19734 VSS.n5521 VSS.n5520 4.5005
R19735 VSS.n5248 VSS.n5246 4.5005
R19736 VSS.n5260 VSS.n5259 4.5005
R19737 VSS.n5493 VSS.n5492 4.5005
R19738 VSS.n5272 VSS.n5262 4.5005
R19739 VSS.n5522 VSS.n5241 4.5005
R19740 VSS.n5553 VSS.n5221 4.5005
R19741 VSS.n5467 VSS.n5466 4.5005
R19742 VSS.n5229 VSS.n5228 4.5005
R19743 VSS.n5542 VSS.n5229 4.5005
R19744 VSS.n5258 VSS.n5256 4.5005
R19745 VSS.n5256 VSS.n5255 4.5005
R19746 VSS.n5482 VSS.n5271 4.5005
R19747 VSS.n5534 VSS.n5533 4.5005
R19748 VSS.n5534 VSS.n5235 4.5005
R19749 VSS.n5589 VSS.n5588 4.5005
R19750 VSS.n5588 VSS.n5587 4.5005
R19751 VSS.n5712 VSS.n5152 4.5005
R19752 VSS.n5653 VSS.n5179 4.5005
R19753 VSS.n5616 VSS.n5615 4.5005
R19754 VSS.n5566 VSS.n5564 4.5005
R19755 VSS.n5595 VSS.n5594 4.5005
R19756 VSS.n5606 VSS.n5605 4.5005
R19757 VSS.n5607 VSS.n5606 4.5005
R19758 VSS.n5640 VSS.n5639 4.5005
R19759 VSS.n5613 VSS.n5612 4.5005
R19760 VSS.n5188 VSS.n5187 4.5005
R19761 VSS.n5197 VSS.n5188 4.5005
R19762 VSS.n5707 VSS.n5706 4.5005
R19763 VSS.n5680 VSS.n5168 4.5005
R19764 VSS.n5680 VSS.n5162 4.5005
R19765 VSS.n5687 VSS.n5164 4.5005
R19766 VSS.n5658 VSS.n5654 4.5005
R19767 VSS.n5658 VSS.n5657 4.5005
R19768 VSS.n5661 VSS.n5652 4.5005
R19769 VSS.n5645 VSS.n5644 4.5005
R19770 VSS.n5644 VSS.n5174 4.5005
R19771 VSS.n5711 VSS.n5710 4.5005
R19772 VSS.n5153 VSS.n5151 4.5005
R19773 VSS.n5151 VSS.n5150 4.5005
R19774 VSS.n5668 VSS.n5667 4.5005
R19775 VSS.n5669 VSS.n5668 4.5005
R19776 VSS.n5165 VSS.n5163 4.5005
R19777 VSS.n5726 VSS.n5725 4.5005
R19778 VSS.n5597 VSS.n5596 4.5005
R19779 VSS.n5598 VSS.n5208 4.5005
R19780 VSS.n5449 VSS.n5296 4.5005
R19781 VSS.n5448 VSS.n5447 4.5005
R19782 VSS.n5318 VSS.n5317 4.5005
R19783 VSS.n5400 VSS.n5399 4.5005
R19784 VSS.n5373 VSS.n5371 4.5005
R19785 VSS.n5372 VSS.n5349 4.5005
R19786 VSS.n5375 VSS.n5374 4.5005
R19787 VSS.n5307 VSS.n5306 4.5005
R19788 VSS.n5438 VSS.n5437 4.5005
R19789 VSS.n5330 VSS.n5329 4.5005
R19790 VSS.n5409 VSS.n5408 4.5005
R19791 VSS.n5407 VSS.n5406 4.5005
R19792 VSS.n5352 VSS.n5336 4.5005
R19793 VSS.n5311 VSS.n5309 4.5005
R19794 VSS.n5446 VSS.n5298 4.5005
R19795 VSS.n5369 VSS.n5368 4.5005
R19796 VSS.n5451 VSS.n5450 4.5005
R19797 VSS.n5451 VSS.n5294 4.5005
R19798 VSS.n5419 VSS.n5327 4.5005
R19799 VSS.n5398 VSS.n5337 4.5005
R19800 VSS.n5398 VSS.n5397 4.5005
R19801 VSS.n5384 VSS.n5350 4.5005
R19802 VSS.n5316 VSS.n5312 4.5005
R19803 VSS.n5314 VSS.n5312 4.5005
R19804 VSS.n5463 VSS.n5462 4.5005
R19805 VSS.n5462 VSS.n5461 4.5005
R19806 VSS.n5819 VSS.n5814 4.5005
R19807 VSS.n6147 VSS.n6146 4.5005
R19808 VSS.n6124 VSS.n5829 4.5005
R19809 VSS.n5857 VSS.n5855 4.5005
R19810 VSS.n6063 VSS.n6061 4.5005
R19811 VSS.n6062 VSS.n5862 4.5005
R19812 VSS.n6065 VSS.n6064 4.5005
R19813 VSS.n6123 VSS.n6122 4.5005
R19814 VSS.n5831 VSS.n5818 4.5005
R19815 VSS.n6113 VSS.n6112 4.5005
R19816 VSS.n5840 VSS.n5838 4.5005
R19817 VSS.n5852 VSS.n5851 4.5005
R19818 VSS.n6085 VSS.n6084 4.5005
R19819 VSS.n5864 VSS.n5854 4.5005
R19820 VSS.n6114 VSS.n5833 4.5005
R19821 VSS.n6145 VSS.n5813 4.5005
R19822 VSS.n6059 VSS.n6058 4.5005
R19823 VSS.n5821 VSS.n5820 4.5005
R19824 VSS.n6134 VSS.n5821 4.5005
R19825 VSS.n5850 VSS.n5848 4.5005
R19826 VSS.n5848 VSS.n5847 4.5005
R19827 VSS.n6074 VSS.n5863 4.5005
R19828 VSS.n6126 VSS.n6125 4.5005
R19829 VSS.n6126 VSS.n5827 4.5005
R19830 VSS.n6181 VSS.n6180 4.5005
R19831 VSS.n6180 VSS.n6179 4.5005
R19832 VSS.n6304 VSS.n5744 4.5005
R19833 VSS.n6245 VSS.n5771 4.5005
R19834 VSS.n6208 VSS.n6207 4.5005
R19835 VSS.n6158 VSS.n6156 4.5005
R19836 VSS.n6187 VSS.n6186 4.5005
R19837 VSS.n6198 VSS.n6197 4.5005
R19838 VSS.n6199 VSS.n6198 4.5005
R19839 VSS.n6232 VSS.n6231 4.5005
R19840 VSS.n6205 VSS.n6204 4.5005
R19841 VSS.n5780 VSS.n5779 4.5005
R19842 VSS.n5789 VSS.n5780 4.5005
R19843 VSS.n6299 VSS.n6298 4.5005
R19844 VSS.n6272 VSS.n5760 4.5005
R19845 VSS.n6272 VSS.n5754 4.5005
R19846 VSS.n6279 VSS.n5756 4.5005
R19847 VSS.n6250 VSS.n6246 4.5005
R19848 VSS.n6250 VSS.n6249 4.5005
R19849 VSS.n6253 VSS.n6244 4.5005
R19850 VSS.n6237 VSS.n6236 4.5005
R19851 VSS.n6236 VSS.n5766 4.5005
R19852 VSS.n6303 VSS.n6302 4.5005
R19853 VSS.n5745 VSS.n5743 4.5005
R19854 VSS.n5743 VSS.n5742 4.5005
R19855 VSS.n6260 VSS.n6259 4.5005
R19856 VSS.n6261 VSS.n6260 4.5005
R19857 VSS.n5757 VSS.n5755 4.5005
R19858 VSS.n6318 VSS.n6317 4.5005
R19859 VSS.n6189 VSS.n6188 4.5005
R19860 VSS.n6190 VSS.n5800 4.5005
R19861 VSS.n6041 VSS.n5888 4.5005
R19862 VSS.n6040 VSS.n6039 4.5005
R19863 VSS.n5910 VSS.n5909 4.5005
R19864 VSS.n5992 VSS.n5991 4.5005
R19865 VSS.n5965 VSS.n5963 4.5005
R19866 VSS.n5964 VSS.n5941 4.5005
R19867 VSS.n5967 VSS.n5966 4.5005
R19868 VSS.n5899 VSS.n5898 4.5005
R19869 VSS.n6030 VSS.n6029 4.5005
R19870 VSS.n5922 VSS.n5921 4.5005
R19871 VSS.n6001 VSS.n6000 4.5005
R19872 VSS.n5999 VSS.n5998 4.5005
R19873 VSS.n5944 VSS.n5928 4.5005
R19874 VSS.n5903 VSS.n5901 4.5005
R19875 VSS.n6038 VSS.n5890 4.5005
R19876 VSS.n5961 VSS.n5960 4.5005
R19877 VSS.n6043 VSS.n6042 4.5005
R19878 VSS.n6043 VSS.n5886 4.5005
R19879 VSS.n6011 VSS.n5919 4.5005
R19880 VSS.n5990 VSS.n5929 4.5005
R19881 VSS.n5990 VSS.n5989 4.5005
R19882 VSS.n5976 VSS.n5942 4.5005
R19883 VSS.n5908 VSS.n5904 4.5005
R19884 VSS.n5906 VSS.n5904 4.5005
R19885 VSS.n6055 VSS.n6054 4.5005
R19886 VSS.n6054 VSS.n6053 4.5005
R19887 VSS.n6411 VSS.n6406 4.5005
R19888 VSS.n6739 VSS.n6738 4.5005
R19889 VSS.n6716 VSS.n6421 4.5005
R19890 VSS.n6449 VSS.n6447 4.5005
R19891 VSS.n6655 VSS.n6653 4.5005
R19892 VSS.n6654 VSS.n6454 4.5005
R19893 VSS.n6657 VSS.n6656 4.5005
R19894 VSS.n6715 VSS.n6714 4.5005
R19895 VSS.n6423 VSS.n6410 4.5005
R19896 VSS.n6705 VSS.n6704 4.5005
R19897 VSS.n6432 VSS.n6430 4.5005
R19898 VSS.n6444 VSS.n6443 4.5005
R19899 VSS.n6677 VSS.n6676 4.5005
R19900 VSS.n6456 VSS.n6446 4.5005
R19901 VSS.n6706 VSS.n6425 4.5005
R19902 VSS.n6737 VSS.n6405 4.5005
R19903 VSS.n6651 VSS.n6650 4.5005
R19904 VSS.n6413 VSS.n6412 4.5005
R19905 VSS.n6726 VSS.n6413 4.5005
R19906 VSS.n6442 VSS.n6440 4.5005
R19907 VSS.n6440 VSS.n6439 4.5005
R19908 VSS.n6666 VSS.n6455 4.5005
R19909 VSS.n6718 VSS.n6717 4.5005
R19910 VSS.n6718 VSS.n6419 4.5005
R19911 VSS.n6773 VSS.n6772 4.5005
R19912 VSS.n6772 VSS.n6771 4.5005
R19913 VSS.n6896 VSS.n6336 4.5005
R19914 VSS.n6837 VSS.n6363 4.5005
R19915 VSS.n6800 VSS.n6799 4.5005
R19916 VSS.n6750 VSS.n6748 4.5005
R19917 VSS.n6779 VSS.n6778 4.5005
R19918 VSS.n6790 VSS.n6789 4.5005
R19919 VSS.n6791 VSS.n6790 4.5005
R19920 VSS.n6824 VSS.n6823 4.5005
R19921 VSS.n6797 VSS.n6796 4.5005
R19922 VSS.n6372 VSS.n6371 4.5005
R19923 VSS.n6381 VSS.n6372 4.5005
R19924 VSS.n6891 VSS.n6890 4.5005
R19925 VSS.n6864 VSS.n6352 4.5005
R19926 VSS.n6864 VSS.n6346 4.5005
R19927 VSS.n6871 VSS.n6348 4.5005
R19928 VSS.n6842 VSS.n6838 4.5005
R19929 VSS.n6842 VSS.n6841 4.5005
R19930 VSS.n6845 VSS.n6836 4.5005
R19931 VSS.n6829 VSS.n6828 4.5005
R19932 VSS.n6828 VSS.n6358 4.5005
R19933 VSS.n6895 VSS.n6894 4.5005
R19934 VSS.n6337 VSS.n6335 4.5005
R19935 VSS.n6335 VSS.n6334 4.5005
R19936 VSS.n6852 VSS.n6851 4.5005
R19937 VSS.n6853 VSS.n6852 4.5005
R19938 VSS.n6349 VSS.n6347 4.5005
R19939 VSS.n6910 VSS.n6909 4.5005
R19940 VSS.n6781 VSS.n6780 4.5005
R19941 VSS.n6782 VSS.n6392 4.5005
R19942 VSS.n6633 VSS.n6480 4.5005
R19943 VSS.n6632 VSS.n6631 4.5005
R19944 VSS.n6502 VSS.n6501 4.5005
R19945 VSS.n6584 VSS.n6583 4.5005
R19946 VSS.n6557 VSS.n6555 4.5005
R19947 VSS.n6556 VSS.n6533 4.5005
R19948 VSS.n6559 VSS.n6558 4.5005
R19949 VSS.n6491 VSS.n6490 4.5005
R19950 VSS.n6622 VSS.n6621 4.5005
R19951 VSS.n6514 VSS.n6513 4.5005
R19952 VSS.n6593 VSS.n6592 4.5005
R19953 VSS.n6591 VSS.n6590 4.5005
R19954 VSS.n6536 VSS.n6520 4.5005
R19955 VSS.n6495 VSS.n6493 4.5005
R19956 VSS.n6630 VSS.n6482 4.5005
R19957 VSS.n6553 VSS.n6552 4.5005
R19958 VSS.n6635 VSS.n6634 4.5005
R19959 VSS.n6635 VSS.n6478 4.5005
R19960 VSS.n6603 VSS.n6511 4.5005
R19961 VSS.n6582 VSS.n6521 4.5005
R19962 VSS.n6582 VSS.n6581 4.5005
R19963 VSS.n6568 VSS.n6534 4.5005
R19964 VSS.n6500 VSS.n6496 4.5005
R19965 VSS.n6498 VSS.n6496 4.5005
R19966 VSS.n6647 VSS.n6646 4.5005
R19967 VSS.n6646 VSS.n6645 4.5005
R19968 VSS.n2611 VSS.n2610 4.5005
R19969 VSS.n2614 VSS.n2613 4.5005
R19970 VSS.n2597 VSS.n2596 4.5005
R19971 VSS.n2572 VSS.n2571 4.5005
R19972 VSS.n2563 VSS.n2562 4.5005
R19973 VSS.n2564 VSS.n2556 4.5005
R19974 VSS.n2560 VSS.n2557 4.5005
R19975 VSS.n2521 VSS.n2519 4.5005
R19976 VSS.n7013 VSS.n7012 4.5005
R19977 VSS.n7020 VSS.n2511 4.5005
R19978 VSS.n7027 VSS.n7026 4.5005
R19979 VSS.n7028 VSS.n2503 4.5005
R19980 VSS.n2568 VSS.n2500 4.5005
R19981 VSS.n7035 VSS.n7034 4.5005
R19982 VSS.n7019 VSS.n7018 4.5005
R19983 VSS.n2612 VSS.n2536 4.5005
R19984 VSS.n7043 VSS.n7042 4.5005
R19985 VSS.n2609 VSS.n2537 4.5005
R19986 VSS.n2609 VSS.n2608 4.5005
R19987 VSS.n2570 VSS.n2569 4.5005
R19988 VSS.n2569 VSS.n2547 4.5005
R19989 VSS.n2566 VSS.n2565 4.5005
R19990 VSS.n2599 VSS.n2598 4.5005
R19991 VSS.n2599 VSS.n2592 4.5005
R19992 VSS.n7005 VSS.n2529 4.5005
R19993 VSS.n7005 VSS.n7004 4.5005
R19994 VSS.n2762 VSS.n2761 4.5005
R19995 VSS.n2732 VSS.n2681 4.5005
R19996 VSS.n6972 VSS.n6971 4.5005
R19997 VSS.n2639 VSS.n2623 4.5005
R19998 VSS.n2647 VSS.n2646 4.5005
R19999 VSS.n6986 VSS.n2631 4.5005
R20000 VSS.n2631 VSS.n2629 4.5005
R20001 VSS.n2694 VSS.n2693 4.5005
R20002 VSS.n2665 VSS.n2664 4.5005
R20003 VSS.n6970 VSS.n2660 4.5005
R20004 VSS.n2660 VSS.n2658 4.5005
R20005 VSS.n2767 VSS.n2751 4.5005
R20006 VSS.n6944 VSS.n6943 4.5005
R20007 VSS.n6945 VSS.n6944 4.5005
R20008 VSS.n6939 VSS.n2712 4.5005
R20009 VSS.n2734 VSS.n2733 4.5005
R20010 VSS.n2734 VSS.n2729 4.5005
R20011 VSS.n6949 VSS.n2705 4.5005
R20012 VSS.n2699 VSS.n2698 4.5005
R20013 VSS.n2698 VSS.n2676 4.5005
R20014 VSS.n2763 VSS.n2759 4.5005
R20015 VSS.n6931 VSS.n2721 4.5005
R20016 VSS.n6931 VSS.n6930 4.5005
R20017 VSS.n6956 VSS.n6955 4.5005
R20018 VSS.n6957 VSS.n6956 4.5005
R20019 VSS.n6942 VSS.n2710 4.5005
R20020 VSS.n2752 VSS.n2750 4.5005
R20021 VSS.n2632 VSS.n2630 4.5005
R20022 VSS.n2648 VSS.n2636 4.5005
R20023 VSS.n2477 VSS.n2324 4.5005
R20024 VSS.n2476 VSS.n2475 4.5005
R20025 VSS.n2346 VSS.n2345 4.5005
R20026 VSS.n2428 VSS.n2427 4.5005
R20027 VSS.n2401 VSS.n2399 4.5005
R20028 VSS.n2400 VSS.n2377 4.5005
R20029 VSS.n2403 VSS.n2402 4.5005
R20030 VSS.n2335 VSS.n2334 4.5005
R20031 VSS.n2466 VSS.n2465 4.5005
R20032 VSS.n2358 VSS.n2357 4.5005
R20033 VSS.n2437 VSS.n2436 4.5005
R20034 VSS.n2435 VSS.n2434 4.5005
R20035 VSS.n2380 VSS.n2364 4.5005
R20036 VSS.n2339 VSS.n2337 4.5005
R20037 VSS.n2474 VSS.n2326 4.5005
R20038 VSS.n2397 VSS.n2396 4.5005
R20039 VSS.n2479 VSS.n2478 4.5005
R20040 VSS.n2479 VSS.n2322 4.5005
R20041 VSS.n2447 VSS.n2355 4.5005
R20042 VSS.n2426 VSS.n2365 4.5005
R20043 VSS.n2426 VSS.n2425 4.5005
R20044 VSS.n2412 VSS.n2378 4.5005
R20045 VSS.n2344 VSS.n2340 4.5005
R20046 VSS.n2342 VSS.n2340 4.5005
R20047 VSS.n2491 VSS.n2490 4.5005
R20048 VSS.n2490 VSS.n2489 4.5005
R20049 VSS.n2858 VSS.n2853 4.5005
R20050 VSS.n3187 VSS.n3186 4.5005
R20051 VSS.n3164 VSS.n2868 4.5005
R20052 VSS.n2896 VSS.n2894 4.5005
R20053 VSS.n3103 VSS.n3101 4.5005
R20054 VSS.n3102 VSS.n2901 4.5005
R20055 VSS.n3105 VSS.n3104 4.5005
R20056 VSS.n3163 VSS.n3162 4.5005
R20057 VSS.n2870 VSS.n2857 4.5005
R20058 VSS.n3153 VSS.n3152 4.5005
R20059 VSS.n2879 VSS.n2877 4.5005
R20060 VSS.n2891 VSS.n2890 4.5005
R20061 VSS.n3125 VSS.n3124 4.5005
R20062 VSS.n2903 VSS.n2893 4.5005
R20063 VSS.n3154 VSS.n2872 4.5005
R20064 VSS.n3185 VSS.n2852 4.5005
R20065 VSS.n3099 VSS.n3098 4.5005
R20066 VSS.n2860 VSS.n2859 4.5005
R20067 VSS.n3174 VSS.n2860 4.5005
R20068 VSS.n2889 VSS.n2887 4.5005
R20069 VSS.n2887 VSS.n2886 4.5005
R20070 VSS.n3114 VSS.n2902 4.5005
R20071 VSS.n3166 VSS.n3165 4.5005
R20072 VSS.n3166 VSS.n2866 4.5005
R20073 VSS.n3221 VSS.n3220 4.5005
R20074 VSS.n3220 VSS.n3219 4.5005
R20075 VSS.n3344 VSS.n2783 4.5005
R20076 VSS.n3285 VSS.n2810 4.5005
R20077 VSS.n3248 VSS.n3247 4.5005
R20078 VSS.n3198 VSS.n3196 4.5005
R20079 VSS.n3227 VSS.n3226 4.5005
R20080 VSS.n3238 VSS.n3237 4.5005
R20081 VSS.n3239 VSS.n3238 4.5005
R20082 VSS.n3272 VSS.n3271 4.5005
R20083 VSS.n3245 VSS.n3244 4.5005
R20084 VSS.n2819 VSS.n2818 4.5005
R20085 VSS.n2828 VSS.n2819 4.5005
R20086 VSS.n3339 VSS.n3338 4.5005
R20087 VSS.n3312 VSS.n2799 4.5005
R20088 VSS.n3312 VSS.n2793 4.5005
R20089 VSS.n3319 VSS.n2795 4.5005
R20090 VSS.n3290 VSS.n3286 4.5005
R20091 VSS.n3290 VSS.n3289 4.5005
R20092 VSS.n3293 VSS.n3284 4.5005
R20093 VSS.n3277 VSS.n3276 4.5005
R20094 VSS.n3276 VSS.n2805 4.5005
R20095 VSS.n3343 VSS.n3342 4.5005
R20096 VSS.n2784 VSS.n2782 4.5005
R20097 VSS.n2782 VSS.n2781 4.5005
R20098 VSS.n3300 VSS.n3299 4.5005
R20099 VSS.n3301 VSS.n3300 4.5005
R20100 VSS.n2796 VSS.n2794 4.5005
R20101 VSS.n3358 VSS.n3357 4.5005
R20102 VSS.n3229 VSS.n3228 4.5005
R20103 VSS.n3230 VSS.n2839 4.5005
R20104 VSS.n2933 VSS.n2928 4.5005
R20105 VSS.n3083 VSS.n3082 4.5005
R20106 VSS.n3059 VSS.n2943 4.5005
R20107 VSS.n3020 VSS.n3019 4.5005
R20108 VSS.n2998 VSS.n2996 4.5005
R20109 VSS.n2997 VSS.n2976 4.5005
R20110 VSS.n3000 VSS.n2999 4.5005
R20111 VSS.n3058 VSS.n3057 4.5005
R20112 VSS.n2945 VSS.n2932 4.5005
R20113 VSS.n3048 VSS.n3047 4.5005
R20114 VSS.n2954 VSS.n2952 4.5005
R20115 VSS.n2968 VSS.n2967 4.5005
R20116 VSS.n2978 VSS.n2970 4.5005
R20117 VSS.n3049 VSS.n2947 4.5005
R20118 VSS.n3081 VSS.n2927 4.5005
R20119 VSS.n2994 VSS.n2993 4.5005
R20120 VSS.n2935 VSS.n2934 4.5005
R20121 VSS.n3070 VSS.n2935 4.5005
R20122 VSS.n3040 VSS.n2953 4.5005
R20123 VSS.n2966 VSS.n2964 4.5005
R20124 VSS.n2964 VSS.n2963 4.5005
R20125 VSS.n3009 VSS.n2977 4.5005
R20126 VSS.n3061 VSS.n3060 4.5005
R20127 VSS.n3061 VSS.n2941 4.5005
R20128 VSS.n3095 VSS.n3094 4.5005
R20129 VSS.n3094 VSS.n3093 4.5005
R20130 VSS.n125 VSS.n120 4.5005
R20131 VSS.n9147 VSS.n9146 4.5005
R20132 VSS.n9124 VSS.n135 4.5005
R20133 VSS.n163 VSS.n161 4.5005
R20134 VSS.n9063 VSS.n9061 4.5005
R20135 VSS.n9062 VSS.n168 4.5005
R20136 VSS.n9065 VSS.n9064 4.5005
R20137 VSS.n9123 VSS.n9122 4.5005
R20138 VSS.n137 VSS.n124 4.5005
R20139 VSS.n9113 VSS.n9112 4.5005
R20140 VSS.n146 VSS.n144 4.5005
R20141 VSS.n158 VSS.n157 4.5005
R20142 VSS.n9085 VSS.n9084 4.5005
R20143 VSS.n170 VSS.n160 4.5005
R20144 VSS.n9114 VSS.n139 4.5005
R20145 VSS.n9145 VSS.n119 4.5005
R20146 VSS.n9059 VSS.n9058 4.5005
R20147 VSS.n127 VSS.n126 4.5005
R20148 VSS.n9134 VSS.n127 4.5005
R20149 VSS.n156 VSS.n154 4.5005
R20150 VSS.n154 VSS.n153 4.5005
R20151 VSS.n9074 VSS.n169 4.5005
R20152 VSS.n9126 VSS.n9125 4.5005
R20153 VSS.n9126 VSS.n133 4.5005
R20154 VSS.n9181 VSS.n9180 4.5005
R20155 VSS.n9180 VSS.n9179 4.5005
R20156 VSS.n9304 VSS.n50 4.5005
R20157 VSS.n9245 VSS.n77 4.5005
R20158 VSS.n9208 VSS.n9207 4.5005
R20159 VSS.n9158 VSS.n9156 4.5005
R20160 VSS.n9187 VSS.n9186 4.5005
R20161 VSS.n9198 VSS.n9197 4.5005
R20162 VSS.n9199 VSS.n9198 4.5005
R20163 VSS.n9232 VSS.n9231 4.5005
R20164 VSS.n9205 VSS.n9204 4.5005
R20165 VSS.n86 VSS.n85 4.5005
R20166 VSS.n95 VSS.n86 4.5005
R20167 VSS.n9299 VSS.n9298 4.5005
R20168 VSS.n9272 VSS.n66 4.5005
R20169 VSS.n9272 VSS.n60 4.5005
R20170 VSS.n9279 VSS.n62 4.5005
R20171 VSS.n9250 VSS.n9246 4.5005
R20172 VSS.n9250 VSS.n9249 4.5005
R20173 VSS.n9253 VSS.n9244 4.5005
R20174 VSS.n9237 VSS.n9236 4.5005
R20175 VSS.n9236 VSS.n72 4.5005
R20176 VSS.n9303 VSS.n9302 4.5005
R20177 VSS.n51 VSS.n49 4.5005
R20178 VSS.n49 VSS.n48 4.5005
R20179 VSS.n9260 VSS.n9259 4.5005
R20180 VSS.n9261 VSS.n9260 4.5005
R20181 VSS.n63 VSS.n61 4.5005
R20182 VSS.n9318 VSS.n9317 4.5005
R20183 VSS.n9189 VSS.n9188 4.5005
R20184 VSS.n9190 VSS.n106 4.5005
R20185 VSS.n392 VSS.n391 4.5005
R20186 VSS.n394 VSS.n393 4.5005
R20187 VSS.n375 VSS.n374 4.5005
R20188 VSS.n351 VSS.n283 4.5005
R20189 VSS.n335 VSS.n329 4.5005
R20190 VSS.n338 VSS.n337 4.5005
R20191 VSS.n334 VSS.n333 4.5005
R20192 VSS.n305 VSS.n303 4.5005
R20193 VSS.n404 VSS.n403 4.5005
R20194 VSS.n411 VSS.n295 4.5005
R20195 VSS.n418 VSS.n417 4.5005
R20196 VSS.n419 VSS.n286 4.5005
R20197 VSS.n426 VSS.n425 4.5005
R20198 VSS.n410 VSS.n409 4.5005
R20199 VSS.n395 VSS.n308 4.5005
R20200 VSS.n434 VSS.n433 4.5005
R20201 VSS.n311 VSS.n310 4.5005
R20202 VSS.n312 VSS.n311 4.5005
R20203 VSS.n362 VSS.n291 4.5005
R20204 VSS.n353 VSS.n352 4.5005
R20205 VSS.n353 VSS.n326 4.5005
R20206 VSS.n336 VSS.n330 4.5005
R20207 VSS.n373 VSS.n372 4.5005
R20208 VSS.n372 VSS.n316 4.5005
R20209 VSS.n9055 VSS.n9054 4.5005
R20210 VSS.n9054 VSS.n9053 4.5005
R20211 VSS.n603 VSS.n602 4.5005
R20212 VSS.n606 VSS.n605 4.5005
R20213 VSS.n589 VSS.n588 4.5005
R20214 VSS.n564 VSS.n563 4.5005
R20215 VSS.n555 VSS.n554 4.5005
R20216 VSS.n556 VSS.n550 4.5005
R20217 VSS.n552 VSS.n551 4.5005
R20218 VSS.n510 VSS.n508 4.5005
R20219 VSS.n832 VSS.n831 4.5005
R20220 VSS.n839 VSS.n500 4.5005
R20221 VSS.n846 VSS.n845 4.5005
R20222 VSS.n847 VSS.n492 4.5005
R20223 VSS.n560 VSS.n489 4.5005
R20224 VSS.n854 VSS.n853 4.5005
R20225 VSS.n838 VSS.n837 4.5005
R20226 VSS.n604 VSS.n525 4.5005
R20227 VSS.n862 VSS.n861 4.5005
R20228 VSS.n601 VSS.n526 4.5005
R20229 VSS.n601 VSS.n600 4.5005
R20230 VSS.n562 VSS.n561 4.5005
R20231 VSS.n561 VSS.n536 4.5005
R20232 VSS.n558 VSS.n557 4.5005
R20233 VSS.n591 VSS.n590 4.5005
R20234 VSS.n591 VSS.n584 4.5005
R20235 VSS.n824 VSS.n518 4.5005
R20236 VSS.n824 VSS.n823 4.5005
R20237 VSS.n716 VSS.n33 4.5005
R20238 VSS.n723 VSS.n722 4.5005
R20239 VSS.n768 VSS.n697 4.5005
R20240 VSS.n789 VSS.n652 4.5005
R20241 VSS.n652 VSS.n650 4.5005
R20242 VSS.n639 VSS.n638 4.5005
R20243 VSS.n631 VSS.n615 4.5005
R20244 VSS.n657 VSS.n656 4.5005
R20245 VSS.n640 VSS.n628 4.5005
R20246 VSS.n805 VSS.n623 4.5005
R20247 VSS.n623 VSS.n621 4.5005
R20248 VSS.n686 VSS.n685 4.5005
R20249 VSS.n691 VSS.n690 4.5005
R20250 VSS.n690 VSS.n668 4.5005
R20251 VSS.n775 VSS.n774 4.5005
R20252 VSS.n776 VSS.n775 4.5005
R20253 VSS.n735 VSS.n734 4.5005
R20254 VSS.n735 VSS.n730 4.5005
R20255 VSS.n763 VSS.n762 4.5005
R20256 VSS.n764 VSS.n763 4.5005
R20257 VSS.n758 VSS.n704 4.5005
R20258 VSS.n750 VSS.n713 4.5005
R20259 VSS.n750 VSS.n749 4.5005
R20260 VSS.n34 VSS.n27 4.5005
R20261 VSS.n761 VSS.n702 4.5005
R20262 VSS.n624 VSS.n622 4.5005
R20263 VSS.n724 VSS.n715 4.5005
R20264 VSS.n733 VSS.n673 4.5005
R20265 VSS.n791 VSS.n790 4.5005
R20266 VSS.n947 VSS.n946 4.5005
R20267 VSS.n950 VSS.n949 4.5005
R20268 VSS.n932 VSS.n931 4.5005
R20269 VSS.n907 VSS.n449 4.5005
R20270 VSS.n900 VSS.n899 4.5005
R20271 VSS.n901 VSS.n893 4.5005
R20272 VSS.n897 VSS.n894 4.5005
R20273 VSS.n471 VSS.n469 4.5005
R20274 VSS.n969 VSS.n968 4.5005
R20275 VSS.n976 VSS.n461 4.5005
R20276 VSS.n983 VSS.n982 4.5005
R20277 VSS.n984 VSS.n452 4.5005
R20278 VSS.n991 VSS.n990 4.5005
R20279 VSS.n975 VSS.n974 4.5005
R20280 VSS.n948 VSS.n872 4.5005
R20281 VSS.n999 VSS.n998 4.5005
R20282 VSS.n945 VSS.n873 4.5005
R20283 VSS.n945 VSS.n944 4.5005
R20284 VSS.n879 VSS.n457 4.5005
R20285 VSS.n906 VSS.n905 4.5005
R20286 VSS.n906 VSS.n884 4.5005
R20287 VSS.n903 VSS.n902 4.5005
R20288 VSS.n934 VSS.n933 4.5005
R20289 VSS.n934 VSS.n927 4.5005
R20290 VSS.n961 VSS.n865 4.5005
R20291 VSS.n961 VSS.n960 4.5005
R20292 VSS.n7330 VSS.n7329 4.5005
R20293 VSS.n7300 VSS.n7249 4.5005
R20294 VSS.n8400 VSS.n8399 4.5005
R20295 VSS.n7207 VSS.n7191 4.5005
R20296 VSS.n7215 VSS.n7214 4.5005
R20297 VSS.n8414 VSS.n7199 4.5005
R20298 VSS.n7199 VSS.n7197 4.5005
R20299 VSS.n7262 VSS.n7261 4.5005
R20300 VSS.n7233 VSS.n7232 4.5005
R20301 VSS.n8398 VSS.n7228 4.5005
R20302 VSS.n7228 VSS.n7226 4.5005
R20303 VSS.n7335 VSS.n7319 4.5005
R20304 VSS.n8372 VSS.n8371 4.5005
R20305 VSS.n8373 VSS.n8372 4.5005
R20306 VSS.n8367 VSS.n7280 4.5005
R20307 VSS.n7302 VSS.n7301 4.5005
R20308 VSS.n7302 VSS.n7297 4.5005
R20309 VSS.n8377 VSS.n7273 4.5005
R20310 VSS.n7267 VSS.n7266 4.5005
R20311 VSS.n7266 VSS.n7244 4.5005
R20312 VSS.n7331 VSS.n7327 4.5005
R20313 VSS.n8359 VSS.n7289 4.5005
R20314 VSS.n8359 VSS.n8358 4.5005
R20315 VSS.n8384 VSS.n8383 4.5005
R20316 VSS.n8385 VSS.n8384 4.5005
R20317 VSS.n8370 VSS.n7278 4.5005
R20318 VSS.n7320 VSS.n7318 4.5005
R20319 VSS.n7200 VSS.n7198 4.5005
R20320 VSS.n7216 VSS.n7204 4.5005
R20321 VSS.n7608 VSS.n7414 3.69976
R20322 VSS.n8200 VSS.n7828 3.69976
R20323 VSS.n1667 VSS.n1357 3.69976
R20324 VSS.n2259 VSS.n1930 3.69976
R20325 VSS.n3810 VSS.n3438 3.69976
R20326 VSS.n4402 VSS.n4030 3.69976
R20327 VSS.n4994 VSS.n4622 3.69976
R20328 VSS.n5586 VSS.n5214 3.69976
R20329 VSS.n6178 VSS.n5806 3.69976
R20330 VSS.n6770 VSS.n6398 3.69976
R20331 VSS.n7003 VSS.n2528 3.69976
R20332 VSS.n3218 VSS.n2845 3.69976
R20333 VSS.n9178 VSS.n112 3.69976
R20334 VSS.n9004 VSS.n8675 3.69976
R20335 VSS.n822 VSS.n517 3.69976
R20336 VSS.n8431 VSS.n7096 3.69976
R20337 VSS.n8635 VSS.n200 3.69922
R20338 VSS.n1317 VSS.n1146 3.69922
R20339 VSS.n1890 VSS.n1719 3.69922
R20340 VSS.n3684 VSS.n3513 3.69922
R20341 VSS.n4276 VSS.n4105 3.69922
R20342 VSS.n4868 VSS.n4697 3.69922
R20343 VSS.n5460 VSS.n5289 3.69922
R20344 VSS.n6052 VSS.n5881 3.69922
R20345 VSS.n6644 VSS.n6473 3.69922
R20346 VSS.n2488 VSS.n2317 3.69922
R20347 VSS.n3092 VSS.n2920 3.69922
R20348 VSS.n9052 VSS.n180 3.69922
R20349 VSS.n959 VSS.n478 3.69922
R20350 VSS.n8480 VSS.n1045 3.69922
R20351 VSS.n8074 VSS.n7903 3.69922
R20352 VSS.n8470 VSS.n7061 3.42389
R20353 VSS.n7486 VSS.n1046 3.42389
R20354 VSS.n7488 VSS.n7487 3.42389
R20355 VSS.n8078 VSS.n8077 3.42389
R20356 VSS.n8080 VSS.n8079 3.42389
R20357 VSS.n9043 VSS.n8640 3.42389
R20358 VSS.n8639 VSS.n8638 3.42389
R20359 VSS.n1706 VSS.n1322 3.42389
R20360 VSS.n1321 VSS.n1320 3.42389
R20361 VSS.n2298 VSS.n1895 3.42389
R20362 VSS.n1894 VSS.n1893 3.42389
R20363 VSS.n3690 VSS.n3689 3.42389
R20364 VSS.n3688 VSS.n3687 3.42389
R20365 VSS.n4282 VSS.n4281 3.42389
R20366 VSS.n4280 VSS.n4279 3.42389
R20367 VSS.n4874 VSS.n4873 3.42389
R20368 VSS.n4872 VSS.n4871 3.42389
R20369 VSS.n5466 VSS.n5465 3.42389
R20370 VSS.n5464 VSS.n5463 3.42389
R20371 VSS.n6058 VSS.n6057 3.42389
R20372 VSS.n6056 VSS.n6055 3.42389
R20373 VSS.n6650 VSS.n6649 3.42389
R20374 VSS.n6648 VSS.n6647 3.42389
R20375 VSS.n7042 VSS.n2493 3.42389
R20376 VSS.n2492 VSS.n2491 3.42389
R20377 VSS.n3098 VSS.n3097 3.42389
R20378 VSS.n3096 VSS.n3095 3.42389
R20379 VSS.n9058 VSS.n9057 3.42389
R20380 VSS.n9056 VSS.n9055 3.42389
R20381 VSS.n863 VSS.n862 3.42389
R20382 VSS.n865 VSS.n864 3.42389
R20383 VSS.n7210 VSS.n7097 3.423
R20384 VSS.n8519 VSS.n1009 3.423
R20385 VSS.n7612 VSS.n7611 3.423
R20386 VSS.n7982 VSS.n7981 3.423
R20387 VSS.n8204 VSS.n8203 3.423
R20388 VSS.n8790 VSS.n8676 3.423
R20389 VSS.n8543 VSS.n8542 3.423
R20390 VSS.n1471 VSS.n1358 3.423
R20391 VSS.n1225 VSS.n1224 3.423
R20392 VSS.n2044 VSS.n1931 3.423
R20393 VSS.n1798 VSS.n1797 3.423
R20394 VSS.n3814 VSS.n3813 3.423
R20395 VSS.n3592 VSS.n3591 3.423
R20396 VSS.n4406 VSS.n4405 3.423
R20397 VSS.n4184 VSS.n4183 3.423
R20398 VSS.n4998 VSS.n4997 3.423
R20399 VSS.n4776 VSS.n4775 3.423
R20400 VSS.n5590 VSS.n5589 3.423
R20401 VSS.n5368 VSS.n5367 3.423
R20402 VSS.n6182 VSS.n6181 3.423
R20403 VSS.n5960 VSS.n5959 3.423
R20404 VSS.n6774 VSS.n6773 3.423
R20405 VSS.n6552 VSS.n6551 3.423
R20406 VSS.n2642 VSS.n2529 3.423
R20407 VSS.n2396 VSS.n2395 3.423
R20408 VSS.n3222 VSS.n3221 3.423
R20409 VSS.n2993 VSS.n2992 3.423
R20410 VSS.n9182 VSS.n9181 3.423
R20411 VSS.n433 VSS.n276 3.423
R20412 VSS.n634 VSS.n518 3.423
R20413 VSS.n998 VSS.n442 3.423
R20414 VSS.n7731 VSS.n7726 3.4105
R20415 VSS.n7731 VSS.n7730 3.4105
R20416 VSS.n7725 VSS.n7353 3.4105
R20417 VSS.n7750 VSS.n7749 3.4105
R20418 VSS.n7749 VSS.n7748 3.4105
R20419 VSS.n7708 VSS.n7706 3.4105
R20420 VSS.n7708 VSS.n7707 3.4105
R20421 VSS.n7724 VSS.n7723 3.4105
R20422 VSS.n7723 VSS.n7722 3.4105
R20423 VSS.n7686 VSS.n7685 3.4105
R20424 VSS.n7685 VSS.n7684 3.4105
R20425 VSS.n7367 VSS.n7366 3.4105
R20426 VSS.n7705 VSS.n7704 3.4105
R20427 VSS.n7704 VSS.n7703 3.4105
R20428 VSS.n7669 VSS.n7668 3.4105
R20429 VSS.n7688 VSS.n7687 3.4105
R20430 VSS.n7653 VSS.n7652 3.4105
R20431 VSS.n7652 VSS.n7651 3.4105
R20432 VSS.n7654 VSS.n7385 3.4105
R20433 VSS.n7657 VSS.n7380 3.4105
R20434 VSS.n7626 VSS.n7625 3.4105
R20435 VSS.n7626 VSS.n7403 3.4105
R20436 VSS.n7399 VSS.n7386 3.4105
R20437 VSS.n7633 VSS.n7399 3.4105
R20438 VSS.n8485 VSS.n8484 3.4105
R20439 VSS.n8484 VSS.n8483 3.4105
R20440 VSS.n8492 VSS.n8491 3.4105
R20441 VSS.n8487 VSS.n8486 3.4105
R20442 VSS.n8488 VSS.n8487 3.4105
R20443 VSS.n8500 VSS.n8499 3.4105
R20444 VSS.n8499 VSS.n8498 3.4105
R20445 VSS.n1031 VSS.n1026 3.4105
R20446 VSS.n8494 VSS.n8493 3.4105
R20447 VSS.n8494 VSS.n1030 3.4105
R20448 VSS.n8508 VSS.n8507 3.4105
R20449 VSS.n8507 VSS.n8506 3.4105
R20450 VSS.n1025 VSS.n1023 3.4105
R20451 VSS.n8502 VSS.n8501 3.4105
R20452 VSS.n8502 VSS.n1021 3.4105
R20453 VSS.n8515 VSS.n8514 3.4105
R20454 VSS.n8514 VSS.n8513 3.4105
R20455 VSS.n8510 VSS.n8509 3.4105
R20456 VSS.n8516 VSS.n1010 3.4105
R20457 VSS.n1010 VSS.n1008 3.4105
R20458 VSS.n7613 VSS.n7410 3.4105
R20459 VSS.n7587 VSS.n7410 3.4105
R20460 VSS.n7407 VSS.n7406 3.4105
R20461 VSS.n7623 VSS.n7622 3.4105
R20462 VSS.n7622 VSS.n7621 3.4105
R20463 VSS.n7572 VSS.n7571 3.4105
R20464 VSS.n7572 VSS.n7413 3.4105
R20465 VSS.n7549 VSS.n7548 3.4105
R20466 VSS.n7570 VSS.n7569 3.4105
R20467 VSS.n7569 VSS.n7568 3.4105
R20468 VSS.n7539 VSS.n7443 3.4105
R20469 VSS.n7443 VSS.n7442 3.4105
R20470 VSS.n7541 VSS.n7540 3.4105
R20471 VSS.n7547 VSS.n7546 3.4105
R20472 VSS.n7546 VSS.n7545 3.4105
R20473 VSS.n7522 VSS.n7521 3.4105
R20474 VSS.n7522 VSS.n7457 3.4105
R20475 VSS.n7518 VSS.n7445 3.4105
R20476 VSS.n7538 VSS.n7537 3.4105
R20477 VSS.n7537 VSS.n7536 3.4105
R20478 VSS.n7501 VSS.n7500 3.4105
R20479 VSS.n7501 VSS.n7473 3.4105
R20480 VSS.n7517 VSS.n7516 3.4105
R20481 VSS.n7499 VSS.n7498 3.4105
R20482 VSS.n7498 VSS.n7497 3.4105
R20483 VSS.n8323 VSS.n8318 3.4105
R20484 VSS.n8323 VSS.n8322 3.4105
R20485 VSS.n8317 VSS.n7767 3.4105
R20486 VSS.n8342 VSS.n8341 3.4105
R20487 VSS.n8341 VSS.n8340 3.4105
R20488 VSS.n8300 VSS.n8298 3.4105
R20489 VSS.n8300 VSS.n8299 3.4105
R20490 VSS.n8316 VSS.n8315 3.4105
R20491 VSS.n8315 VSS.n8314 3.4105
R20492 VSS.n8278 VSS.n8277 3.4105
R20493 VSS.n8277 VSS.n8276 3.4105
R20494 VSS.n7781 VSS.n7780 3.4105
R20495 VSS.n8297 VSS.n8296 3.4105
R20496 VSS.n8296 VSS.n8295 3.4105
R20497 VSS.n8261 VSS.n8260 3.4105
R20498 VSS.n8280 VSS.n8279 3.4105
R20499 VSS.n8245 VSS.n8244 3.4105
R20500 VSS.n8244 VSS.n8243 3.4105
R20501 VSS.n8246 VSS.n7799 3.4105
R20502 VSS.n8249 VSS.n7794 3.4105
R20503 VSS.n8218 VSS.n8217 3.4105
R20504 VSS.n8218 VSS.n7817 3.4105
R20505 VSS.n7813 VSS.n7800 3.4105
R20506 VSS.n8225 VSS.n7813 3.4105
R20507 VSS.n8057 VSS.n8056 3.4105
R20508 VSS.n8057 VSS.n7902 3.4105
R20509 VSS.n8050 VSS.n8049 3.4105
R20510 VSS.n8055 VSS.n8054 3.4105
R20511 VSS.n8054 VSS.n8053 3.4105
R20512 VSS.n8030 VSS.n8029 3.4105
R20513 VSS.n8030 VSS.n7942 3.4105
R20514 VSS.n8028 VSS.n8027 3.4105
R20515 VSS.n8048 VSS.n8047 3.4105
R20516 VSS.n8047 VSS.n8046 3.4105
R20517 VSS.n8017 VSS.n7948 3.4105
R20518 VSS.n7948 VSS.n7947 3.4105
R20519 VSS.n7946 VSS.n7945 3.4105
R20520 VSS.n8025 VSS.n8024 3.4105
R20521 VSS.n8024 VSS.n7940 3.4105
R20522 VSS.n7995 VSS.n7994 3.4105
R20523 VSS.n7995 VSS.n7967 3.4105
R20524 VSS.n8016 VSS.n8015 3.4105
R20525 VSS.n7993 VSS.n7992 3.4105
R20526 VSS.n7992 VSS.n7991 3.4105
R20527 VSS.n8205 VSS.n7824 3.4105
R20528 VSS.n8179 VSS.n7824 3.4105
R20529 VSS.n7821 VSS.n7820 3.4105
R20530 VSS.n8215 VSS.n8214 3.4105
R20531 VSS.n8214 VSS.n8213 3.4105
R20532 VSS.n8164 VSS.n8163 3.4105
R20533 VSS.n8164 VSS.n7827 3.4105
R20534 VSS.n8141 VSS.n8140 3.4105
R20535 VSS.n8162 VSS.n8161 3.4105
R20536 VSS.n8161 VSS.n8160 3.4105
R20537 VSS.n8131 VSS.n7857 3.4105
R20538 VSS.n7857 VSS.n7856 3.4105
R20539 VSS.n8133 VSS.n8132 3.4105
R20540 VSS.n8139 VSS.n8138 3.4105
R20541 VSS.n8138 VSS.n8137 3.4105
R20542 VSS.n8114 VSS.n8113 3.4105
R20543 VSS.n8114 VSS.n7871 3.4105
R20544 VSS.n8110 VSS.n7859 3.4105
R20545 VSS.n8130 VSS.n8129 3.4105
R20546 VSS.n8129 VSS.n8128 3.4105
R20547 VSS.n8093 VSS.n8092 3.4105
R20548 VSS.n8093 VSS.n7887 3.4105
R20549 VSS.n8109 VSS.n8108 3.4105
R20550 VSS.n8091 VSS.n8090 3.4105
R20551 VSS.n8090 VSS.n8089 3.4105
R20552 VSS.n8934 VSS.n8933 3.4105
R20553 VSS.n8935 VSS.n8934 3.4105
R20554 VSS.n8932 VSS.n8890 3.4105
R20555 VSS.n8929 VSS.n8893 3.4105
R20556 VSS.n8929 VSS.n8928 3.4105
R20557 VSS.n8948 VSS.n8947 3.4105
R20558 VSS.n8947 VSS.n8946 3.4105
R20559 VSS.n8891 VSS.n8887 3.4105
R20560 VSS.n8887 VSS.n8885 3.4105
R20561 VSS.n8873 VSS.n8855 3.4105
R20562 VSS.n8873 VSS.n8872 3.4105
R20563 VSS.n8877 VSS.n8853 3.4105
R20564 VSS.n8950 VSS.n8949 3.4105
R20565 VSS.n8951 VSS.n8950 3.4105
R20566 VSS.n8966 VSS.n8965 3.4105
R20567 VSS.n8862 VSS.n8861 3.4105
R20568 VSS.n8811 VSS.n8800 3.4105
R20569 VSS.n8811 VSS.n8805 3.4105
R20570 VSS.n8813 VSS.n8812 3.4105
R20571 VSS.n8968 VSS.n8967 3.4105
R20572 VSS.n8986 VSS.n8985 3.4105
R20573 VSS.n8986 VSS.n8779 3.4105
R20574 VSS.n8983 VSS.n8982 3.4105
R20575 VSS.n8982 VSS.n8981 3.4105
R20576 VSS.n9009 VSS.n9008 3.4105
R20577 VSS.n9008 VSS.n9007 3.4105
R20578 VSS.n9016 VSS.n9015 3.4105
R20579 VSS.n9011 VSS.n9010 3.4105
R20580 VSS.n9012 VSS.n9011 3.4105
R20581 VSS.n9024 VSS.n9023 3.4105
R20582 VSS.n9023 VSS.n9022 3.4105
R20583 VSS.n8661 VSS.n8657 3.4105
R20584 VSS.n9018 VSS.n9017 3.4105
R20585 VSS.n9018 VSS.n8660 3.4105
R20586 VSS.n9032 VSS.n9031 3.4105
R20587 VSS.n9031 VSS.n9030 3.4105
R20588 VSS.n8656 VSS.n8654 3.4105
R20589 VSS.n9026 VSS.n9025 3.4105
R20590 VSS.n9026 VSS.n8652 3.4105
R20591 VSS.n9039 VSS.n9038 3.4105
R20592 VSS.n9038 VSS.n9037 3.4105
R20593 VSS.n9034 VSS.n9033 3.4105
R20594 VSS.n9040 VSS.n8641 3.4105
R20595 VSS.n8641 VSS.n196 3.4105
R20596 VSS.n8791 VSS.n8789 3.4105
R20597 VSS.n8789 VSS.n8788 3.4105
R20598 VSS.n8782 VSS.n8781 3.4105
R20599 VSS.n8799 VSS.n8798 3.4105
R20600 VSS.n8798 VSS.n8797 3.4105
R20601 VSS.n8618 VSS.n8617 3.4105
R20602 VSS.n8618 VSS.n199 3.4105
R20603 VSS.n8611 VSS.n8610 3.4105
R20604 VSS.n8616 VSS.n8615 3.4105
R20605 VSS.n8615 VSS.n8614 3.4105
R20606 VSS.n8591 VSS.n8590 3.4105
R20607 VSS.n8591 VSS.n239 3.4105
R20608 VSS.n8589 VSS.n8588 3.4105
R20609 VSS.n8609 VSS.n8608 3.4105
R20610 VSS.n8608 VSS.n8607 3.4105
R20611 VSS.n8578 VSS.n245 3.4105
R20612 VSS.n245 VSS.n244 3.4105
R20613 VSS.n243 VSS.n242 3.4105
R20614 VSS.n8586 VSS.n8585 3.4105
R20615 VSS.n8585 VSS.n237 3.4105
R20616 VSS.n8556 VSS.n8555 3.4105
R20617 VSS.n8556 VSS.n264 3.4105
R20618 VSS.n8577 VSS.n8576 3.4105
R20619 VSS.n8554 VSS.n8553 3.4105
R20620 VSS.n8553 VSS.n8552 3.4105
R20621 VSS.n1553 VSS.n1549 3.4105
R20622 VSS.n1559 VSS.n1553 3.4105
R20623 VSS.n1555 VSS.n1554 3.4105
R20624 VSS.n9350 VSS.n9349 3.4105
R20625 VSS.n9349 VSS.n9348 3.4105
R20626 VSS.n1601 VSS.n1600 3.4105
R20627 VSS.n1602 VSS.n1601 3.4105
R20628 VSS.n1598 VSS.n1597 3.4105
R20629 VSS.n1597 VSS.n1596 3.4105
R20630 VSS.n1616 VSS.n1615 3.4105
R20631 VSS.n1615 VSS.n1614 3.4105
R20632 VSS.n1547 VSS.n1546 3.4105
R20633 VSS.n1548 VSS.n1540 3.4105
R20634 VSS.n1540 VSS.n1536 3.4105
R20635 VSS.n1530 VSS.n1529 3.4105
R20636 VSS.n1618 VSS.n1617 3.4105
R20637 VSS.n1633 VSS.n1498 3.4105
R20638 VSS.n1633 VSS.n1632 3.4105
R20639 VSS.n1515 VSS.n1491 3.4105
R20640 VSS.n1518 VSS.n1511 3.4105
R20641 VSS.n1649 VSS.n1481 3.4105
R20642 VSS.n1649 VSS.n1648 3.4105
R20643 VSS.n1497 VSS.n1496 3.4105
R20644 VSS.n1496 VSS.n1495 3.4105
R20645 VSS.n1672 VSS.n1671 3.4105
R20646 VSS.n1671 VSS.n1670 3.4105
R20647 VSS.n1679 VSS.n1678 3.4105
R20648 VSS.n1674 VSS.n1673 3.4105
R20649 VSS.n1675 VSS.n1674 3.4105
R20650 VSS.n1687 VSS.n1686 3.4105
R20651 VSS.n1686 VSS.n1685 3.4105
R20652 VSS.n1343 VSS.n1339 3.4105
R20653 VSS.n1681 VSS.n1680 3.4105
R20654 VSS.n1681 VSS.n1342 3.4105
R20655 VSS.n1695 VSS.n1694 3.4105
R20656 VSS.n1694 VSS.n1693 3.4105
R20657 VSS.n1338 VSS.n1336 3.4105
R20658 VSS.n1689 VSS.n1688 3.4105
R20659 VSS.n1689 VSS.n1334 3.4105
R20660 VSS.n1702 VSS.n1701 3.4105
R20661 VSS.n1701 VSS.n1700 3.4105
R20662 VSS.n1697 VSS.n1696 3.4105
R20663 VSS.n1703 VSS.n1323 3.4105
R20664 VSS.n1323 VSS.n1142 3.4105
R20665 VSS.n1472 VSS.n1470 3.4105
R20666 VSS.n1470 VSS.n1469 3.4105
R20667 VSS.n1464 VSS.n1463 3.4105
R20668 VSS.n1480 VSS.n1479 3.4105
R20669 VSS.n1479 VSS.n1478 3.4105
R20670 VSS.n1300 VSS.n1299 3.4105
R20671 VSS.n1300 VSS.n1145 3.4105
R20672 VSS.n1293 VSS.n1292 3.4105
R20673 VSS.n1298 VSS.n1297 3.4105
R20674 VSS.n1297 VSS.n1296 3.4105
R20675 VSS.n1273 VSS.n1272 3.4105
R20676 VSS.n1273 VSS.n1185 3.4105
R20677 VSS.n1271 VSS.n1270 3.4105
R20678 VSS.n1291 VSS.n1290 3.4105
R20679 VSS.n1290 VSS.n1289 3.4105
R20680 VSS.n1260 VSS.n1191 3.4105
R20681 VSS.n1191 VSS.n1190 3.4105
R20682 VSS.n1189 VSS.n1188 3.4105
R20683 VSS.n1268 VSS.n1267 3.4105
R20684 VSS.n1267 VSS.n1183 3.4105
R20685 VSS.n1238 VSS.n1237 3.4105
R20686 VSS.n1238 VSS.n1210 3.4105
R20687 VSS.n1259 VSS.n1258 3.4105
R20688 VSS.n1236 VSS.n1235 3.4105
R20689 VSS.n1235 VSS.n1234 3.4105
R20690 VSS.n2168 VSS.n2122 3.4105
R20691 VSS.n2168 VSS.n2167 3.4105
R20692 VSS.n2171 VSS.n2170 3.4105
R20693 VSS.n2175 VSS.n2174 3.4105
R20694 VSS.n2176 VSS.n2175 3.4105
R20695 VSS.n2193 VSS.n2192 3.4105
R20696 VSS.n2194 VSS.n2193 3.4105
R20697 VSS.n2190 VSS.n2189 3.4105
R20698 VSS.n2189 VSS.n2188 3.4105
R20699 VSS.n2208 VSS.n2207 3.4105
R20700 VSS.n2207 VSS.n2206 3.4105
R20701 VSS.n2120 VSS.n2119 3.4105
R20702 VSS.n2121 VSS.n2113 3.4105
R20703 VSS.n2113 VSS.n2109 3.4105
R20704 VSS.n2103 VSS.n2102 3.4105
R20705 VSS.n2210 VSS.n2209 3.4105
R20706 VSS.n2225 VSS.n2071 3.4105
R20707 VSS.n2225 VSS.n2224 3.4105
R20708 VSS.n2088 VSS.n2064 3.4105
R20709 VSS.n2091 VSS.n2084 3.4105
R20710 VSS.n2241 VSS.n2054 3.4105
R20711 VSS.n2241 VSS.n2240 3.4105
R20712 VSS.n2070 VSS.n2069 3.4105
R20713 VSS.n2069 VSS.n2068 3.4105
R20714 VSS.n2264 VSS.n2263 3.4105
R20715 VSS.n2263 VSS.n2262 3.4105
R20716 VSS.n2271 VSS.n2270 3.4105
R20717 VSS.n2266 VSS.n2265 3.4105
R20718 VSS.n2267 VSS.n2266 3.4105
R20719 VSS.n2279 VSS.n2278 3.4105
R20720 VSS.n2278 VSS.n2277 3.4105
R20721 VSS.n1916 VSS.n1912 3.4105
R20722 VSS.n2273 VSS.n2272 3.4105
R20723 VSS.n2273 VSS.n1915 3.4105
R20724 VSS.n2287 VSS.n2286 3.4105
R20725 VSS.n2286 VSS.n2285 3.4105
R20726 VSS.n1911 VSS.n1909 3.4105
R20727 VSS.n2281 VSS.n2280 3.4105
R20728 VSS.n2281 VSS.n1907 3.4105
R20729 VSS.n2294 VSS.n2293 3.4105
R20730 VSS.n2293 VSS.n2292 3.4105
R20731 VSS.n2289 VSS.n2288 3.4105
R20732 VSS.n2295 VSS.n1896 3.4105
R20733 VSS.n1896 VSS.n1715 3.4105
R20734 VSS.n2045 VSS.n2043 3.4105
R20735 VSS.n2043 VSS.n2042 3.4105
R20736 VSS.n2037 VSS.n2036 3.4105
R20737 VSS.n2053 VSS.n2052 3.4105
R20738 VSS.n2052 VSS.n2051 3.4105
R20739 VSS.n1873 VSS.n1872 3.4105
R20740 VSS.n1873 VSS.n1718 3.4105
R20741 VSS.n1866 VSS.n1865 3.4105
R20742 VSS.n1871 VSS.n1870 3.4105
R20743 VSS.n1870 VSS.n1869 3.4105
R20744 VSS.n1846 VSS.n1845 3.4105
R20745 VSS.n1846 VSS.n1758 3.4105
R20746 VSS.n1844 VSS.n1843 3.4105
R20747 VSS.n1864 VSS.n1863 3.4105
R20748 VSS.n1863 VSS.n1862 3.4105
R20749 VSS.n1833 VSS.n1764 3.4105
R20750 VSS.n1764 VSS.n1763 3.4105
R20751 VSS.n1762 VSS.n1761 3.4105
R20752 VSS.n1841 VSS.n1840 3.4105
R20753 VSS.n1840 VSS.n1756 3.4105
R20754 VSS.n1811 VSS.n1810 3.4105
R20755 VSS.n1811 VSS.n1783 3.4105
R20756 VSS.n1832 VSS.n1831 3.4105
R20757 VSS.n1809 VSS.n1808 3.4105
R20758 VSS.n1808 VSS.n1807 3.4105
R20759 VSS.n3927 VSS.n3378 3.4105
R20760 VSS.n3933 VSS.n3378 3.4105
R20761 VSS.n3929 VSS.n3928 3.4105
R20762 VSS.n3953 VSS.n3952 3.4105
R20763 VSS.n3952 VSS.n3951 3.4105
R20764 VSS.n3910 VSS.n3908 3.4105
R20765 VSS.n3910 VSS.n3909 3.4105
R20766 VSS.n3926 VSS.n3925 3.4105
R20767 VSS.n3925 VSS.n3924 3.4105
R20768 VSS.n3888 VSS.n3887 3.4105
R20769 VSS.n3887 VSS.n3886 3.4105
R20770 VSS.n3391 VSS.n3390 3.4105
R20771 VSS.n3907 VSS.n3906 3.4105
R20772 VSS.n3906 VSS.n3905 3.4105
R20773 VSS.n3871 VSS.n3870 3.4105
R20774 VSS.n3890 VSS.n3889 3.4105
R20775 VSS.n3855 VSS.n3854 3.4105
R20776 VSS.n3854 VSS.n3853 3.4105
R20777 VSS.n3856 VSS.n3409 3.4105
R20778 VSS.n3859 VSS.n3404 3.4105
R20779 VSS.n3828 VSS.n3827 3.4105
R20780 VSS.n3828 VSS.n3427 3.4105
R20781 VSS.n3423 VSS.n3410 3.4105
R20782 VSS.n3835 VSS.n3423 3.4105
R20783 VSS.n3774 VSS.n3773 3.4105
R20784 VSS.n3774 VSS.n3437 3.4105
R20785 VSS.n3751 VSS.n3750 3.4105
R20786 VSS.n3772 VSS.n3771 3.4105
R20787 VSS.n3771 VSS.n3770 3.4105
R20788 VSS.n3741 VSS.n3467 3.4105
R20789 VSS.n3467 VSS.n3466 3.4105
R20790 VSS.n3743 VSS.n3742 3.4105
R20791 VSS.n3749 VSS.n3748 3.4105
R20792 VSS.n3748 VSS.n3747 3.4105
R20793 VSS.n3724 VSS.n3723 3.4105
R20794 VSS.n3724 VSS.n3481 3.4105
R20795 VSS.n3720 VSS.n3469 3.4105
R20796 VSS.n3740 VSS.n3739 3.4105
R20797 VSS.n3739 VSS.n3738 3.4105
R20798 VSS.n3703 VSS.n3702 3.4105
R20799 VSS.n3703 VSS.n3497 3.4105
R20800 VSS.n3719 VSS.n3718 3.4105
R20801 VSS.n3701 VSS.n3700 3.4105
R20802 VSS.n3700 VSS.n3699 3.4105
R20803 VSS.n3815 VSS.n3434 3.4105
R20804 VSS.n3789 VSS.n3434 3.4105
R20805 VSS.n3431 VSS.n3430 3.4105
R20806 VSS.n3825 VSS.n3824 3.4105
R20807 VSS.n3824 VSS.n3823 3.4105
R20808 VSS.n3667 VSS.n3666 3.4105
R20809 VSS.n3667 VSS.n3512 3.4105
R20810 VSS.n3660 VSS.n3659 3.4105
R20811 VSS.n3665 VSS.n3664 3.4105
R20812 VSS.n3664 VSS.n3663 3.4105
R20813 VSS.n3640 VSS.n3639 3.4105
R20814 VSS.n3640 VSS.n3552 3.4105
R20815 VSS.n3638 VSS.n3637 3.4105
R20816 VSS.n3658 VSS.n3657 3.4105
R20817 VSS.n3657 VSS.n3656 3.4105
R20818 VSS.n3627 VSS.n3558 3.4105
R20819 VSS.n3558 VSS.n3557 3.4105
R20820 VSS.n3556 VSS.n3555 3.4105
R20821 VSS.n3635 VSS.n3634 3.4105
R20822 VSS.n3634 VSS.n3550 3.4105
R20823 VSS.n3605 VSS.n3604 3.4105
R20824 VSS.n3605 VSS.n3577 3.4105
R20825 VSS.n3626 VSS.n3625 3.4105
R20826 VSS.n3603 VSS.n3602 3.4105
R20827 VSS.n3602 VSS.n3601 3.4105
R20828 VSS.n4519 VSS.n3970 3.4105
R20829 VSS.n4525 VSS.n3970 3.4105
R20830 VSS.n4521 VSS.n4520 3.4105
R20831 VSS.n4545 VSS.n4544 3.4105
R20832 VSS.n4544 VSS.n4543 3.4105
R20833 VSS.n4502 VSS.n4500 3.4105
R20834 VSS.n4502 VSS.n4501 3.4105
R20835 VSS.n4518 VSS.n4517 3.4105
R20836 VSS.n4517 VSS.n4516 3.4105
R20837 VSS.n4480 VSS.n4479 3.4105
R20838 VSS.n4479 VSS.n4478 3.4105
R20839 VSS.n3983 VSS.n3982 3.4105
R20840 VSS.n4499 VSS.n4498 3.4105
R20841 VSS.n4498 VSS.n4497 3.4105
R20842 VSS.n4463 VSS.n4462 3.4105
R20843 VSS.n4482 VSS.n4481 3.4105
R20844 VSS.n4447 VSS.n4446 3.4105
R20845 VSS.n4446 VSS.n4445 3.4105
R20846 VSS.n4448 VSS.n4001 3.4105
R20847 VSS.n4451 VSS.n3996 3.4105
R20848 VSS.n4420 VSS.n4419 3.4105
R20849 VSS.n4420 VSS.n4019 3.4105
R20850 VSS.n4015 VSS.n4002 3.4105
R20851 VSS.n4427 VSS.n4015 3.4105
R20852 VSS.n4366 VSS.n4365 3.4105
R20853 VSS.n4366 VSS.n4029 3.4105
R20854 VSS.n4343 VSS.n4342 3.4105
R20855 VSS.n4364 VSS.n4363 3.4105
R20856 VSS.n4363 VSS.n4362 3.4105
R20857 VSS.n4333 VSS.n4059 3.4105
R20858 VSS.n4059 VSS.n4058 3.4105
R20859 VSS.n4335 VSS.n4334 3.4105
R20860 VSS.n4341 VSS.n4340 3.4105
R20861 VSS.n4340 VSS.n4339 3.4105
R20862 VSS.n4316 VSS.n4315 3.4105
R20863 VSS.n4316 VSS.n4073 3.4105
R20864 VSS.n4312 VSS.n4061 3.4105
R20865 VSS.n4332 VSS.n4331 3.4105
R20866 VSS.n4331 VSS.n4330 3.4105
R20867 VSS.n4295 VSS.n4294 3.4105
R20868 VSS.n4295 VSS.n4089 3.4105
R20869 VSS.n4311 VSS.n4310 3.4105
R20870 VSS.n4293 VSS.n4292 3.4105
R20871 VSS.n4292 VSS.n4291 3.4105
R20872 VSS.n4407 VSS.n4026 3.4105
R20873 VSS.n4381 VSS.n4026 3.4105
R20874 VSS.n4023 VSS.n4022 3.4105
R20875 VSS.n4417 VSS.n4416 3.4105
R20876 VSS.n4416 VSS.n4415 3.4105
R20877 VSS.n4259 VSS.n4258 3.4105
R20878 VSS.n4259 VSS.n4104 3.4105
R20879 VSS.n4252 VSS.n4251 3.4105
R20880 VSS.n4257 VSS.n4256 3.4105
R20881 VSS.n4256 VSS.n4255 3.4105
R20882 VSS.n4232 VSS.n4231 3.4105
R20883 VSS.n4232 VSS.n4144 3.4105
R20884 VSS.n4230 VSS.n4229 3.4105
R20885 VSS.n4250 VSS.n4249 3.4105
R20886 VSS.n4249 VSS.n4248 3.4105
R20887 VSS.n4219 VSS.n4150 3.4105
R20888 VSS.n4150 VSS.n4149 3.4105
R20889 VSS.n4148 VSS.n4147 3.4105
R20890 VSS.n4227 VSS.n4226 3.4105
R20891 VSS.n4226 VSS.n4142 3.4105
R20892 VSS.n4197 VSS.n4196 3.4105
R20893 VSS.n4197 VSS.n4169 3.4105
R20894 VSS.n4218 VSS.n4217 3.4105
R20895 VSS.n4195 VSS.n4194 3.4105
R20896 VSS.n4194 VSS.n4193 3.4105
R20897 VSS.n5111 VSS.n4562 3.4105
R20898 VSS.n5117 VSS.n4562 3.4105
R20899 VSS.n5113 VSS.n5112 3.4105
R20900 VSS.n5137 VSS.n5136 3.4105
R20901 VSS.n5136 VSS.n5135 3.4105
R20902 VSS.n5094 VSS.n5092 3.4105
R20903 VSS.n5094 VSS.n5093 3.4105
R20904 VSS.n5110 VSS.n5109 3.4105
R20905 VSS.n5109 VSS.n5108 3.4105
R20906 VSS.n5072 VSS.n5071 3.4105
R20907 VSS.n5071 VSS.n5070 3.4105
R20908 VSS.n4575 VSS.n4574 3.4105
R20909 VSS.n5091 VSS.n5090 3.4105
R20910 VSS.n5090 VSS.n5089 3.4105
R20911 VSS.n5055 VSS.n5054 3.4105
R20912 VSS.n5074 VSS.n5073 3.4105
R20913 VSS.n5039 VSS.n5038 3.4105
R20914 VSS.n5038 VSS.n5037 3.4105
R20915 VSS.n5040 VSS.n4593 3.4105
R20916 VSS.n5043 VSS.n4588 3.4105
R20917 VSS.n5012 VSS.n5011 3.4105
R20918 VSS.n5012 VSS.n4611 3.4105
R20919 VSS.n4607 VSS.n4594 3.4105
R20920 VSS.n5019 VSS.n4607 3.4105
R20921 VSS.n4958 VSS.n4957 3.4105
R20922 VSS.n4958 VSS.n4621 3.4105
R20923 VSS.n4935 VSS.n4934 3.4105
R20924 VSS.n4956 VSS.n4955 3.4105
R20925 VSS.n4955 VSS.n4954 3.4105
R20926 VSS.n4925 VSS.n4651 3.4105
R20927 VSS.n4651 VSS.n4650 3.4105
R20928 VSS.n4927 VSS.n4926 3.4105
R20929 VSS.n4933 VSS.n4932 3.4105
R20930 VSS.n4932 VSS.n4931 3.4105
R20931 VSS.n4908 VSS.n4907 3.4105
R20932 VSS.n4908 VSS.n4665 3.4105
R20933 VSS.n4904 VSS.n4653 3.4105
R20934 VSS.n4924 VSS.n4923 3.4105
R20935 VSS.n4923 VSS.n4922 3.4105
R20936 VSS.n4887 VSS.n4886 3.4105
R20937 VSS.n4887 VSS.n4681 3.4105
R20938 VSS.n4903 VSS.n4902 3.4105
R20939 VSS.n4885 VSS.n4884 3.4105
R20940 VSS.n4884 VSS.n4883 3.4105
R20941 VSS.n4999 VSS.n4618 3.4105
R20942 VSS.n4973 VSS.n4618 3.4105
R20943 VSS.n4615 VSS.n4614 3.4105
R20944 VSS.n5009 VSS.n5008 3.4105
R20945 VSS.n5008 VSS.n5007 3.4105
R20946 VSS.n4851 VSS.n4850 3.4105
R20947 VSS.n4851 VSS.n4696 3.4105
R20948 VSS.n4844 VSS.n4843 3.4105
R20949 VSS.n4849 VSS.n4848 3.4105
R20950 VSS.n4848 VSS.n4847 3.4105
R20951 VSS.n4824 VSS.n4823 3.4105
R20952 VSS.n4824 VSS.n4736 3.4105
R20953 VSS.n4822 VSS.n4821 3.4105
R20954 VSS.n4842 VSS.n4841 3.4105
R20955 VSS.n4841 VSS.n4840 3.4105
R20956 VSS.n4811 VSS.n4742 3.4105
R20957 VSS.n4742 VSS.n4741 3.4105
R20958 VSS.n4740 VSS.n4739 3.4105
R20959 VSS.n4819 VSS.n4818 3.4105
R20960 VSS.n4818 VSS.n4734 3.4105
R20961 VSS.n4789 VSS.n4788 3.4105
R20962 VSS.n4789 VSS.n4761 3.4105
R20963 VSS.n4810 VSS.n4809 3.4105
R20964 VSS.n4787 VSS.n4786 3.4105
R20965 VSS.n4786 VSS.n4785 3.4105
R20966 VSS.n5703 VSS.n5154 3.4105
R20967 VSS.n5709 VSS.n5154 3.4105
R20968 VSS.n5705 VSS.n5704 3.4105
R20969 VSS.n5729 VSS.n5728 3.4105
R20970 VSS.n5728 VSS.n5727 3.4105
R20971 VSS.n5686 VSS.n5684 3.4105
R20972 VSS.n5686 VSS.n5685 3.4105
R20973 VSS.n5702 VSS.n5701 3.4105
R20974 VSS.n5701 VSS.n5700 3.4105
R20975 VSS.n5664 VSS.n5663 3.4105
R20976 VSS.n5663 VSS.n5662 3.4105
R20977 VSS.n5167 VSS.n5166 3.4105
R20978 VSS.n5683 VSS.n5682 3.4105
R20979 VSS.n5682 VSS.n5681 3.4105
R20980 VSS.n5647 VSS.n5646 3.4105
R20981 VSS.n5666 VSS.n5665 3.4105
R20982 VSS.n5631 VSS.n5630 3.4105
R20983 VSS.n5630 VSS.n5629 3.4105
R20984 VSS.n5632 VSS.n5185 3.4105
R20985 VSS.n5635 VSS.n5180 3.4105
R20986 VSS.n5604 VSS.n5603 3.4105
R20987 VSS.n5604 VSS.n5203 3.4105
R20988 VSS.n5199 VSS.n5186 3.4105
R20989 VSS.n5611 VSS.n5199 3.4105
R20990 VSS.n5550 VSS.n5549 3.4105
R20991 VSS.n5550 VSS.n5213 3.4105
R20992 VSS.n5527 VSS.n5526 3.4105
R20993 VSS.n5548 VSS.n5547 3.4105
R20994 VSS.n5547 VSS.n5546 3.4105
R20995 VSS.n5517 VSS.n5243 3.4105
R20996 VSS.n5243 VSS.n5242 3.4105
R20997 VSS.n5519 VSS.n5518 3.4105
R20998 VSS.n5525 VSS.n5524 3.4105
R20999 VSS.n5524 VSS.n5523 3.4105
R21000 VSS.n5500 VSS.n5499 3.4105
R21001 VSS.n5500 VSS.n5257 3.4105
R21002 VSS.n5496 VSS.n5245 3.4105
R21003 VSS.n5516 VSS.n5515 3.4105
R21004 VSS.n5515 VSS.n5514 3.4105
R21005 VSS.n5479 VSS.n5478 3.4105
R21006 VSS.n5479 VSS.n5273 3.4105
R21007 VSS.n5495 VSS.n5494 3.4105
R21008 VSS.n5477 VSS.n5476 3.4105
R21009 VSS.n5476 VSS.n5475 3.4105
R21010 VSS.n5591 VSS.n5210 3.4105
R21011 VSS.n5565 VSS.n5210 3.4105
R21012 VSS.n5207 VSS.n5206 3.4105
R21013 VSS.n5601 VSS.n5600 3.4105
R21014 VSS.n5600 VSS.n5599 3.4105
R21015 VSS.n5443 VSS.n5442 3.4105
R21016 VSS.n5443 VSS.n5288 3.4105
R21017 VSS.n5436 VSS.n5435 3.4105
R21018 VSS.n5441 VSS.n5440 3.4105
R21019 VSS.n5440 VSS.n5439 3.4105
R21020 VSS.n5416 VSS.n5415 3.4105
R21021 VSS.n5416 VSS.n5328 3.4105
R21022 VSS.n5414 VSS.n5413 3.4105
R21023 VSS.n5434 VSS.n5433 3.4105
R21024 VSS.n5433 VSS.n5432 3.4105
R21025 VSS.n5403 VSS.n5334 3.4105
R21026 VSS.n5334 VSS.n5333 3.4105
R21027 VSS.n5332 VSS.n5331 3.4105
R21028 VSS.n5411 VSS.n5410 3.4105
R21029 VSS.n5410 VSS.n5326 3.4105
R21030 VSS.n5381 VSS.n5380 3.4105
R21031 VSS.n5381 VSS.n5353 3.4105
R21032 VSS.n5402 VSS.n5401 3.4105
R21033 VSS.n5379 VSS.n5378 3.4105
R21034 VSS.n5378 VSS.n5377 3.4105
R21035 VSS.n6295 VSS.n5746 3.4105
R21036 VSS.n6301 VSS.n5746 3.4105
R21037 VSS.n6297 VSS.n6296 3.4105
R21038 VSS.n6321 VSS.n6320 3.4105
R21039 VSS.n6320 VSS.n6319 3.4105
R21040 VSS.n6278 VSS.n6276 3.4105
R21041 VSS.n6278 VSS.n6277 3.4105
R21042 VSS.n6294 VSS.n6293 3.4105
R21043 VSS.n6293 VSS.n6292 3.4105
R21044 VSS.n6256 VSS.n6255 3.4105
R21045 VSS.n6255 VSS.n6254 3.4105
R21046 VSS.n5759 VSS.n5758 3.4105
R21047 VSS.n6275 VSS.n6274 3.4105
R21048 VSS.n6274 VSS.n6273 3.4105
R21049 VSS.n6239 VSS.n6238 3.4105
R21050 VSS.n6258 VSS.n6257 3.4105
R21051 VSS.n6223 VSS.n6222 3.4105
R21052 VSS.n6222 VSS.n6221 3.4105
R21053 VSS.n6224 VSS.n5777 3.4105
R21054 VSS.n6227 VSS.n5772 3.4105
R21055 VSS.n6196 VSS.n6195 3.4105
R21056 VSS.n6196 VSS.n5795 3.4105
R21057 VSS.n5791 VSS.n5778 3.4105
R21058 VSS.n6203 VSS.n5791 3.4105
R21059 VSS.n6142 VSS.n6141 3.4105
R21060 VSS.n6142 VSS.n5805 3.4105
R21061 VSS.n6119 VSS.n6118 3.4105
R21062 VSS.n6140 VSS.n6139 3.4105
R21063 VSS.n6139 VSS.n6138 3.4105
R21064 VSS.n6109 VSS.n5835 3.4105
R21065 VSS.n5835 VSS.n5834 3.4105
R21066 VSS.n6111 VSS.n6110 3.4105
R21067 VSS.n6117 VSS.n6116 3.4105
R21068 VSS.n6116 VSS.n6115 3.4105
R21069 VSS.n6092 VSS.n6091 3.4105
R21070 VSS.n6092 VSS.n5849 3.4105
R21071 VSS.n6088 VSS.n5837 3.4105
R21072 VSS.n6108 VSS.n6107 3.4105
R21073 VSS.n6107 VSS.n6106 3.4105
R21074 VSS.n6071 VSS.n6070 3.4105
R21075 VSS.n6071 VSS.n5865 3.4105
R21076 VSS.n6087 VSS.n6086 3.4105
R21077 VSS.n6069 VSS.n6068 3.4105
R21078 VSS.n6068 VSS.n6067 3.4105
R21079 VSS.n6183 VSS.n5802 3.4105
R21080 VSS.n6157 VSS.n5802 3.4105
R21081 VSS.n5799 VSS.n5798 3.4105
R21082 VSS.n6193 VSS.n6192 3.4105
R21083 VSS.n6192 VSS.n6191 3.4105
R21084 VSS.n6035 VSS.n6034 3.4105
R21085 VSS.n6035 VSS.n5880 3.4105
R21086 VSS.n6028 VSS.n6027 3.4105
R21087 VSS.n6033 VSS.n6032 3.4105
R21088 VSS.n6032 VSS.n6031 3.4105
R21089 VSS.n6008 VSS.n6007 3.4105
R21090 VSS.n6008 VSS.n5920 3.4105
R21091 VSS.n6006 VSS.n6005 3.4105
R21092 VSS.n6026 VSS.n6025 3.4105
R21093 VSS.n6025 VSS.n6024 3.4105
R21094 VSS.n5995 VSS.n5926 3.4105
R21095 VSS.n5926 VSS.n5925 3.4105
R21096 VSS.n5924 VSS.n5923 3.4105
R21097 VSS.n6003 VSS.n6002 3.4105
R21098 VSS.n6002 VSS.n5918 3.4105
R21099 VSS.n5973 VSS.n5972 3.4105
R21100 VSS.n5973 VSS.n5945 3.4105
R21101 VSS.n5994 VSS.n5993 3.4105
R21102 VSS.n5971 VSS.n5970 3.4105
R21103 VSS.n5970 VSS.n5969 3.4105
R21104 VSS.n6887 VSS.n6338 3.4105
R21105 VSS.n6893 VSS.n6338 3.4105
R21106 VSS.n6889 VSS.n6888 3.4105
R21107 VSS.n6913 VSS.n6912 3.4105
R21108 VSS.n6912 VSS.n6911 3.4105
R21109 VSS.n6870 VSS.n6868 3.4105
R21110 VSS.n6870 VSS.n6869 3.4105
R21111 VSS.n6886 VSS.n6885 3.4105
R21112 VSS.n6885 VSS.n6884 3.4105
R21113 VSS.n6848 VSS.n6847 3.4105
R21114 VSS.n6847 VSS.n6846 3.4105
R21115 VSS.n6351 VSS.n6350 3.4105
R21116 VSS.n6867 VSS.n6866 3.4105
R21117 VSS.n6866 VSS.n6865 3.4105
R21118 VSS.n6831 VSS.n6830 3.4105
R21119 VSS.n6850 VSS.n6849 3.4105
R21120 VSS.n6815 VSS.n6814 3.4105
R21121 VSS.n6814 VSS.n6813 3.4105
R21122 VSS.n6816 VSS.n6369 3.4105
R21123 VSS.n6819 VSS.n6364 3.4105
R21124 VSS.n6788 VSS.n6787 3.4105
R21125 VSS.n6788 VSS.n6387 3.4105
R21126 VSS.n6383 VSS.n6370 3.4105
R21127 VSS.n6795 VSS.n6383 3.4105
R21128 VSS.n6734 VSS.n6733 3.4105
R21129 VSS.n6734 VSS.n6397 3.4105
R21130 VSS.n6711 VSS.n6710 3.4105
R21131 VSS.n6732 VSS.n6731 3.4105
R21132 VSS.n6731 VSS.n6730 3.4105
R21133 VSS.n6701 VSS.n6427 3.4105
R21134 VSS.n6427 VSS.n6426 3.4105
R21135 VSS.n6703 VSS.n6702 3.4105
R21136 VSS.n6709 VSS.n6708 3.4105
R21137 VSS.n6708 VSS.n6707 3.4105
R21138 VSS.n6684 VSS.n6683 3.4105
R21139 VSS.n6684 VSS.n6441 3.4105
R21140 VSS.n6680 VSS.n6429 3.4105
R21141 VSS.n6700 VSS.n6699 3.4105
R21142 VSS.n6699 VSS.n6698 3.4105
R21143 VSS.n6663 VSS.n6662 3.4105
R21144 VSS.n6663 VSS.n6457 3.4105
R21145 VSS.n6679 VSS.n6678 3.4105
R21146 VSS.n6661 VSS.n6660 3.4105
R21147 VSS.n6660 VSS.n6659 3.4105
R21148 VSS.n6775 VSS.n6394 3.4105
R21149 VSS.n6749 VSS.n6394 3.4105
R21150 VSS.n6391 VSS.n6390 3.4105
R21151 VSS.n6785 VSS.n6784 3.4105
R21152 VSS.n6784 VSS.n6783 3.4105
R21153 VSS.n6627 VSS.n6626 3.4105
R21154 VSS.n6627 VSS.n6472 3.4105
R21155 VSS.n6620 VSS.n6619 3.4105
R21156 VSS.n6625 VSS.n6624 3.4105
R21157 VSS.n6624 VSS.n6623 3.4105
R21158 VSS.n6600 VSS.n6599 3.4105
R21159 VSS.n6600 VSS.n6512 3.4105
R21160 VSS.n6598 VSS.n6597 3.4105
R21161 VSS.n6618 VSS.n6617 3.4105
R21162 VSS.n6617 VSS.n6616 3.4105
R21163 VSS.n6587 VSS.n6518 3.4105
R21164 VSS.n6518 VSS.n6517 3.4105
R21165 VSS.n6516 VSS.n6515 3.4105
R21166 VSS.n6595 VSS.n6594 3.4105
R21167 VSS.n6594 VSS.n6510 3.4105
R21168 VSS.n6565 VSS.n6564 3.4105
R21169 VSS.n6565 VSS.n6537 3.4105
R21170 VSS.n6586 VSS.n6585 3.4105
R21171 VSS.n6563 VSS.n6562 3.4105
R21172 VSS.n6562 VSS.n6561 3.4105
R21173 VSS.n2766 VSS.n2720 3.4105
R21174 VSS.n2766 VSS.n2765 3.4105
R21175 VSS.n2769 VSS.n2768 3.4105
R21176 VSS.n6919 VSS.n6918 3.4105
R21177 VSS.n6920 VSS.n6919 3.4105
R21178 VSS.n6937 VSS.n6936 3.4105
R21179 VSS.n6938 VSS.n6937 3.4105
R21180 VSS.n6934 VSS.n6933 3.4105
R21181 VSS.n6933 VSS.n6932 3.4105
R21182 VSS.n6952 VSS.n6951 3.4105
R21183 VSS.n6951 VSS.n6950 3.4105
R21184 VSS.n2718 VSS.n2717 3.4105
R21185 VSS.n2719 VSS.n2711 3.4105
R21186 VSS.n2711 VSS.n2707 3.4105
R21187 VSS.n2701 VSS.n2700 3.4105
R21188 VSS.n6954 VSS.n6953 3.4105
R21189 VSS.n6969 VSS.n2669 3.4105
R21190 VSS.n6969 VSS.n6968 3.4105
R21191 VSS.n2686 VSS.n2662 3.4105
R21192 VSS.n2689 VSS.n2682 3.4105
R21193 VSS.n6985 VSS.n2652 3.4105
R21194 VSS.n6985 VSS.n6984 3.4105
R21195 VSS.n2668 VSS.n2667 3.4105
R21196 VSS.n2667 VSS.n2666 3.4105
R21197 VSS.n7008 VSS.n7007 3.4105
R21198 VSS.n7007 VSS.n7006 3.4105
R21199 VSS.n7015 VSS.n7014 3.4105
R21200 VSS.n7010 VSS.n7009 3.4105
R21201 VSS.n7011 VSS.n7010 3.4105
R21202 VSS.n7023 VSS.n7022 3.4105
R21203 VSS.n7022 VSS.n7021 3.4105
R21204 VSS.n2514 VSS.n2510 3.4105
R21205 VSS.n7017 VSS.n7016 3.4105
R21206 VSS.n7017 VSS.n2513 3.4105
R21207 VSS.n7031 VSS.n7030 3.4105
R21208 VSS.n7030 VSS.n7029 3.4105
R21209 VSS.n2509 VSS.n2507 3.4105
R21210 VSS.n7025 VSS.n7024 3.4105
R21211 VSS.n7025 VSS.n2505 3.4105
R21212 VSS.n7038 VSS.n7037 3.4105
R21213 VSS.n7037 VSS.n7036 3.4105
R21214 VSS.n7033 VSS.n7032 3.4105
R21215 VSS.n7039 VSS.n2494 3.4105
R21216 VSS.n2494 VSS.n2313 3.4105
R21217 VSS.n2643 VSS.n2641 3.4105
R21218 VSS.n2641 VSS.n2640 3.4105
R21219 VSS.n2635 VSS.n2634 3.4105
R21220 VSS.n2651 VSS.n2650 3.4105
R21221 VSS.n2650 VSS.n2649 3.4105
R21222 VSS.n2471 VSS.n2470 3.4105
R21223 VSS.n2471 VSS.n2316 3.4105
R21224 VSS.n2464 VSS.n2463 3.4105
R21225 VSS.n2469 VSS.n2468 3.4105
R21226 VSS.n2468 VSS.n2467 3.4105
R21227 VSS.n2444 VSS.n2443 3.4105
R21228 VSS.n2444 VSS.n2356 3.4105
R21229 VSS.n2442 VSS.n2441 3.4105
R21230 VSS.n2462 VSS.n2461 3.4105
R21231 VSS.n2461 VSS.n2460 3.4105
R21232 VSS.n2431 VSS.n2362 3.4105
R21233 VSS.n2362 VSS.n2361 3.4105
R21234 VSS.n2360 VSS.n2359 3.4105
R21235 VSS.n2439 VSS.n2438 3.4105
R21236 VSS.n2438 VSS.n2354 3.4105
R21237 VSS.n2409 VSS.n2408 3.4105
R21238 VSS.n2409 VSS.n2381 3.4105
R21239 VSS.n2430 VSS.n2429 3.4105
R21240 VSS.n2407 VSS.n2406 3.4105
R21241 VSS.n2406 VSS.n2405 3.4105
R21242 VSS.n3335 VSS.n2785 3.4105
R21243 VSS.n3341 VSS.n2785 3.4105
R21244 VSS.n3337 VSS.n3336 3.4105
R21245 VSS.n3361 VSS.n3360 3.4105
R21246 VSS.n3360 VSS.n3359 3.4105
R21247 VSS.n3318 VSS.n3316 3.4105
R21248 VSS.n3318 VSS.n3317 3.4105
R21249 VSS.n3334 VSS.n3333 3.4105
R21250 VSS.n3333 VSS.n3332 3.4105
R21251 VSS.n3296 VSS.n3295 3.4105
R21252 VSS.n3295 VSS.n3294 3.4105
R21253 VSS.n2798 VSS.n2797 3.4105
R21254 VSS.n3315 VSS.n3314 3.4105
R21255 VSS.n3314 VSS.n3313 3.4105
R21256 VSS.n3279 VSS.n3278 3.4105
R21257 VSS.n3298 VSS.n3297 3.4105
R21258 VSS.n3263 VSS.n3262 3.4105
R21259 VSS.n3262 VSS.n3261 3.4105
R21260 VSS.n3264 VSS.n2816 3.4105
R21261 VSS.n3267 VSS.n2811 3.4105
R21262 VSS.n3236 VSS.n3235 3.4105
R21263 VSS.n3236 VSS.n2834 3.4105
R21264 VSS.n2830 VSS.n2817 3.4105
R21265 VSS.n3243 VSS.n2830 3.4105
R21266 VSS.n3182 VSS.n3181 3.4105
R21267 VSS.n3182 VSS.n2844 3.4105
R21268 VSS.n3159 VSS.n3158 3.4105
R21269 VSS.n3180 VSS.n3179 3.4105
R21270 VSS.n3179 VSS.n3178 3.4105
R21271 VSS.n3149 VSS.n2874 3.4105
R21272 VSS.n2874 VSS.n2873 3.4105
R21273 VSS.n3151 VSS.n3150 3.4105
R21274 VSS.n3157 VSS.n3156 3.4105
R21275 VSS.n3156 VSS.n3155 3.4105
R21276 VSS.n3132 VSS.n3131 3.4105
R21277 VSS.n3132 VSS.n2888 3.4105
R21278 VSS.n3128 VSS.n2876 3.4105
R21279 VSS.n3148 VSS.n3147 3.4105
R21280 VSS.n3147 VSS.n3146 3.4105
R21281 VSS.n3111 VSS.n3110 3.4105
R21282 VSS.n3111 VSS.n2904 3.4105
R21283 VSS.n3127 VSS.n3126 3.4105
R21284 VSS.n3109 VSS.n3108 3.4105
R21285 VSS.n3108 VSS.n3107 3.4105
R21286 VSS.n3223 VSS.n2841 3.4105
R21287 VSS.n3197 VSS.n2841 3.4105
R21288 VSS.n2838 VSS.n2837 3.4105
R21289 VSS.n3233 VSS.n3232 3.4105
R21290 VSS.n3232 VSS.n3231 3.4105
R21291 VSS.n3078 VSS.n3077 3.4105
R21292 VSS.n3078 VSS.n2919 3.4105
R21293 VSS.n3054 VSS.n3053 3.4105
R21294 VSS.n3076 VSS.n3075 3.4105
R21295 VSS.n3075 VSS.n3074 3.4105
R21296 VSS.n3044 VSS.n2949 3.4105
R21297 VSS.n2949 VSS.n2948 3.4105
R21298 VSS.n3046 VSS.n3045 3.4105
R21299 VSS.n3052 VSS.n3051 3.4105
R21300 VSS.n3051 VSS.n3050 3.4105
R21301 VSS.n3027 VSS.n3026 3.4105
R21302 VSS.n3027 VSS.n2965 3.4105
R21303 VSS.n3023 VSS.n2951 3.4105
R21304 VSS.n3043 VSS.n3042 3.4105
R21305 VSS.n3042 VSS.n3041 3.4105
R21306 VSS.n3006 VSS.n3005 3.4105
R21307 VSS.n3006 VSS.n2979 3.4105
R21308 VSS.n3022 VSS.n3021 3.4105
R21309 VSS.n3004 VSS.n3003 3.4105
R21310 VSS.n3003 VSS.n3002 3.4105
R21311 VSS.n9295 VSS.n52 3.4105
R21312 VSS.n9301 VSS.n52 3.4105
R21313 VSS.n9297 VSS.n9296 3.4105
R21314 VSS.n9321 VSS.n9320 3.4105
R21315 VSS.n9320 VSS.n9319 3.4105
R21316 VSS.n9278 VSS.n9276 3.4105
R21317 VSS.n9278 VSS.n9277 3.4105
R21318 VSS.n9294 VSS.n9293 3.4105
R21319 VSS.n9293 VSS.n9292 3.4105
R21320 VSS.n9256 VSS.n9255 3.4105
R21321 VSS.n9255 VSS.n9254 3.4105
R21322 VSS.n65 VSS.n64 3.4105
R21323 VSS.n9275 VSS.n9274 3.4105
R21324 VSS.n9274 VSS.n9273 3.4105
R21325 VSS.n9239 VSS.n9238 3.4105
R21326 VSS.n9258 VSS.n9257 3.4105
R21327 VSS.n9223 VSS.n9222 3.4105
R21328 VSS.n9222 VSS.n9221 3.4105
R21329 VSS.n9224 VSS.n83 3.4105
R21330 VSS.n9227 VSS.n78 3.4105
R21331 VSS.n9196 VSS.n9195 3.4105
R21332 VSS.n9196 VSS.n101 3.4105
R21333 VSS.n97 VSS.n84 3.4105
R21334 VSS.n9203 VSS.n97 3.4105
R21335 VSS.n9142 VSS.n9141 3.4105
R21336 VSS.n9142 VSS.n111 3.4105
R21337 VSS.n9119 VSS.n9118 3.4105
R21338 VSS.n9140 VSS.n9139 3.4105
R21339 VSS.n9139 VSS.n9138 3.4105
R21340 VSS.n9109 VSS.n141 3.4105
R21341 VSS.n141 VSS.n140 3.4105
R21342 VSS.n9111 VSS.n9110 3.4105
R21343 VSS.n9117 VSS.n9116 3.4105
R21344 VSS.n9116 VSS.n9115 3.4105
R21345 VSS.n9092 VSS.n9091 3.4105
R21346 VSS.n9092 VSS.n155 3.4105
R21347 VSS.n9088 VSS.n143 3.4105
R21348 VSS.n9108 VSS.n9107 3.4105
R21349 VSS.n9107 VSS.n9106 3.4105
R21350 VSS.n9071 VSS.n9070 3.4105
R21351 VSS.n9071 VSS.n171 3.4105
R21352 VSS.n9087 VSS.n9086 3.4105
R21353 VSS.n9069 VSS.n9068 3.4105
R21354 VSS.n9068 VSS.n9067 3.4105
R21355 VSS.n9183 VSS.n108 3.4105
R21356 VSS.n9157 VSS.n108 3.4105
R21357 VSS.n105 VSS.n104 3.4105
R21358 VSS.n9193 VSS.n9192 3.4105
R21359 VSS.n9192 VSS.n9191 3.4105
R21360 VSS.n399 VSS.n398 3.4105
R21361 VSS.n398 VSS.n179 3.4105
R21362 VSS.n406 VSS.n405 3.4105
R21363 VSS.n401 VSS.n400 3.4105
R21364 VSS.n402 VSS.n401 3.4105
R21365 VSS.n414 VSS.n413 3.4105
R21366 VSS.n413 VSS.n412 3.4105
R21367 VSS.n298 VSS.n293 3.4105
R21368 VSS.n408 VSS.n407 3.4105
R21369 VSS.n408 VSS.n297 3.4105
R21370 VSS.n422 VSS.n421 3.4105
R21371 VSS.n421 VSS.n420 3.4105
R21372 VSS.n292 VSS.n290 3.4105
R21373 VSS.n416 VSS.n415 3.4105
R21374 VSS.n416 VSS.n288 3.4105
R21375 VSS.n429 VSS.n428 3.4105
R21376 VSS.n428 VSS.n427 3.4105
R21377 VSS.n424 VSS.n423 3.4105
R21378 VSS.n430 VSS.n277 3.4105
R21379 VSS.n277 VSS.n275 3.4105
R21380 VSS.n718 VSS.n717 3.4105
R21381 VSS.n756 VSS.n755 3.4105
R21382 VSS.n757 VSS.n756 3.4105
R21383 VSS.n753 VSS.n752 3.4105
R21384 VSS.n752 VSS.n751 3.4105
R21385 VSS.n771 VSS.n770 3.4105
R21386 VSS.n770 VSS.n769 3.4105
R21387 VSS.n710 VSS.n709 3.4105
R21388 VSS.n711 VSS.n703 3.4105
R21389 VSS.n703 VSS.n699 3.4105
R21390 VSS.n693 VSS.n692 3.4105
R21391 VSS.n773 VSS.n772 3.4105
R21392 VSS.n788 VSS.n661 3.4105
R21393 VSS.n788 VSS.n787 3.4105
R21394 VSS.n678 VSS.n654 3.4105
R21395 VSS.n681 VSS.n674 3.4105
R21396 VSS.n804 VSS.n644 3.4105
R21397 VSS.n804 VSS.n803 3.4105
R21398 VSS.n660 VSS.n659 3.4105
R21399 VSS.n659 VSS.n658 3.4105
R21400 VSS.n635 VSS.n633 3.4105
R21401 VSS.n633 VSS.n632 3.4105
R21402 VSS.n627 VSS.n626 3.4105
R21403 VSS.n643 VSS.n642 3.4105
R21404 VSS.n642 VSS.n641 3.4105
R21405 VSS.n719 VSS.n712 3.4105
R21406 VSS.n721 VSS.n719 3.4105
R21407 VSS.n827 VSS.n826 3.4105
R21408 VSS.n826 VSS.n825 3.4105
R21409 VSS.n834 VSS.n833 3.4105
R21410 VSS.n829 VSS.n828 3.4105
R21411 VSS.n830 VSS.n829 3.4105
R21412 VSS.n842 VSS.n841 3.4105
R21413 VSS.n841 VSS.n840 3.4105
R21414 VSS.n503 VSS.n499 3.4105
R21415 VSS.n836 VSS.n835 3.4105
R21416 VSS.n836 VSS.n502 3.4105
R21417 VSS.n850 VSS.n849 3.4105
R21418 VSS.n849 VSS.n848 3.4105
R21419 VSS.n498 VSS.n496 3.4105
R21420 VSS.n844 VSS.n843 3.4105
R21421 VSS.n844 VSS.n494 3.4105
R21422 VSS.n857 VSS.n856 3.4105
R21423 VSS.n856 VSS.n855 3.4105
R21424 VSS.n852 VSS.n851 3.4105
R21425 VSS.n859 VSS.n858 3.4105
R21426 VSS.n860 VSS.n859 3.4105
R21427 VSS.n9326 VSS.n9325 3.4105
R21428 VSS.n9327 VSS.n9326 3.4105
R21429 VSS.n964 VSS.n963 3.4105
R21430 VSS.n963 VSS.n962 3.4105
R21431 VSS.n971 VSS.n970 3.4105
R21432 VSS.n966 VSS.n965 3.4105
R21433 VSS.n967 VSS.n966 3.4105
R21434 VSS.n979 VSS.n978 3.4105
R21435 VSS.n978 VSS.n977 3.4105
R21436 VSS.n464 VSS.n459 3.4105
R21437 VSS.n973 VSS.n972 3.4105
R21438 VSS.n973 VSS.n463 3.4105
R21439 VSS.n987 VSS.n986 3.4105
R21440 VSS.n986 VSS.n985 3.4105
R21441 VSS.n458 VSS.n456 3.4105
R21442 VSS.n981 VSS.n980 3.4105
R21443 VSS.n981 VSS.n454 3.4105
R21444 VSS.n994 VSS.n993 3.4105
R21445 VSS.n993 VSS.n992 3.4105
R21446 VSS.n989 VSS.n988 3.4105
R21447 VSS.n995 VSS.n443 3.4105
R21448 VSS.n443 VSS.n441 3.4105
R21449 VSS.n7334 VSS.n7288 3.4105
R21450 VSS.n7334 VSS.n7333 3.4105
R21451 VSS.n7337 VSS.n7336 3.4105
R21452 VSS.n8347 VSS.n8346 3.4105
R21453 VSS.n8348 VSS.n8347 3.4105
R21454 VSS.n8365 VSS.n8364 3.4105
R21455 VSS.n8366 VSS.n8365 3.4105
R21456 VSS.n8362 VSS.n8361 3.4105
R21457 VSS.n8361 VSS.n8360 3.4105
R21458 VSS.n8380 VSS.n8379 3.4105
R21459 VSS.n8379 VSS.n8378 3.4105
R21460 VSS.n7286 VSS.n7285 3.4105
R21461 VSS.n7287 VSS.n7279 3.4105
R21462 VSS.n7279 VSS.n7275 3.4105
R21463 VSS.n7269 VSS.n7268 3.4105
R21464 VSS.n8382 VSS.n8381 3.4105
R21465 VSS.n8397 VSS.n7237 3.4105
R21466 VSS.n8397 VSS.n8396 3.4105
R21467 VSS.n7254 VSS.n7230 3.4105
R21468 VSS.n7257 VSS.n7250 3.4105
R21469 VSS.n8413 VSS.n7220 3.4105
R21470 VSS.n8413 VSS.n8412 3.4105
R21471 VSS.n7236 VSS.n7235 3.4105
R21472 VSS.n7235 VSS.n7234 3.4105
R21473 VSS.n8436 VSS.n8435 3.4105
R21474 VSS.n8435 VSS.n8434 3.4105
R21475 VSS.n8443 VSS.n8442 3.4105
R21476 VSS.n8438 VSS.n8437 3.4105
R21477 VSS.n8439 VSS.n8438 3.4105
R21478 VSS.n8451 VSS.n8450 3.4105
R21479 VSS.n8450 VSS.n8449 3.4105
R21480 VSS.n7082 VSS.n7078 3.4105
R21481 VSS.n8445 VSS.n8444 3.4105
R21482 VSS.n8445 VSS.n7081 3.4105
R21483 VSS.n8459 VSS.n8458 3.4105
R21484 VSS.n8458 VSS.n8457 3.4105
R21485 VSS.n7077 VSS.n7075 3.4105
R21486 VSS.n8453 VSS.n8452 3.4105
R21487 VSS.n8453 VSS.n7073 3.4105
R21488 VSS.n8466 VSS.n8465 3.4105
R21489 VSS.n8465 VSS.n8464 3.4105
R21490 VSS.n8461 VSS.n8460 3.4105
R21491 VSS.n8467 VSS.n7062 3.4105
R21492 VSS.n7062 VSS.n7060 3.4105
R21493 VSS.n7211 VSS.n7209 3.4105
R21494 VSS.n7209 VSS.n7208 3.4105
R21495 VSS.n7203 VSS.n7202 3.4105
R21496 VSS.n7219 VSS.n7218 3.4105
R21497 VSS.n7218 VSS.n7217 3.4105
R21498 VSS.n7123 VSS.n7122 3.29193
R21499 VSS.n7143 VSS.n7142 3.29193
R21500 VSS.n7162 VSS.n7107 3.29193
R21501 VSS.n1073 VSS.n1072 3.29193
R21502 VSS.n1091 VSS.n1090 3.29193
R21503 VSS.n1110 VSS.n1056 3.29193
R21504 VSS.n7594 VSS.n7593 3.29193
R21505 VSS.n7737 VSS.n7343 3.29193
R21506 VSS.n7479 VSS.n7469 3.29193
R21507 VSS.n7512 VSS.n7511 3.29193
R21508 VSS.n7550 VSS.n7430 3.29193
R21509 VSS.n7973 VSS.n7962 3.29193
R21510 VSS.n8000 VSS.n7956 3.29193
R21511 VSS.n7935 VSS.n7934 3.29193
R21512 VSS.n8186 VSS.n8185 3.29193
R21513 VSS.n8329 VSS.n7757 3.29193
R21514 VSS.n7893 VSS.n7883 3.29193
R21515 VSS.n8104 VSS.n8103 3.29193
R21516 VSS.n8142 VSS.n7844 3.29193
R21517 VSS.n8702 VSS.n8701 3.29193
R21518 VSS.n8722 VSS.n8721 3.29193
R21519 VSS.n8741 VSS.n8686 3.29193
R21520 VSS.n8785 VSS.n8775 3.29193
R21521 VSS.n8917 VSS.n8898 3.29193
R21522 VSS.n270 VSS.n259 3.29193
R21523 VSS.n8561 VSS.n253 3.29193
R21524 VSS.n232 VSS.n231 3.29193
R21525 VSS.n1384 VSS.n1383 3.29193
R21526 VSS.n1404 VSS.n1403 3.29193
R21527 VSS.n1423 VSS.n1368 3.29193
R21528 VSS.n1466 VSS.n1457 3.29193
R21529 VSS.n1566 VSS.n5 3.29193
R21530 VSS.n1216 VSS.n1205 3.29193
R21531 VSS.n1243 VSS.n1199 3.29193
R21532 VSS.n1178 VSS.n1177 3.29193
R21533 VSS.n1957 VSS.n1956 3.29193
R21534 VSS.n1977 VSS.n1976 3.29193
R21535 VSS.n1996 VSS.n1941 3.29193
R21536 VSS.n2039 VSS.n2030 3.29193
R21537 VSS.n2179 VSS.n2178 3.29193
R21538 VSS.n1789 VSS.n1778 3.29193
R21539 VSS.n1816 VSS.n1772 3.29193
R21540 VSS.n1751 VSS.n1750 3.29193
R21541 VSS.n3503 VSS.n3493 3.29193
R21542 VSS.n3714 VSS.n3713 3.29193
R21543 VSS.n3752 VSS.n3454 3.29193
R21544 VSS.n3796 VSS.n3795 3.29193
R21545 VSS.n3940 VSS.n3368 3.29193
R21546 VSS.n3583 VSS.n3572 3.29193
R21547 VSS.n3610 VSS.n3566 3.29193
R21548 VSS.n3545 VSS.n3544 3.29193
R21549 VSS.n4095 VSS.n4085 3.29193
R21550 VSS.n4306 VSS.n4305 3.29193
R21551 VSS.n4344 VSS.n4046 3.29193
R21552 VSS.n4388 VSS.n4387 3.29193
R21553 VSS.n4532 VSS.n3960 3.29193
R21554 VSS.n4175 VSS.n4164 3.29193
R21555 VSS.n4202 VSS.n4158 3.29193
R21556 VSS.n4137 VSS.n4136 3.29193
R21557 VSS.n4687 VSS.n4677 3.29193
R21558 VSS.n4898 VSS.n4897 3.29193
R21559 VSS.n4936 VSS.n4638 3.29193
R21560 VSS.n4980 VSS.n4979 3.29193
R21561 VSS.n5124 VSS.n4552 3.29193
R21562 VSS.n4767 VSS.n4756 3.29193
R21563 VSS.n4794 VSS.n4750 3.29193
R21564 VSS.n4729 VSS.n4728 3.29193
R21565 VSS.n5279 VSS.n5269 3.29193
R21566 VSS.n5490 VSS.n5489 3.29193
R21567 VSS.n5528 VSS.n5230 3.29193
R21568 VSS.n5572 VSS.n5571 3.29193
R21569 VSS.n5716 VSS.n5144 3.29193
R21570 VSS.n5359 VSS.n5348 3.29193
R21571 VSS.n5386 VSS.n5342 3.29193
R21572 VSS.n5321 VSS.n5320 3.29193
R21573 VSS.n5871 VSS.n5861 3.29193
R21574 VSS.n6082 VSS.n6081 3.29193
R21575 VSS.n6120 VSS.n5822 3.29193
R21576 VSS.n6164 VSS.n6163 3.29193
R21577 VSS.n6308 VSS.n5736 3.29193
R21578 VSS.n5951 VSS.n5940 3.29193
R21579 VSS.n5978 VSS.n5934 3.29193
R21580 VSS.n5913 VSS.n5912 3.29193
R21581 VSS.n6463 VSS.n6453 3.29193
R21582 VSS.n6674 VSS.n6673 3.29193
R21583 VSS.n6712 VSS.n6414 3.29193
R21584 VSS.n6756 VSS.n6755 3.29193
R21585 VSS.n6900 VSS.n6328 3.29193
R21586 VSS.n6543 VSS.n6532 3.29193
R21587 VSS.n6570 VSS.n6526 3.29193
R21588 VSS.n6505 VSS.n6504 3.29193
R21589 VSS.n2555 VSS.n2554 3.29193
R21590 VSS.n2575 VSS.n2574 3.29193
R21591 VSS.n2594 VSS.n2539 3.29193
R21592 VSS.n2637 VSS.n2628 3.29193
R21593 VSS.n6923 VSS.n6922 3.29193
R21594 VSS.n2387 VSS.n2376 3.29193
R21595 VSS.n2414 VSS.n2370 3.29193
R21596 VSS.n2349 VSS.n2348 3.29193
R21597 VSS.n2910 VSS.n2900 3.29193
R21598 VSS.n3122 VSS.n3121 3.29193
R21599 VSS.n3160 VSS.n2861 3.29193
R21600 VSS.n3204 VSS.n3203 3.29193
R21601 VSS.n3348 VSS.n2775 3.29193
R21602 VSS.n2985 VSS.n2975 3.29193
R21603 VSS.n3017 VSS.n3016 3.29193
R21604 VSS.n3055 VSS.n2936 3.29193
R21605 VSS.n186 VSS.n167 3.29193
R21606 VSS.n9082 VSS.n9081 3.29193
R21607 VSS.n9120 VSS.n128 3.29193
R21608 VSS.n9164 VSS.n9163 3.29193
R21609 VSS.n9308 VSS.n42 3.29193
R21610 VSS.n341 VSS.n340 3.29193
R21611 VSS.n349 VSS.n348 3.29193
R21612 VSS.n378 VSS.n377 3.29193
R21613 VSS.n549 VSS.n548 3.29193
R21614 VSS.n567 VSS.n566 3.29193
R21615 VSS.n586 VSS.n528 3.29193
R21616 VSS.n629 VSS.n620 3.29193
R21617 VSS.n9330 VSS.n9329 3.29193
R21618 VSS.n892 VSS.n891 3.29193
R21619 VSS.n910 VSS.n909 3.29193
R21620 VSS.n929 VSS.n875 3.29193
R21621 VSS.n7205 VSS.n7196 3.29193
R21622 VSS.n8351 VSS.n8350 3.29193
R21623 VSS.n7185 VSS.n7184 3.2005
R21624 VSS.n1134 VSS.n1133 3.2005
R21625 VSS.n7580 VSS.n7579 3.2005
R21626 VSS.n7916 VSS.n7915 3.2005
R21627 VSS.n8172 VSS.n8171 3.2005
R21628 VSS.n8764 VSS.n8763 3.2005
R21629 VSS.n213 VSS.n212 3.2005
R21630 VSS.n1446 VSS.n1445 3.2005
R21631 VSS.n1159 VSS.n1158 3.2005
R21632 VSS.n2019 VSS.n2018 3.2005
R21633 VSS.n1732 VSS.n1731 3.2005
R21634 VSS.n3782 VSS.n3781 3.2005
R21635 VSS.n3526 VSS.n3525 3.2005
R21636 VSS.n4374 VSS.n4373 3.2005
R21637 VSS.n4118 VSS.n4117 3.2005
R21638 VSS.n4966 VSS.n4965 3.2005
R21639 VSS.n4710 VSS.n4709 3.2005
R21640 VSS.n5558 VSS.n5557 3.2005
R21641 VSS.n5302 VSS.n5301 3.2005
R21642 VSS.n6150 VSS.n6149 3.2005
R21643 VSS.n5894 VSS.n5893 3.2005
R21644 VSS.n6742 VSS.n6741 3.2005
R21645 VSS.n6486 VSS.n6485 3.2005
R21646 VSS.n2617 VSS.n2616 3.2005
R21647 VSS.n2330 VSS.n2329 3.2005
R21648 VSS.n3190 VSS.n3189 3.2005
R21649 VSS.n3086 VSS.n3085 3.2005
R21650 VSS.n9150 VSS.n9149 3.2005
R21651 VSS.n388 VSS.n387 3.2005
R21652 VSS.n609 VSS.n608 3.2005
R21653 VSS.n953 VSS.n952 3.2005
R21654 VSS.n7535 VSS.n7534 3.03311
R21655 VSS.n7505 VSS.n7504 3.03311
R21656 VSS.n8127 VSS.n8126 3.03311
R21657 VSS.n8097 VSS.n8096 3.03311
R21658 VSS.n8595 VSS.n8594 3.03311
R21659 VSS.n8560 VSS.n8559 3.03311
R21660 VSS.n1372 VSS.n1341 3.03311
R21661 VSS.n1396 VSS.n1395 3.03311
R21662 VSS.n1277 VSS.n1276 3.03311
R21663 VSS.n1242 VSS.n1241 3.03311
R21664 VSS.n1945 VSS.n1914 3.03311
R21665 VSS.n1969 VSS.n1968 3.03311
R21666 VSS.n1850 VSS.n1849 3.03311
R21667 VSS.n1815 VSS.n1814 3.03311
R21668 VSS.n3737 VSS.n3736 3.03311
R21669 VSS.n3707 VSS.n3706 3.03311
R21670 VSS.n3644 VSS.n3643 3.03311
R21671 VSS.n3609 VSS.n3608 3.03311
R21672 VSS.n4329 VSS.n4328 3.03311
R21673 VSS.n4299 VSS.n4298 3.03311
R21674 VSS.n4236 VSS.n4235 3.03311
R21675 VSS.n4201 VSS.n4200 3.03311
R21676 VSS.n4921 VSS.n4920 3.03311
R21677 VSS.n4891 VSS.n4890 3.03311
R21678 VSS.n4828 VSS.n4827 3.03311
R21679 VSS.n4793 VSS.n4792 3.03311
R21680 VSS.n5513 VSS.n5512 3.03311
R21681 VSS.n5483 VSS.n5482 3.03311
R21682 VSS.n5420 VSS.n5419 3.03311
R21683 VSS.n5385 VSS.n5384 3.03311
R21684 VSS.n6105 VSS.n6104 3.03311
R21685 VSS.n6075 VSS.n6074 3.03311
R21686 VSS.n6012 VSS.n6011 3.03311
R21687 VSS.n5977 VSS.n5976 3.03311
R21688 VSS.n6697 VSS.n6696 3.03311
R21689 VSS.n6667 VSS.n6666 3.03311
R21690 VSS.n6604 VSS.n6603 3.03311
R21691 VSS.n6569 VSS.n6568 3.03311
R21692 VSS.n2543 VSS.n2512 3.03311
R21693 VSS.n2567 VSS.n2566 3.03311
R21694 VSS.n2448 VSS.n2447 3.03311
R21695 VSS.n2413 VSS.n2412 3.03311
R21696 VSS.n3145 VSS.n3144 3.03311
R21697 VSS.n3115 VSS.n3114 3.03311
R21698 VSS.n3040 VSS.n3039 3.03311
R21699 VSS.n3010 VSS.n3009 3.03311
R21700 VSS.n9105 VSS.n9104 3.03311
R21701 VSS.n9075 VSS.n9074 3.03311
R21702 VSS.n363 VSS.n362 3.03311
R21703 VSS.n330 VSS.n327 3.03311
R21704 VSS.n8690 VSS.n8659 3.03311
R21705 VSS.n8714 VSS.n8713 3.03311
R21706 VSS.n532 VSS.n501 3.03311
R21707 VSS.n559 VSS.n558 3.03311
R21708 VSS.n880 VSS.n879 3.03311
R21709 VSS.n904 VSS.n903 3.03311
R21710 VSS.n1061 VSS.n1060 3.03311
R21711 VSS.n1085 VSS.n1084 3.03311
R21712 VSS.n8034 VSS.n8033 3.03311
R21713 VSS.n7999 VSS.n7998 3.03311
R21714 VSS.n7111 VSS.n7080 3.03311
R21715 VSS.n7135 VSS.n7134 3.03311
R21716 VSS.n7149 VSS.n7114 2.81479
R21717 VSS.n7170 VSS.n7110 2.81479
R21718 VSS.n8009 VSS.n7959 2.81479
R21719 VSS.n8042 VSS.n7929 2.81479
R21720 VSS.n1097 VSS.n1064 2.81479
R21721 VSS.n1118 VSS.n1059 2.81479
R21722 VSS.n916 VSS.n883 2.81479
R21723 VSS.n937 VSS.n878 2.81479
R21724 VSS.n7528 VSS.n7454 2.81479
R21725 VSS.n7559 VSS.n7433 2.81479
R21726 VSS.n8120 VSS.n7868 2.81479
R21727 VSS.n8151 VSS.n7847 2.81479
R21728 VSS.n8728 VSS.n8693 2.81479
R21729 VSS.n8749 VSS.n8689 2.81479
R21730 VSS.n8570 VSS.n256 2.81479
R21731 VSS.n8603 VSS.n226 2.81479
R21732 VSS.n1252 VSS.n1202 2.81479
R21733 VSS.n1285 VSS.n1172 2.81479
R21734 VSS.n1410 VSS.n1375 2.81479
R21735 VSS.n1431 VSS.n1371 2.81479
R21736 VSS.n1825 VSS.n1775 2.81479
R21737 VSS.n1858 VSS.n1745 2.81479
R21738 VSS.n1983 VSS.n1948 2.81479
R21739 VSS.n2004 VSS.n1944 2.81479
R21740 VSS.n3619 VSS.n3569 2.81479
R21741 VSS.n3652 VSS.n3539 2.81479
R21742 VSS.n3730 VSS.n3478 2.81479
R21743 VSS.n3761 VSS.n3457 2.81479
R21744 VSS.n4211 VSS.n4161 2.81479
R21745 VSS.n4244 VSS.n4131 2.81479
R21746 VSS.n4322 VSS.n4070 2.81479
R21747 VSS.n4353 VSS.n4049 2.81479
R21748 VSS.n4803 VSS.n4753 2.81479
R21749 VSS.n4836 VSS.n4723 2.81479
R21750 VSS.n4914 VSS.n4662 2.81479
R21751 VSS.n4945 VSS.n4641 2.81479
R21752 VSS.n5395 VSS.n5345 2.81479
R21753 VSS.n5428 VSS.n5315 2.81479
R21754 VSS.n5506 VSS.n5254 2.81479
R21755 VSS.n5537 VSS.n5233 2.81479
R21756 VSS.n5987 VSS.n5937 2.81479
R21757 VSS.n6020 VSS.n5907 2.81479
R21758 VSS.n6098 VSS.n5846 2.81479
R21759 VSS.n6129 VSS.n5825 2.81479
R21760 VSS.n6579 VSS.n6529 2.81479
R21761 VSS.n6612 VSS.n6499 2.81479
R21762 VSS.n6690 VSS.n6438 2.81479
R21763 VSS.n6721 VSS.n6417 2.81479
R21764 VSS.n2423 VSS.n2373 2.81479
R21765 VSS.n2456 VSS.n2343 2.81479
R21766 VSS.n2581 VSS.n2546 2.81479
R21767 VSS.n2602 VSS.n2542 2.81479
R21768 VSS.n3033 VSS.n2962 2.81479
R21769 VSS.n3064 VSS.n2939 2.81479
R21770 VSS.n3138 VSS.n2885 2.81479
R21771 VSS.n3169 VSS.n2864 2.81479
R21772 VSS.n356 VSS.n323 2.81479
R21773 VSS.n369 VSS.n319 2.81479
R21774 VSS.n9098 VSS.n152 2.81479
R21775 VSS.n9129 VSS.n131 2.81479
R21776 VSS.n573 VSS.n535 2.81479
R21777 VSS.n594 VSS.n531 2.81479
R21778 VSS.n7700 VSS.n7699 2.5605
R21779 VSS.n8292 VSS.n8291 2.5605
R21780 VSS.n8954 VSS.n8953 2.5605
R21781 VSS.n1611 VSS.n1537 2.5605
R21782 VSS.n2203 VSS.n2110 2.5605
R21783 VSS.n3902 VSS.n3901 2.5605
R21784 VSS.n4494 VSS.n4493 2.5605
R21785 VSS.n5086 VSS.n5085 2.5605
R21786 VSS.n5678 VSS.n5677 2.5605
R21787 VSS.n6270 VSS.n6269 2.5605
R21788 VSS.n6862 VSS.n6861 2.5605
R21789 VSS.n6947 VSS.n2708 2.5605
R21790 VSS.n3310 VSS.n3309 2.5605
R21791 VSS.n9270 VSS.n9269 2.5605
R21792 VSS.n766 VSS.n700 2.5605
R21793 VSS.n8375 VSS.n7276 2.5605
R21794 VSS.n7649 VSS.n7648 2.46907
R21795 VSS.n8241 VSS.n8240 2.46907
R21796 VSS.n8972 VSS.n8807 2.46907
R21797 VSS.n1630 VSS.n1629 2.46907
R21798 VSS.n2222 VSS.n2221 2.46907
R21799 VSS.n3851 VSS.n3850 2.46907
R21800 VSS.n4443 VSS.n4442 2.46907
R21801 VSS.n5035 VSS.n5034 2.46907
R21802 VSS.n5627 VSS.n5626 2.46907
R21803 VSS.n6219 VSS.n6218 2.46907
R21804 VSS.n6811 VSS.n6810 2.46907
R21805 VSS.n6966 VSS.n6965 2.46907
R21806 VSS.n3259 VSS.n3258 2.46907
R21807 VSS.n9219 VSS.n9218 2.46907
R21808 VSS.n785 VSS.n784 2.46907
R21809 VSS.n8394 VSS.n8393 2.46907
R21810 VSS.n8039 VSS.t212 2.42341
R21811 VSS.n7719 VSS.n7718 2.37764
R21812 VSS.n8311 VSS.n8310 2.37764
R21813 VSS.n8944 VSS.n8883 2.37764
R21814 VSS.n1586 VSS.n1585 2.37764
R21815 VSS.n2146 VSS.n2145 2.37764
R21816 VSS.n3921 VSS.n3920 2.37764
R21817 VSS.n4513 VSS.n4512 2.37764
R21818 VSS.n5105 VSS.n5104 2.37764
R21819 VSS.n5697 VSS.n5696 2.37764
R21820 VSS.n6289 VSS.n6288 2.37764
R21821 VSS.n6881 VSS.n6880 2.37764
R21822 VSS.n2744 VSS.n2743 2.37764
R21823 VSS.n3329 VSS.n3328 2.37764
R21824 VSS.n9289 VSS.n9288 2.37764
R21825 VSS.n747 VSS.n746 2.37764
R21826 VSS.n7312 VSS.n7311 2.37764
R21827 VSS.n7631 VSS.n7396 2.28621
R21828 VSS.n8223 VSS.n7810 2.28621
R21829 VSS.n8830 VSS.n8828 2.28621
R21830 VSS.n1645 VSS.n1644 2.28621
R21831 VSS.n2237 VSS.n2236 2.28621
R21832 VSS.n3833 VSS.n3420 2.28621
R21833 VSS.n4425 VSS.n4012 2.28621
R21834 VSS.n5017 VSS.n4604 2.28621
R21835 VSS.n5609 VSS.n5196 2.28621
R21836 VSS.n6201 VSS.n5788 2.28621
R21837 VSS.n6793 VSS.n6380 2.28621
R21838 VSS.n6981 VSS.n6980 2.28621
R21839 VSS.n3241 VSS.n2827 2.28621
R21840 VSS.n9201 VSS.n94 2.28621
R21841 VSS.n800 VSS.n799 2.28621
R21842 VSS.n8409 VSS.n8408 2.28621
R21843 VSS.n8345 VSS.n8344 2.27261
R21844 VSS.n3363 VSS.n37 2.27256
R21845 VSS.n6323 VSS.n5731 2.27256
R21846 VSS.n3955 VSS.n0 2.27256
R21847 VSS.n7095 VSS.n7093 2.2505
R21848 VSS.n7161 VSS.n7084 2.2505
R21849 VSS.n7091 VSS.n7090 2.2505
R21850 VSS.n7066 VSS.n7064 2.2505
R21851 VSS.n7072 VSS.n7070 2.2505
R21852 VSS.n7127 VSS.n7126 2.2505
R21853 VSS.n1044 VSS.n1042 2.2505
R21854 VSS.n1109 VSS.n1033 2.2505
R21855 VSS.n1040 VSS.n1039 2.2505
R21856 VSS.n1014 VSS.n1012 2.2505
R21857 VSS.n1020 VSS.n1018 2.2505
R21858 VSS.n1077 VSS.n1076 2.2505
R21859 VSS.n7735 VSS.n7351 2.2505
R21860 VSS.n7682 VSS.n7672 2.2505
R21861 VSS.n7711 VSS.n7710 2.2505
R21862 VSS.n7636 VSS.n7398 2.2505
R21863 VSS.n7659 VSS.n7658 2.2505
R21864 VSS.n7661 VSS.n7381 2.2505
R21865 VSS.n7404 VSS.n7402 2.2505
R21866 VSS.n7574 VSS.n7573 2.2505
R21867 VSS.n7438 VSS.n7436 2.2505
R21868 VSS.n7567 VSS.n7425 2.2505
R21869 VSS.n7503 VSS.n7502 2.2505
R21870 VSS.n7524 VSS.n7523 2.2505
R21871 VSS.n7496 VSS.n7477 2.2505
R21872 VSS.n8059 VSS.n8058 2.2505
R21873 VSS.n8045 VSS.n7924 2.2505
R21874 VSS.n7911 VSS.n7909 2.2505
R21875 VSS.n7997 VSS.n7996 2.2505
R21876 VSS.n7954 VSS.n7953 2.2505
R21877 VSS.n7990 VSS.n7971 2.2505
R21878 VSS.n8327 VSS.n7765 2.2505
R21879 VSS.n8274 VSS.n8264 2.2505
R21880 VSS.n8303 VSS.n8302 2.2505
R21881 VSS.n8228 VSS.n7812 2.2505
R21882 VSS.n8251 VSS.n8250 2.2505
R21883 VSS.n8253 VSS.n7795 2.2505
R21884 VSS.n7818 VSS.n7816 2.2505
R21885 VSS.n8166 VSS.n8165 2.2505
R21886 VSS.n7852 VSS.n7850 2.2505
R21887 VSS.n8159 VSS.n7839 2.2505
R21888 VSS.n8095 VSS.n8094 2.2505
R21889 VSS.n8116 VSS.n8115 2.2505
R21890 VSS.n8088 VSS.n7891 2.2505
R21891 VSS.n8674 VSS.n8672 2.2505
R21892 VSS.n8740 VSS.n8663 2.2505
R21893 VSS.n8670 VSS.n8669 2.2505
R21894 VSS.n8645 VSS.n8643 2.2505
R21895 VSS.n8651 VSS.n8649 2.2505
R21896 VSS.n8706 VSS.n8705 2.2505
R21897 VSS.n8939 VSS.n8886 2.2505
R21898 VSS.n8871 VSS.n8856 2.2505
R21899 VSS.n8909 VSS.n8908 2.2505
R21900 VSS.n8979 VSS.n8978 2.2505
R21901 VSS.n8810 VSS.n8808 2.2505
R21902 VSS.n8840 VSS.n8816 2.2505
R21903 VSS.n8989 VSS.n8778 2.2505
R21904 VSS.n8620 VSS.n8619 2.2505
R21905 VSS.n8606 VSS.n221 2.2505
R21906 VSS.n208 VSS.n206 2.2505
R21907 VSS.n8558 VSS.n8557 2.2505
R21908 VSS.n251 VSS.n250 2.2505
R21909 VSS.n8551 VSS.n268 2.2505
R21910 VSS.n1356 VSS.n1354 2.2505
R21911 VSS.n1422 VSS.n1345 2.2505
R21912 VSS.n1352 VSS.n1351 2.2505
R21913 VSS.n1327 VSS.n1325 2.2505
R21914 VSS.n1333 VSS.n1331 2.2505
R21915 VSS.n1388 VSS.n1387 2.2505
R21916 VSS.n1564 VSS.n1563 2.2505
R21917 VSS.n1535 VSS.n1533 2.2505
R21918 VSS.n1605 VSS.n1604 2.2505
R21919 VSS.n1490 VSS.n1488 2.2505
R21920 VSS.n1520 VSS.n1519 2.2505
R21921 VSS.n1522 VSS.n1512 2.2505
R21922 VSS.n1652 VSS.n1651 2.2505
R21923 VSS.n1302 VSS.n1301 2.2505
R21924 VSS.n1288 VSS.n1167 2.2505
R21925 VSS.n1154 VSS.n1152 2.2505
R21926 VSS.n1240 VSS.n1239 2.2505
R21927 VSS.n1197 VSS.n1196 2.2505
R21928 VSS.n1233 VSS.n1214 2.2505
R21929 VSS.n1929 VSS.n1927 2.2505
R21930 VSS.n1995 VSS.n1918 2.2505
R21931 VSS.n1925 VSS.n1924 2.2505
R21932 VSS.n1900 VSS.n1898 2.2505
R21933 VSS.n1906 VSS.n1904 2.2505
R21934 VSS.n1961 VSS.n1960 2.2505
R21935 VSS.n2162 VSS.n2125 2.2505
R21936 VSS.n2108 VSS.n2106 2.2505
R21937 VSS.n2197 VSS.n2196 2.2505
R21938 VSS.n2063 VSS.n2061 2.2505
R21939 VSS.n2093 VSS.n2092 2.2505
R21940 VSS.n2095 VSS.n2085 2.2505
R21941 VSS.n2244 VSS.n2243 2.2505
R21942 VSS.n1875 VSS.n1874 2.2505
R21943 VSS.n1861 VSS.n1740 2.2505
R21944 VSS.n1727 VSS.n1725 2.2505
R21945 VSS.n1813 VSS.n1812 2.2505
R21946 VSS.n1770 VSS.n1769 2.2505
R21947 VSS.n1806 VSS.n1787 2.2505
R21948 VSS.n3776 VSS.n3775 2.2505
R21949 VSS.n3462 VSS.n3460 2.2505
R21950 VSS.n3769 VSS.n3449 2.2505
R21951 VSS.n3705 VSS.n3704 2.2505
R21952 VSS.n3726 VSS.n3725 2.2505
R21953 VSS.n3698 VSS.n3501 2.2505
R21954 VSS.n3938 VSS.n3937 2.2505
R21955 VSS.n3884 VSS.n3874 2.2505
R21956 VSS.n3913 VSS.n3912 2.2505
R21957 VSS.n3838 VSS.n3422 2.2505
R21958 VSS.n3861 VSS.n3860 2.2505
R21959 VSS.n3863 VSS.n3405 2.2505
R21960 VSS.n3428 VSS.n3426 2.2505
R21961 VSS.n3669 VSS.n3668 2.2505
R21962 VSS.n3655 VSS.n3534 2.2505
R21963 VSS.n3521 VSS.n3519 2.2505
R21964 VSS.n3607 VSS.n3606 2.2505
R21965 VSS.n3564 VSS.n3563 2.2505
R21966 VSS.n3600 VSS.n3581 2.2505
R21967 VSS.n4368 VSS.n4367 2.2505
R21968 VSS.n4054 VSS.n4052 2.2505
R21969 VSS.n4361 VSS.n4041 2.2505
R21970 VSS.n4297 VSS.n4296 2.2505
R21971 VSS.n4318 VSS.n4317 2.2505
R21972 VSS.n4290 VSS.n4093 2.2505
R21973 VSS.n4530 VSS.n4529 2.2505
R21974 VSS.n4476 VSS.n4466 2.2505
R21975 VSS.n4505 VSS.n4504 2.2505
R21976 VSS.n4430 VSS.n4014 2.2505
R21977 VSS.n4453 VSS.n4452 2.2505
R21978 VSS.n4455 VSS.n3997 2.2505
R21979 VSS.n4020 VSS.n4018 2.2505
R21980 VSS.n4261 VSS.n4260 2.2505
R21981 VSS.n4247 VSS.n4126 2.2505
R21982 VSS.n4113 VSS.n4111 2.2505
R21983 VSS.n4199 VSS.n4198 2.2505
R21984 VSS.n4156 VSS.n4155 2.2505
R21985 VSS.n4192 VSS.n4173 2.2505
R21986 VSS.n4960 VSS.n4959 2.2505
R21987 VSS.n4646 VSS.n4644 2.2505
R21988 VSS.n4953 VSS.n4633 2.2505
R21989 VSS.n4889 VSS.n4888 2.2505
R21990 VSS.n4910 VSS.n4909 2.2505
R21991 VSS.n4882 VSS.n4685 2.2505
R21992 VSS.n5122 VSS.n5121 2.2505
R21993 VSS.n5068 VSS.n5058 2.2505
R21994 VSS.n5097 VSS.n5096 2.2505
R21995 VSS.n5022 VSS.n4606 2.2505
R21996 VSS.n5045 VSS.n5044 2.2505
R21997 VSS.n5047 VSS.n4589 2.2505
R21998 VSS.n4612 VSS.n4610 2.2505
R21999 VSS.n4853 VSS.n4852 2.2505
R22000 VSS.n4839 VSS.n4718 2.2505
R22001 VSS.n4705 VSS.n4703 2.2505
R22002 VSS.n4791 VSS.n4790 2.2505
R22003 VSS.n4748 VSS.n4747 2.2505
R22004 VSS.n4784 VSS.n4765 2.2505
R22005 VSS.n5552 VSS.n5551 2.2505
R22006 VSS.n5238 VSS.n5236 2.2505
R22007 VSS.n5545 VSS.n5225 2.2505
R22008 VSS.n5481 VSS.n5480 2.2505
R22009 VSS.n5502 VSS.n5501 2.2505
R22010 VSS.n5474 VSS.n5277 2.2505
R22011 VSS.n5714 VSS.n5713 2.2505
R22012 VSS.n5660 VSS.n5650 2.2505
R22013 VSS.n5689 VSS.n5688 2.2505
R22014 VSS.n5614 VSS.n5198 2.2505
R22015 VSS.n5637 VSS.n5636 2.2505
R22016 VSS.n5639 VSS.n5181 2.2505
R22017 VSS.n5204 VSS.n5202 2.2505
R22018 VSS.n5445 VSS.n5444 2.2505
R22019 VSS.n5431 VSS.n5310 2.2505
R22020 VSS.n5297 VSS.n5295 2.2505
R22021 VSS.n5383 VSS.n5382 2.2505
R22022 VSS.n5340 VSS.n5339 2.2505
R22023 VSS.n5376 VSS.n5357 2.2505
R22024 VSS.n6144 VSS.n6143 2.2505
R22025 VSS.n5830 VSS.n5828 2.2505
R22026 VSS.n6137 VSS.n5817 2.2505
R22027 VSS.n6073 VSS.n6072 2.2505
R22028 VSS.n6094 VSS.n6093 2.2505
R22029 VSS.n6066 VSS.n5869 2.2505
R22030 VSS.n6306 VSS.n6305 2.2505
R22031 VSS.n6252 VSS.n6242 2.2505
R22032 VSS.n6281 VSS.n6280 2.2505
R22033 VSS.n6206 VSS.n5790 2.2505
R22034 VSS.n6229 VSS.n6228 2.2505
R22035 VSS.n6231 VSS.n5773 2.2505
R22036 VSS.n5796 VSS.n5794 2.2505
R22037 VSS.n6037 VSS.n6036 2.2505
R22038 VSS.n6023 VSS.n5902 2.2505
R22039 VSS.n5889 VSS.n5887 2.2505
R22040 VSS.n5975 VSS.n5974 2.2505
R22041 VSS.n5932 VSS.n5931 2.2505
R22042 VSS.n5968 VSS.n5949 2.2505
R22043 VSS.n6736 VSS.n6735 2.2505
R22044 VSS.n6422 VSS.n6420 2.2505
R22045 VSS.n6729 VSS.n6409 2.2505
R22046 VSS.n6665 VSS.n6664 2.2505
R22047 VSS.n6686 VSS.n6685 2.2505
R22048 VSS.n6658 VSS.n6461 2.2505
R22049 VSS.n6898 VSS.n6897 2.2505
R22050 VSS.n6844 VSS.n6834 2.2505
R22051 VSS.n6873 VSS.n6872 2.2505
R22052 VSS.n6798 VSS.n6382 2.2505
R22053 VSS.n6821 VSS.n6820 2.2505
R22054 VSS.n6823 VSS.n6365 2.2505
R22055 VSS.n6388 VSS.n6386 2.2505
R22056 VSS.n6629 VSS.n6628 2.2505
R22057 VSS.n6615 VSS.n6494 2.2505
R22058 VSS.n6481 VSS.n6479 2.2505
R22059 VSS.n6567 VSS.n6566 2.2505
R22060 VSS.n6524 VSS.n6523 2.2505
R22061 VSS.n6560 VSS.n6541 2.2505
R22062 VSS.n2527 VSS.n2525 2.2505
R22063 VSS.n2593 VSS.n2516 2.2505
R22064 VSS.n2523 VSS.n2522 2.2505
R22065 VSS.n2498 VSS.n2496 2.2505
R22066 VSS.n2504 VSS.n2502 2.2505
R22067 VSS.n2559 VSS.n2558 2.2505
R22068 VSS.n2760 VSS.n2723 2.2505
R22069 VSS.n2706 VSS.n2704 2.2505
R22070 VSS.n6941 VSS.n6940 2.2505
R22071 VSS.n2661 VSS.n2659 2.2505
R22072 VSS.n2691 VSS.n2690 2.2505
R22073 VSS.n2693 VSS.n2683 2.2505
R22074 VSS.n6988 VSS.n6987 2.2505
R22075 VSS.n2473 VSS.n2472 2.2505
R22076 VSS.n2459 VSS.n2338 2.2505
R22077 VSS.n2325 VSS.n2323 2.2505
R22078 VSS.n2411 VSS.n2410 2.2505
R22079 VSS.n2368 VSS.n2367 2.2505
R22080 VSS.n2404 VSS.n2385 2.2505
R22081 VSS.n3184 VSS.n3183 2.2505
R22082 VSS.n2869 VSS.n2867 2.2505
R22083 VSS.n3177 VSS.n2856 2.2505
R22084 VSS.n3113 VSS.n3112 2.2505
R22085 VSS.n3134 VSS.n3133 2.2505
R22086 VSS.n3106 VSS.n2908 2.2505
R22087 VSS.n3346 VSS.n3345 2.2505
R22088 VSS.n3292 VSS.n3282 2.2505
R22089 VSS.n3321 VSS.n3320 2.2505
R22090 VSS.n3246 VSS.n2829 2.2505
R22091 VSS.n3269 VSS.n3268 2.2505
R22092 VSS.n3271 VSS.n2812 2.2505
R22093 VSS.n2835 VSS.n2833 2.2505
R22094 VSS.n3080 VSS.n3079 2.2505
R22095 VSS.n2944 VSS.n2942 2.2505
R22096 VSS.n3073 VSS.n2931 2.2505
R22097 VSS.n3008 VSS.n3007 2.2505
R22098 VSS.n3029 VSS.n3028 2.2505
R22099 VSS.n3001 VSS.n2983 2.2505
R22100 VSS.n9144 VSS.n9143 2.2505
R22101 VSS.n136 VSS.n134 2.2505
R22102 VSS.n9137 VSS.n123 2.2505
R22103 VSS.n9073 VSS.n9072 2.2505
R22104 VSS.n9094 VSS.n9093 2.2505
R22105 VSS.n9066 VSS.n175 2.2505
R22106 VSS.n9306 VSS.n9305 2.2505
R22107 VSS.n9252 VSS.n9242 2.2505
R22108 VSS.n9281 VSS.n9280 2.2505
R22109 VSS.n9206 VSS.n96 2.2505
R22110 VSS.n9229 VSS.n9228 2.2505
R22111 VSS.n9231 VSS.n79 2.2505
R22112 VSS.n102 VSS.n100 2.2505
R22113 VSS.n397 VSS.n396 2.2505
R22114 VSS.n317 VSS.n300 2.2505
R22115 VSS.n307 VSS.n306 2.2505
R22116 VSS.n281 VSS.n279 2.2505
R22117 VSS.n287 VSS.n285 2.2505
R22118 VSS.n332 VSS.n331 2.2505
R22119 VSS.n516 VSS.n514 2.2505
R22120 VSS.n585 VSS.n505 2.2505
R22121 VSS.n512 VSS.n511 2.2505
R22122 VSS.n487 VSS.n485 2.2505
R22123 VSS.n493 VSS.n491 2.2505
R22124 VSS.n483 VSS.n482 2.2505
R22125 VSS.n807 VSS.n806 2.2505
R22126 VSS.n653 VSS.n651 2.2505
R22127 VSS.n683 VSS.n682 2.2505
R22128 VSS.n698 VSS.n696 2.2505
R22129 VSS.n760 VSS.n759 2.2505
R22130 VSS.n726 VSS.n725 2.2505
R22131 VSS.n685 VSS.n675 2.2505
R22132 VSS.n477 VSS.n475 2.2505
R22133 VSS.n928 VSS.n466 2.2505
R22134 VSS.n473 VSS.n472 2.2505
R22135 VSS.n447 VSS.n445 2.2505
R22136 VSS.n453 VSS.n451 2.2505
R22137 VSS.n896 VSS.n895 2.2505
R22138 VSS.n7328 VSS.n7291 2.2505
R22139 VSS.n7274 VSS.n7272 2.2505
R22140 VSS.n8369 VSS.n8368 2.2505
R22141 VSS.n7229 VSS.n7227 2.2505
R22142 VSS.n7259 VSS.n7258 2.2505
R22143 VSS.n7261 VSS.n7251 2.2505
R22144 VSS.n8416 VSS.n8415 2.2505
R22145 VSS.n9323 VSS.n37 2.24315
R22146 VSS.n6915 VSS.n6323 2.24315
R22147 VSS.n4547 VSS.n3955 2.24315
R22148 VSS.n8344 VSS.n7752 2.24315
R22149 VSS.n7692 VSS.n7691 2.10336
R22150 VSS.n8284 VSS.n8283 2.10336
R22151 VSS.n8961 VSS.n8821 2.10336
R22152 VSS.n1622 VSS.n1621 2.10336
R22153 VSS.n2214 VSS.n2213 2.10336
R22154 VSS.n3894 VSS.n3893 2.10336
R22155 VSS.n4486 VSS.n4485 2.10336
R22156 VSS.n5078 VSS.n5077 2.10336
R22157 VSS.n5670 VSS.n5669 2.10336
R22158 VSS.n6262 VSS.n6261 2.10336
R22159 VSS.n6854 VSS.n6853 2.10336
R22160 VSS.n6958 VSS.n6957 2.10336
R22161 VSS.n3302 VSS.n3301 2.10336
R22162 VSS.n9262 VSS.n9261 2.10336
R22163 VSS.n777 VSS.n776 2.10336
R22164 VSS.n8386 VSS.n8385 2.10336
R22165 VSS.n7692 VSS.n7374 2.01193
R22166 VSS.n8284 VSS.n7788 2.01193
R22167 VSS.n8962 VSS.n8961 2.01193
R22168 VSS.n1622 VSS.n1505 2.01193
R22169 VSS.n2214 VSS.n2078 2.01193
R22170 VSS.n3894 VSS.n3398 2.01193
R22171 VSS.n4486 VSS.n3990 2.01193
R22172 VSS.n5078 VSS.n4582 2.01193
R22173 VSS.n5670 VSS.n5174 2.01193
R22174 VSS.n6262 VSS.n5766 2.01193
R22175 VSS.n6854 VSS.n6358 2.01193
R22176 VSS.n6958 VSS.n2676 2.01193
R22177 VSS.n3302 VSS.n2805 2.01193
R22178 VSS.n9262 VSS.n72 2.01193
R22179 VSS.n777 VSS.n668 2.01193
R22180 VSS.n8386 VSS.n7244 2.01193
R22181 VSS.n8472 VSS.n8471 1.98071
R22182 VSS.n1000 VSS.n999 1.98071
R22183 VSS.n7489 VSS.n7485 1.98071
R22184 VSS.n8521 VSS.n8520 1.98071
R22185 VSS.n8081 VSS.n7899 1.98071
R22186 VSS.n7983 VSS.n7980 1.98071
R22187 VSS.n8544 VSS.n8541 1.98071
R22188 VSS.n9045 VSS.n9044 1.98071
R22189 VSS.n1226 VSS.n1223 1.98071
R22190 VSS.n1708 VSS.n1707 1.98071
R22191 VSS.n1799 VSS.n1796 1.98071
R22192 VSS.n2300 VSS.n2299 1.98071
R22193 VSS.n3593 VSS.n3590 1.98071
R22194 VSS.n3691 VSS.n3509 1.98071
R22195 VSS.n4185 VSS.n4182 1.98071
R22196 VSS.n4283 VSS.n4101 1.98071
R22197 VSS.n4777 VSS.n4774 1.98071
R22198 VSS.n4875 VSS.n4693 1.98071
R22199 VSS.n5369 VSS.n5366 1.98071
R22200 VSS.n5467 VSS.n5285 1.98071
R22201 VSS.n5961 VSS.n5958 1.98071
R22202 VSS.n6059 VSS.n5877 1.98071
R22203 VSS.n6553 VSS.n6550 1.98071
R22204 VSS.n6651 VSS.n6469 1.98071
R22205 VSS.n2397 VSS.n2394 1.98071
R22206 VSS.n7044 VSS.n7043 1.98071
R22207 VSS.n2994 VSS.n2991 1.98071
R22208 VSS.n3099 VSS.n2916 1.98071
R22209 VSS.n435 VSS.n434 1.98071
R22210 VSS.n9059 VSS.n176 1.98071
R22211 VSS.n861 VSS.n481 1.98071
R22212 VSS.n7657 VSS.n7384 1.94045
R22213 VSS.n8249 VSS.n7798 1.94045
R22214 VSS.n8969 VSS.n8968 1.94045
R22215 VSS.n1518 VSS.n1514 1.94045
R22216 VSS.n2091 VSS.n2087 1.94045
R22217 VSS.n3859 VSS.n3408 1.94045
R22218 VSS.n4451 VSS.n4000 1.94045
R22219 VSS.n5043 VSS.n4592 1.94045
R22220 VSS.n5635 VSS.n5184 1.94045
R22221 VSS.n6227 VSS.n5776 1.94045
R22222 VSS.n6819 VSS.n6368 1.94045
R22223 VSS.n2689 VSS.n2685 1.94045
R22224 VSS.n3267 VSS.n2815 1.94045
R22225 VSS.n9227 VSS.n82 1.94045
R22226 VSS.n681 VSS.n677 1.94045
R22227 VSS.n7257 VSS.n7253 1.94045
R22228 VSS VSS.n5139 1.86079
R22229 VSS VSS.n9323 1.85712
R22230 VSS VSS.n6915 1.85712
R22231 VSS VSS.n4547 1.85712
R22232 VSS.n7752 VSS 1.85712
R22233 VSS.n6916 VSS 1.563
R22234 VSS VSS.n9352 1.563
R22235 VSS.n7135 VSS.n7123 1.55479
R22236 VSS.n1085 VSS.n1073 1.55479
R22237 VSS.n7505 VSS.n7469 1.55479
R22238 VSS.n7999 VSS.n7962 1.55479
R22239 VSS.n8097 VSS.n7883 1.55479
R22240 VSS.n8714 VSS.n8702 1.55479
R22241 VSS.n8560 VSS.n259 1.55479
R22242 VSS.n1396 VSS.n1384 1.55479
R22243 VSS.n1242 VSS.n1205 1.55479
R22244 VSS.n1969 VSS.n1957 1.55479
R22245 VSS.n1815 VSS.n1778 1.55479
R22246 VSS.n3707 VSS.n3493 1.55479
R22247 VSS.n3609 VSS.n3572 1.55479
R22248 VSS.n4299 VSS.n4085 1.55479
R22249 VSS.n4201 VSS.n4164 1.55479
R22250 VSS.n4891 VSS.n4677 1.55479
R22251 VSS.n4793 VSS.n4756 1.55479
R22252 VSS.n5483 VSS.n5269 1.55479
R22253 VSS.n5385 VSS.n5348 1.55479
R22254 VSS.n6075 VSS.n5861 1.55479
R22255 VSS.n5977 VSS.n5940 1.55479
R22256 VSS.n6667 VSS.n6453 1.55479
R22257 VSS.n6569 VSS.n6532 1.55479
R22258 VSS.n2567 VSS.n2555 1.55479
R22259 VSS.n2413 VSS.n2376 1.55479
R22260 VSS.n3115 VSS.n2900 1.55479
R22261 VSS.n3010 VSS.n2975 1.55479
R22262 VSS.n9075 VSS.n167 1.55479
R22263 VSS.n340 VSS.n327 1.55479
R22264 VSS.n559 VSS.n549 1.55479
R22265 VSS.n904 VSS.n892 1.55479
R22266 VSS.n7647 VSS.n7393 1.53956
R22267 VSS.n7697 VSS.n7361 1.53956
R22268 VSS.n8239 VSS.n7807 1.53956
R22269 VSS.n8289 VSS.n7775 1.53956
R22270 VSS.n8844 VSS.n8836 1.53956
R22271 VSS.n8956 VSS.n8848 1.53956
R22272 VSS.n1627 VSS.n1486 1.53956
R22273 VSS.n1583 VSS.n1580 1.53956
R22274 VSS.n2219 VSS.n2059 1.53956
R22275 VSS.n2143 VSS.n2140 1.53956
R22276 VSS.n3849 VSS.n3417 1.53956
R22277 VSS.n3899 VSS.n3385 1.53956
R22278 VSS.n4441 VSS.n4009 1.53956
R22279 VSS.n4491 VSS.n3977 1.53956
R22280 VSS.n5033 VSS.n4601 1.53956
R22281 VSS.n5083 VSS.n4569 1.53956
R22282 VSS.n5625 VSS.n5193 1.53956
R22283 VSS.n5675 VSS.n5161 1.53956
R22284 VSS.n6217 VSS.n5785 1.53956
R22285 VSS.n6267 VSS.n5753 1.53956
R22286 VSS.n6809 VSS.n6377 1.53956
R22287 VSS.n6859 VSS.n6345 1.53956
R22288 VSS.n6963 VSS.n2657 1.53956
R22289 VSS.n2741 VSS.n2738 1.53956
R22290 VSS.n3257 VSS.n2824 1.53956
R22291 VSS.n3307 VSS.n2792 1.53956
R22292 VSS.n9217 VSS.n91 1.53956
R22293 VSS.n9267 VSS.n59 1.53956
R22294 VSS.n782 VSS.n649 1.53956
R22295 VSS.n741 VSS.n740 1.53956
R22296 VSS.n8391 VSS.n7225 1.53956
R22297 VSS.n7309 VSS.n7306 1.53956
R22298 VSS.n1029 VSS.n1027 1.5005
R22299 VSS.n8032 VSS.n8031 1.5005
R22300 VSS.n8593 VSS.n8592 1.5005
R22301 VSS.n1275 VSS.n1274 1.5005
R22302 VSS.n1848 VSS.n1847 1.5005
R22303 VSS.n3642 VSS.n3641 1.5005
R22304 VSS.n4234 VSS.n4233 1.5005
R22305 VSS.n4826 VSS.n4825 1.5005
R22306 VSS.n5418 VSS.n5417 1.5005
R22307 VSS.n6010 VSS.n6009 1.5005
R22308 VSS.n6602 VSS.n6601 1.5005
R22309 VSS.n2446 VSS.n2445 1.5005
R22310 VSS.n2956 VSS.n2955 1.5005
R22311 VSS.n296 VSS.n294 1.5005
R22312 VSS.n462 VSS.n460 1.5005
R22313 VSS.n7176 VSS.n7102 1.46336
R22314 VSS.n1125 VSS.n1051 1.46336
R22315 VSS.n7391 VSS.n7383 1.46336
R22316 VSS.n7698 VSS.n7370 1.46336
R22317 VSS.n7564 VSS.n7419 1.46336
R22318 VSS.n7914 VSS.n7908 1.46336
R22319 VSS.n7805 VSS.n7797 1.46336
R22320 VSS.n8290 VSS.n7784 1.46336
R22321 VSS.n8156 VSS.n7833 1.46336
R22322 VSS.n8755 VSS.n8681 1.46336
R22323 VSS.n8843 VSS.n8842 1.46336
R22324 VSS.n8955 VSS.n8849 1.46336
R22325 VSS.n211 VSS.n205 1.46336
R22326 VSS.n1437 VSS.n1363 1.46336
R22327 VSS.n1628 VSS.n1501 1.46336
R22328 VSS.n1579 VSS.n1578 1.46336
R22329 VSS.n1157 VSS.n1151 1.46336
R22330 VSS.n2010 VSS.n1936 1.46336
R22331 VSS.n2220 VSS.n2074 1.46336
R22332 VSS.n2139 VSS.n2138 1.46336
R22333 VSS.n1730 VSS.n1724 1.46336
R22334 VSS.n3766 VSS.n3443 1.46336
R22335 VSS.n3415 VSS.n3407 1.46336
R22336 VSS.n3900 VSS.n3394 1.46336
R22337 VSS.n3524 VSS.n3518 1.46336
R22338 VSS.n4358 VSS.n4035 1.46336
R22339 VSS.n4007 VSS.n3999 1.46336
R22340 VSS.n4492 VSS.n3986 1.46336
R22341 VSS.n4116 VSS.n4110 1.46336
R22342 VSS.n4950 VSS.n4627 1.46336
R22343 VSS.n4599 VSS.n4591 1.46336
R22344 VSS.n5084 VSS.n4578 1.46336
R22345 VSS.n4708 VSS.n4702 1.46336
R22346 VSS.n5542 VSS.n5219 1.46336
R22347 VSS.n5191 VSS.n5183 1.46336
R22348 VSS.n5676 VSS.n5170 1.46336
R22349 VSS.n5300 VSS.n5294 1.46336
R22350 VSS.n6134 VSS.n5811 1.46336
R22351 VSS.n5783 VSS.n5775 1.46336
R22352 VSS.n6268 VSS.n5762 1.46336
R22353 VSS.n5892 VSS.n5886 1.46336
R22354 VSS.n6726 VSS.n6403 1.46336
R22355 VSS.n6375 VSS.n6367 1.46336
R22356 VSS.n6860 VSS.n6354 1.46336
R22357 VSS.n6484 VSS.n6478 1.46336
R22358 VSS.n2608 VSS.n2534 1.46336
R22359 VSS.n6964 VSS.n2672 1.46336
R22360 VSS.n2737 VSS.n2736 1.46336
R22361 VSS.n2328 VSS.n2322 1.46336
R22362 VSS.n3174 VSS.n2850 1.46336
R22363 VSS.n2822 VSS.n2814 1.46336
R22364 VSS.n3308 VSS.n2801 1.46336
R22365 VSS.n3070 VSS.n2925 1.46336
R22366 VSS.n9134 VSS.n117 1.46336
R22367 VSS.n89 VSS.n81 1.46336
R22368 VSS.n9268 VSS.n68 1.46336
R22369 VSS.n389 VSS.n312 1.46336
R22370 VSS.n600 VSS.n523 1.46336
R22371 VSS.n783 VSS.n664 1.46336
R22372 VSS.n738 VSS.n737 1.46336
R22373 VSS.n944 VSS.n870 1.46336
R22374 VSS.n8392 VSS.n7240 1.46336
R22375 VSS.n7305 VSS.n7304 1.46336
R22376 VSS.n7142 VSS.n7115 1.37193
R22377 VSS.n7152 VSS.n7151 1.37193
R22378 VSS.n7159 VSS.n7158 1.37193
R22379 VSS.n7162 VSS.n7160 1.37193
R22380 VSS.n1090 VSS.n1065 1.37193
R22381 VSS.n1100 VSS.n1099 1.37193
R22382 VSS.n1107 VSS.n1106 1.37193
R22383 VSS.n1110 VSS.n1108 1.37193
R22384 VSS.n7512 VSS.n7455 1.37193
R22385 VSS.n7527 VSS.n7449 1.37193
R22386 VSS.n7450 VSS.n7434 1.37193
R22387 VSS.n7550 VSS.n7435 1.37193
R22388 VSS.n8011 VSS.n7956 1.37193
R22389 VSS.n7957 VSS.n7939 1.37193
R22390 VSS.n8035 VSS.n7927 1.37193
R22391 VSS.n7934 VSS.n7928 1.37193
R22392 VSS.n8104 VSS.n7869 1.37193
R22393 VSS.n8119 VSS.n7863 1.37193
R22394 VSS.n7864 VSS.n7848 1.37193
R22395 VSS.n8142 VSS.n7849 1.37193
R22396 VSS.n8721 VSS.n8694 1.37193
R22397 VSS.n8731 VSS.n8730 1.37193
R22398 VSS.n8738 VSS.n8737 1.37193
R22399 VSS.n8741 VSS.n8739 1.37193
R22400 VSS.n8572 VSS.n253 1.37193
R22401 VSS.n254 VSS.n236 1.37193
R22402 VSS.n8596 VSS.n224 1.37193
R22403 VSS.n231 VSS.n225 1.37193
R22404 VSS.n1403 VSS.n1376 1.37193
R22405 VSS.n1413 VSS.n1412 1.37193
R22406 VSS.n1420 VSS.n1419 1.37193
R22407 VSS.n1423 VSS.n1421 1.37193
R22408 VSS.n1254 VSS.n1199 1.37193
R22409 VSS.n1200 VSS.n1182 1.37193
R22410 VSS.n1278 VSS.n1170 1.37193
R22411 VSS.n1177 VSS.n1171 1.37193
R22412 VSS.n1976 VSS.n1949 1.37193
R22413 VSS.n1986 VSS.n1985 1.37193
R22414 VSS.n1993 VSS.n1992 1.37193
R22415 VSS.n1996 VSS.n1994 1.37193
R22416 VSS.n1827 VSS.n1772 1.37193
R22417 VSS.n1773 VSS.n1755 1.37193
R22418 VSS.n1851 VSS.n1743 1.37193
R22419 VSS.n1750 VSS.n1744 1.37193
R22420 VSS.n3714 VSS.n3479 1.37193
R22421 VSS.n3729 VSS.n3473 1.37193
R22422 VSS.n3474 VSS.n3458 1.37193
R22423 VSS.n3752 VSS.n3459 1.37193
R22424 VSS.n3621 VSS.n3566 1.37193
R22425 VSS.n3567 VSS.n3549 1.37193
R22426 VSS.n3645 VSS.n3537 1.37193
R22427 VSS.n3544 VSS.n3538 1.37193
R22428 VSS.n4306 VSS.n4071 1.37193
R22429 VSS.n4321 VSS.n4065 1.37193
R22430 VSS.n4066 VSS.n4050 1.37193
R22431 VSS.n4344 VSS.n4051 1.37193
R22432 VSS.n4213 VSS.n4158 1.37193
R22433 VSS.n4159 VSS.n4141 1.37193
R22434 VSS.n4237 VSS.n4129 1.37193
R22435 VSS.n4136 VSS.n4130 1.37193
R22436 VSS.n4898 VSS.n4663 1.37193
R22437 VSS.n4913 VSS.n4657 1.37193
R22438 VSS.n4658 VSS.n4642 1.37193
R22439 VSS.n4936 VSS.n4643 1.37193
R22440 VSS.n4805 VSS.n4750 1.37193
R22441 VSS.n4751 VSS.n4733 1.37193
R22442 VSS.n4829 VSS.n4721 1.37193
R22443 VSS.n4728 VSS.n4722 1.37193
R22444 VSS.n5490 VSS.n5255 1.37193
R22445 VSS.n5505 VSS.n5249 1.37193
R22446 VSS.n5250 VSS.n5234 1.37193
R22447 VSS.n5528 VSS.n5235 1.37193
R22448 VSS.n5397 VSS.n5342 1.37193
R22449 VSS.n5343 VSS.n5325 1.37193
R22450 VSS.n5421 VSS.n5313 1.37193
R22451 VSS.n5320 VSS.n5314 1.37193
R22452 VSS.n6082 VSS.n5847 1.37193
R22453 VSS.n6097 VSS.n5841 1.37193
R22454 VSS.n5842 VSS.n5826 1.37193
R22455 VSS.n6120 VSS.n5827 1.37193
R22456 VSS.n5989 VSS.n5934 1.37193
R22457 VSS.n5935 VSS.n5917 1.37193
R22458 VSS.n6013 VSS.n5905 1.37193
R22459 VSS.n5912 VSS.n5906 1.37193
R22460 VSS.n6674 VSS.n6439 1.37193
R22461 VSS.n6689 VSS.n6433 1.37193
R22462 VSS.n6434 VSS.n6418 1.37193
R22463 VSS.n6712 VSS.n6419 1.37193
R22464 VSS.n6581 VSS.n6526 1.37193
R22465 VSS.n6527 VSS.n6509 1.37193
R22466 VSS.n6605 VSS.n6497 1.37193
R22467 VSS.n6504 VSS.n6498 1.37193
R22468 VSS.n2574 VSS.n2547 1.37193
R22469 VSS.n2584 VSS.n2583 1.37193
R22470 VSS.n2591 VSS.n2590 1.37193
R22471 VSS.n2594 VSS.n2592 1.37193
R22472 VSS.n2425 VSS.n2370 1.37193
R22473 VSS.n2371 VSS.n2353 1.37193
R22474 VSS.n2449 VSS.n2341 1.37193
R22475 VSS.n2348 VSS.n2342 1.37193
R22476 VSS.n3122 VSS.n2886 1.37193
R22477 VSS.n3137 VSS.n2880 1.37193
R22478 VSS.n2881 VSS.n2865 1.37193
R22479 VSS.n3160 VSS.n2866 1.37193
R22480 VSS.n3017 VSS.n2963 1.37193
R22481 VSS.n3032 VSS.n2957 1.37193
R22482 VSS.n2958 VSS.n2940 1.37193
R22483 VSS.n3055 VSS.n2941 1.37193
R22484 VSS.n9082 VSS.n153 1.37193
R22485 VSS.n9097 VSS.n147 1.37193
R22486 VSS.n148 VSS.n132 1.37193
R22487 VSS.n9120 VSS.n133 1.37193
R22488 VSS.n349 VSS.n326 1.37193
R22489 VSS.n361 VSS.n322 1.37193
R22490 VSS.n364 VSS.n318 1.37193
R22491 VSS.n377 VSS.n316 1.37193
R22492 VSS.n566 VSS.n536 1.37193
R22493 VSS.n576 VSS.n575 1.37193
R22494 VSS.n583 VSS.n582 1.37193
R22495 VSS.n586 VSS.n584 1.37193
R22496 VSS.n909 VSS.n884 1.37193
R22497 VSS.n919 VSS.n918 1.37193
R22498 VSS.n926 VSS.n925 1.37193
R22499 VSS.n929 VSS.n927 1.37193
R22500 VSS.n7641 VSS.n7640 1.2805
R22501 VSS.n7713 VSS.n7358 1.2805
R22502 VSS.n8233 VSS.n8232 1.2805
R22503 VSS.n8305 VSS.n7772 1.2805
R22504 VSS.n8829 VSS.n8806 1.2805
R22505 VSS.n8911 VSS.n8905 1.2805
R22506 VSS.n1638 VSS.n1483 1.2805
R22507 VSS.n1587 VSS.n1538 1.2805
R22508 VSS.n2230 VSS.n2056 1.2805
R22509 VSS.n2147 VSS.n2111 1.2805
R22510 VSS.n3843 VSS.n3842 1.2805
R22511 VSS.n3915 VSS.n3382 1.2805
R22512 VSS.n4435 VSS.n4434 1.2805
R22513 VSS.n4507 VSS.n3974 1.2805
R22514 VSS.n5027 VSS.n5026 1.2805
R22515 VSS.n5099 VSS.n4566 1.2805
R22516 VSS.n5619 VSS.n5618 1.2805
R22517 VSS.n5691 VSS.n5158 1.2805
R22518 VSS.n6211 VSS.n6210 1.2805
R22519 VSS.n6283 VSS.n5750 1.2805
R22520 VSS.n6803 VSS.n6802 1.2805
R22521 VSS.n6875 VSS.n6342 1.2805
R22522 VSS.n6974 VSS.n2654 1.2805
R22523 VSS.n2745 VSS.n2709 1.2805
R22524 VSS.n3251 VSS.n3250 1.2805
R22525 VSS.n3323 VSS.n2789 1.2805
R22526 VSS.n9211 VSS.n9210 1.2805
R22527 VSS.n9283 VSS.n56 1.2805
R22528 VSS.n793 VSS.n646 1.2805
R22529 VSS.n727 VSS.n701 1.2805
R22530 VSS.n8402 VSS.n7222 1.2805
R22531 VSS.n7313 VSS.n7277 1.2805
R22532 VSS.n7144 VSS.n7143 1.18907
R22533 VSS.n7174 VSS.n7107 1.18907
R22534 VSS.n1092 VSS.n1091 1.18907
R22535 VSS.n1123 VSS.n1056 1.18907
R22536 VSS.n7511 VSS.n7466 1.18907
R22537 VSS.n7563 VSS.n7430 1.18907
R22538 VSS.n8001 VSS.n8000 1.18907
R22539 VSS.n7935 VSS.n7907 1.18907
R22540 VSS.n8103 VSS.n7880 1.18907
R22541 VSS.n8155 VSS.n7844 1.18907
R22542 VSS.n8723 VSS.n8722 1.18907
R22543 VSS.n8753 VSS.n8686 1.18907
R22544 VSS.n8562 VSS.n8561 1.18907
R22545 VSS.n232 VSS.n204 1.18907
R22546 VSS.n1405 VSS.n1404 1.18907
R22547 VSS.n1435 VSS.n1368 1.18907
R22548 VSS.n1244 VSS.n1243 1.18907
R22549 VSS.n1178 VSS.n1150 1.18907
R22550 VSS.n1978 VSS.n1977 1.18907
R22551 VSS.n2008 VSS.n1941 1.18907
R22552 VSS.n1817 VSS.n1816 1.18907
R22553 VSS.n1751 VSS.n1723 1.18907
R22554 VSS.n3713 VSS.n3490 1.18907
R22555 VSS.n3765 VSS.n3454 1.18907
R22556 VSS.n3611 VSS.n3610 1.18907
R22557 VSS.n3545 VSS.n3517 1.18907
R22558 VSS.n4305 VSS.n4082 1.18907
R22559 VSS.n4357 VSS.n4046 1.18907
R22560 VSS.n4203 VSS.n4202 1.18907
R22561 VSS.n4137 VSS.n4109 1.18907
R22562 VSS.n4897 VSS.n4674 1.18907
R22563 VSS.n4949 VSS.n4638 1.18907
R22564 VSS.n4795 VSS.n4794 1.18907
R22565 VSS.n4729 VSS.n4701 1.18907
R22566 VSS.n5489 VSS.n5266 1.18907
R22567 VSS.n5541 VSS.n5230 1.18907
R22568 VSS.n5387 VSS.n5386 1.18907
R22569 VSS.n5321 VSS.n5293 1.18907
R22570 VSS.n6081 VSS.n5858 1.18907
R22571 VSS.n6133 VSS.n5822 1.18907
R22572 VSS.n5979 VSS.n5978 1.18907
R22573 VSS.n5913 VSS.n5885 1.18907
R22574 VSS.n6673 VSS.n6450 1.18907
R22575 VSS.n6725 VSS.n6414 1.18907
R22576 VSS.n6571 VSS.n6570 1.18907
R22577 VSS.n6505 VSS.n6477 1.18907
R22578 VSS.n2576 VSS.n2575 1.18907
R22579 VSS.n2606 VSS.n2539 1.18907
R22580 VSS.n2415 VSS.n2414 1.18907
R22581 VSS.n2349 VSS.n2321 1.18907
R22582 VSS.n3121 VSS.n2897 1.18907
R22583 VSS.n3173 VSS.n2861 1.18907
R22584 VSS.n3016 VSS.n2972 1.18907
R22585 VSS.n3069 VSS.n2936 1.18907
R22586 VSS.n9081 VSS.n164 1.18907
R22587 VSS.n9133 VSS.n128 1.18907
R22588 VSS.n348 VSS.n347 1.18907
R22589 VSS.n381 VSS.n378 1.18907
R22590 VSS.n568 VSS.n567 1.18907
R22591 VSS.n598 VSS.n528 1.18907
R22592 VSS.n911 VSS.n910 1.18907
R22593 VSS.n942 VSS.n875 1.18907
R22594 VSS.n8518 VSS.n8517 1.13717
R22595 VSS.n1013 VSS.n1011 1.13717
R22596 VSS.n1022 VSS.n1017 1.13717
R22597 VSS.n1034 VSS.n1032 1.13717
R22598 VSS.n1037 VSS.n1035 1.13717
R22599 VSS.n1043 VSS.n1041 1.13717
R22600 VSS.n7615 VSS.n7614 1.13717
R22601 VSS.n7656 VSS.n7655 1.13717
R22602 VSS.n7673 VSS.n7671 1.13717
R22603 VSS.n7340 VSS.n7339 1.13717
R22604 VSS.n7476 VSS.n7475 1.13717
R22605 VSS.n7474 VSS.n7461 1.13717
R22606 VSS.n7520 VSS.n7519 1.13717
R22607 VSS.n7444 VSS.n7440 1.13717
R22608 VSS.n7424 VSS.n7423 1.13717
R22609 VSS.n7412 VSS.n7411 1.13717
R22610 VSS.n7970 VSS.n7969 1.13717
R22611 VSS.n7968 VSS.n7949 1.13717
R22612 VSS.n8019 VSS.n8018 1.13717
R22613 VSS.n8026 VSS.n7922 1.13717
R22614 VSS.n7919 VSS.n7918 1.13717
R22615 VSS.n7901 VSS.n7900 1.13717
R22616 VSS.n8207 VSS.n8206 1.13717
R22617 VSS.n8248 VSS.n8247 1.13717
R22618 VSS.n8265 VSS.n8263 1.13717
R22619 VSS.n7754 VSS.n7753 1.13717
R22620 VSS.n7890 VSS.n7889 1.13717
R22621 VSS.n7888 VSS.n7875 1.13717
R22622 VSS.n8112 VSS.n8111 1.13717
R22623 VSS.n7858 VSS.n7854 1.13717
R22624 VSS.n7838 VSS.n7837 1.13717
R22625 VSS.n7826 VSS.n7825 1.13717
R22626 VSS.n9042 VSS.n9041 1.13717
R22627 VSS.n8644 VSS.n8642 1.13717
R22628 VSS.n8653 VSS.n8648 1.13717
R22629 VSS.n8664 VSS.n8662 1.13717
R22630 VSS.n8667 VSS.n8665 1.13717
R22631 VSS.n8673 VSS.n8671 1.13717
R22632 VSS.n8793 VSS.n8792 1.13717
R22633 VSS.n8814 VSS.n8809 1.13717
R22634 VSS.n8876 VSS.n8875 1.13717
R22635 VSS.n8931 VSS.n8930 1.13717
R22636 VSS.n267 VSS.n266 1.13717
R22637 VSS.n265 VSS.n246 1.13717
R22638 VSS.n8580 VSS.n8579 1.13717
R22639 VSS.n8587 VSS.n219 1.13717
R22640 VSS.n216 VSS.n215 1.13717
R22641 VSS.n198 VSS.n197 1.13717
R22642 VSS.n1705 VSS.n1704 1.13717
R22643 VSS.n1326 VSS.n1324 1.13717
R22644 VSS.n1335 VSS.n1330 1.13717
R22645 VSS.n1346 VSS.n1344 1.13717
R22646 VSS.n1349 VSS.n1347 1.13717
R22647 VSS.n1355 VSS.n1353 1.13717
R22648 VSS.n1474 VSS.n1473 1.13717
R22649 VSS.n1517 VSS.n1516 1.13717
R22650 VSS.n1545 VSS.n1532 1.13717
R22651 VSS.n2 VSS.n1 1.13717
R22652 VSS.n1213 VSS.n1212 1.13717
R22653 VSS.n1211 VSS.n1192 1.13717
R22654 VSS.n1262 VSS.n1261 1.13717
R22655 VSS.n1269 VSS.n1165 1.13717
R22656 VSS.n1162 VSS.n1161 1.13717
R22657 VSS.n1144 VSS.n1143 1.13717
R22658 VSS.n2297 VSS.n2296 1.13717
R22659 VSS.n1899 VSS.n1897 1.13717
R22660 VSS.n1908 VSS.n1903 1.13717
R22661 VSS.n1919 VSS.n1917 1.13717
R22662 VSS.n1922 VSS.n1920 1.13717
R22663 VSS.n1928 VSS.n1926 1.13717
R22664 VSS.n2047 VSS.n2046 1.13717
R22665 VSS.n2090 VSS.n2089 1.13717
R22666 VSS.n2118 VSS.n2105 1.13717
R22667 VSS.n2172 VSS.n2155 1.13717
R22668 VSS.n1786 VSS.n1785 1.13717
R22669 VSS.n1784 VSS.n1765 1.13717
R22670 VSS.n1835 VSS.n1834 1.13717
R22671 VSS.n1842 VSS.n1738 1.13717
R22672 VSS.n1735 VSS.n1734 1.13717
R22673 VSS.n1717 VSS.n1716 1.13717
R22674 VSS.n3500 VSS.n3499 1.13717
R22675 VSS.n3498 VSS.n3485 1.13717
R22676 VSS.n3722 VSS.n3721 1.13717
R22677 VSS.n3468 VSS.n3464 1.13717
R22678 VSS.n3448 VSS.n3447 1.13717
R22679 VSS.n3436 VSS.n3435 1.13717
R22680 VSS.n3817 VSS.n3816 1.13717
R22681 VSS.n3858 VSS.n3857 1.13717
R22682 VSS.n3875 VSS.n3873 1.13717
R22683 VSS.n3365 VSS.n3364 1.13717
R22684 VSS.n3580 VSS.n3579 1.13717
R22685 VSS.n3578 VSS.n3559 1.13717
R22686 VSS.n3629 VSS.n3628 1.13717
R22687 VSS.n3636 VSS.n3532 1.13717
R22688 VSS.n3529 VSS.n3528 1.13717
R22689 VSS.n3511 VSS.n3510 1.13717
R22690 VSS.n4092 VSS.n4091 1.13717
R22691 VSS.n4090 VSS.n4077 1.13717
R22692 VSS.n4314 VSS.n4313 1.13717
R22693 VSS.n4060 VSS.n4056 1.13717
R22694 VSS.n4040 VSS.n4039 1.13717
R22695 VSS.n4028 VSS.n4027 1.13717
R22696 VSS.n4409 VSS.n4408 1.13717
R22697 VSS.n4450 VSS.n4449 1.13717
R22698 VSS.n4467 VSS.n4465 1.13717
R22699 VSS.n3957 VSS.n3956 1.13717
R22700 VSS.n4172 VSS.n4171 1.13717
R22701 VSS.n4170 VSS.n4151 1.13717
R22702 VSS.n4221 VSS.n4220 1.13717
R22703 VSS.n4228 VSS.n4124 1.13717
R22704 VSS.n4121 VSS.n4120 1.13717
R22705 VSS.n4103 VSS.n4102 1.13717
R22706 VSS.n4684 VSS.n4683 1.13717
R22707 VSS.n4682 VSS.n4669 1.13717
R22708 VSS.n4906 VSS.n4905 1.13717
R22709 VSS.n4652 VSS.n4648 1.13717
R22710 VSS.n4632 VSS.n4631 1.13717
R22711 VSS.n4620 VSS.n4619 1.13717
R22712 VSS.n5001 VSS.n5000 1.13717
R22713 VSS.n5042 VSS.n5041 1.13717
R22714 VSS.n5059 VSS.n5057 1.13717
R22715 VSS.n4549 VSS.n4548 1.13717
R22716 VSS.n4764 VSS.n4763 1.13717
R22717 VSS.n4762 VSS.n4743 1.13717
R22718 VSS.n4813 VSS.n4812 1.13717
R22719 VSS.n4820 VSS.n4716 1.13717
R22720 VSS.n4713 VSS.n4712 1.13717
R22721 VSS.n4695 VSS.n4694 1.13717
R22722 VSS.n5276 VSS.n5275 1.13717
R22723 VSS.n5274 VSS.n5261 1.13717
R22724 VSS.n5498 VSS.n5497 1.13717
R22725 VSS.n5244 VSS.n5240 1.13717
R22726 VSS.n5224 VSS.n5223 1.13717
R22727 VSS.n5212 VSS.n5211 1.13717
R22728 VSS.n5593 VSS.n5592 1.13717
R22729 VSS.n5634 VSS.n5633 1.13717
R22730 VSS.n5651 VSS.n5649 1.13717
R22731 VSS.n5141 VSS.n5140 1.13717
R22732 VSS.n5356 VSS.n5355 1.13717
R22733 VSS.n5354 VSS.n5335 1.13717
R22734 VSS.n5405 VSS.n5404 1.13717
R22735 VSS.n5412 VSS.n5308 1.13717
R22736 VSS.n5305 VSS.n5304 1.13717
R22737 VSS.n5287 VSS.n5286 1.13717
R22738 VSS.n5868 VSS.n5867 1.13717
R22739 VSS.n5866 VSS.n5853 1.13717
R22740 VSS.n6090 VSS.n6089 1.13717
R22741 VSS.n5836 VSS.n5832 1.13717
R22742 VSS.n5816 VSS.n5815 1.13717
R22743 VSS.n5804 VSS.n5803 1.13717
R22744 VSS.n6185 VSS.n6184 1.13717
R22745 VSS.n6226 VSS.n6225 1.13717
R22746 VSS.n6243 VSS.n6241 1.13717
R22747 VSS.n5733 VSS.n5732 1.13717
R22748 VSS.n5948 VSS.n5947 1.13717
R22749 VSS.n5946 VSS.n5927 1.13717
R22750 VSS.n5997 VSS.n5996 1.13717
R22751 VSS.n6004 VSS.n5900 1.13717
R22752 VSS.n5897 VSS.n5896 1.13717
R22753 VSS.n5879 VSS.n5878 1.13717
R22754 VSS.n6460 VSS.n6459 1.13717
R22755 VSS.n6458 VSS.n6445 1.13717
R22756 VSS.n6682 VSS.n6681 1.13717
R22757 VSS.n6428 VSS.n6424 1.13717
R22758 VSS.n6408 VSS.n6407 1.13717
R22759 VSS.n6396 VSS.n6395 1.13717
R22760 VSS.n6777 VSS.n6776 1.13717
R22761 VSS.n6818 VSS.n6817 1.13717
R22762 VSS.n6835 VSS.n6833 1.13717
R22763 VSS.n6325 VSS.n6324 1.13717
R22764 VSS.n6540 VSS.n6539 1.13717
R22765 VSS.n6538 VSS.n6519 1.13717
R22766 VSS.n6589 VSS.n6588 1.13717
R22767 VSS.n6596 VSS.n6492 1.13717
R22768 VSS.n6489 VSS.n6488 1.13717
R22769 VSS.n6471 VSS.n6470 1.13717
R22770 VSS.n7041 VSS.n7040 1.13717
R22771 VSS.n2497 VSS.n2495 1.13717
R22772 VSS.n2506 VSS.n2501 1.13717
R22773 VSS.n2517 VSS.n2515 1.13717
R22774 VSS.n2520 VSS.n2518 1.13717
R22775 VSS.n2526 VSS.n2524 1.13717
R22776 VSS.n2645 VSS.n2644 1.13717
R22777 VSS.n2688 VSS.n2687 1.13717
R22778 VSS.n2716 VSS.n2703 1.13717
R22779 VSS.n2770 VSS.n2753 1.13717
R22780 VSS.n2384 VSS.n2383 1.13717
R22781 VSS.n2382 VSS.n2363 1.13717
R22782 VSS.n2433 VSS.n2432 1.13717
R22783 VSS.n2440 VSS.n2336 1.13717
R22784 VSS.n2333 VSS.n2332 1.13717
R22785 VSS.n2315 VSS.n2314 1.13717
R22786 VSS.n2907 VSS.n2906 1.13717
R22787 VSS.n2905 VSS.n2892 1.13717
R22788 VSS.n3130 VSS.n3129 1.13717
R22789 VSS.n2875 VSS.n2871 1.13717
R22790 VSS.n2855 VSS.n2854 1.13717
R22791 VSS.n2843 VSS.n2842 1.13717
R22792 VSS.n3225 VSS.n3224 1.13717
R22793 VSS.n3266 VSS.n3265 1.13717
R22794 VSS.n3283 VSS.n3281 1.13717
R22795 VSS.n2772 VSS.n2771 1.13717
R22796 VSS.n2982 VSS.n2981 1.13717
R22797 VSS.n2980 VSS.n2969 1.13717
R22798 VSS.n3025 VSS.n3024 1.13717
R22799 VSS.n2950 VSS.n2946 1.13717
R22800 VSS.n2930 VSS.n2929 1.13717
R22801 VSS.n2918 VSS.n2917 1.13717
R22802 VSS.n174 VSS.n173 1.13717
R22803 VSS.n172 VSS.n159 1.13717
R22804 VSS.n9090 VSS.n9089 1.13717
R22805 VSS.n142 VSS.n138 1.13717
R22806 VSS.n122 VSS.n121 1.13717
R22807 VSS.n110 VSS.n109 1.13717
R22808 VSS.n9185 VSS.n9184 1.13717
R22809 VSS.n9226 VSS.n9225 1.13717
R22810 VSS.n9243 VSS.n9241 1.13717
R22811 VSS.n39 VSS.n38 1.13717
R22812 VSS.n432 VSS.n431 1.13717
R22813 VSS.n280 VSS.n278 1.13717
R22814 VSS.n289 VSS.n284 1.13717
R22815 VSS.n301 VSS.n299 1.13717
R22816 VSS.n304 VSS.n302 1.13717
R22817 VSS.n178 VSS.n177 1.13717
R22818 VSS.n36 VSS.n35 1.13717
R22819 VSS.n480 VSS.n479 1.13717
R22820 VSS.n486 VSS.n484 1.13717
R22821 VSS.n495 VSS.n490 1.13717
R22822 VSS.n506 VSS.n504 1.13717
R22823 VSS.n509 VSS.n507 1.13717
R22824 VSS.n515 VSS.n513 1.13717
R22825 VSS.n637 VSS.n636 1.13717
R22826 VSS.n680 VSS.n679 1.13717
R22827 VSS.n708 VSS.n695 1.13717
R22828 VSS.n997 VSS.n996 1.13717
R22829 VSS.n446 VSS.n444 1.13717
R22830 VSS.n455 VSS.n450 1.13717
R22831 VSS.n467 VSS.n465 1.13717
R22832 VSS.n470 VSS.n468 1.13717
R22833 VSS.n476 VSS.n474 1.13717
R22834 VSS.n8469 VSS.n8468 1.13717
R22835 VSS.n7065 VSS.n7063 1.13717
R22836 VSS.n7074 VSS.n7069 1.13717
R22837 VSS.n7085 VSS.n7083 1.13717
R22838 VSS.n7088 VSS.n7086 1.13717
R22839 VSS.n7094 VSS.n7092 1.13717
R22840 VSS.n7213 VSS.n7212 1.13717
R22841 VSS.n7256 VSS.n7255 1.13717
R22842 VSS.n7284 VSS.n7271 1.13717
R22843 VSS.n7338 VSS.n7321 1.13717
R22844 VSS.n7080 VSS.n7076 1.1255
R22845 VSS.n7535 VSS.n7447 1.1255
R22846 VSS.n8127 VSS.n7861 1.1255
R22847 VSS.n8659 VSS.n8655 1.1255
R22848 VSS.n1341 VSS.n1337 1.1255
R22849 VSS.n1914 VSS.n1910 1.1255
R22850 VSS.n3737 VSS.n3471 1.1255
R22851 VSS.n4329 VSS.n4063 1.1255
R22852 VSS.n4921 VSS.n4655 1.1255
R22853 VSS.n5513 VSS.n5247 1.1255
R22854 VSS.n6105 VSS.n5839 1.1255
R22855 VSS.n6697 VSS.n6431 1.1255
R22856 VSS.n2512 VSS.n2508 1.1255
R22857 VSS.n3145 VSS.n2878 1.1255
R22858 VSS.n9105 VSS.n145 1.1255
R22859 VSS.n501 VSS.n497 1.1255
R22860 VSS.n7595 VSS.n7401 1.09764
R22861 VSS.n7738 VSS.n7736 1.09764
R22862 VSS.n8187 VSS.n7815 1.09764
R22863 VSS.n8330 VSS.n8328 1.09764
R22864 VSS.n8991 VSS.n8990 1.09764
R22865 VSS.n8918 VSS.n8884 1.09764
R22866 VSS.n1654 VSS.n1653 1.09764
R22867 VSS.n1593 VSS.n1567 1.09764
R22868 VSS.n2246 VSS.n2245 1.09764
R22869 VSS.n2185 VSS.n2127 1.09764
R22870 VSS.n3797 VSS.n3425 1.09764
R22871 VSS.n3941 VSS.n3939 1.09764
R22872 VSS.n4389 VSS.n4017 1.09764
R22873 VSS.n4533 VSS.n4531 1.09764
R22874 VSS.n4981 VSS.n4609 1.09764
R22875 VSS.n5125 VSS.n5123 1.09764
R22876 VSS.n5573 VSS.n5201 1.09764
R22877 VSS.n5717 VSS.n5715 1.09764
R22878 VSS.n6165 VSS.n5793 1.09764
R22879 VSS.n6309 VSS.n6307 1.09764
R22880 VSS.n6757 VSS.n6385 1.09764
R22881 VSS.n6901 VSS.n6899 1.09764
R22882 VSS.n6990 VSS.n6989 1.09764
R22883 VSS.n6929 VSS.n2725 1.09764
R22884 VSS.n3205 VSS.n2832 1.09764
R22885 VSS.n3349 VSS.n3347 1.09764
R22886 VSS.n9165 VSS.n99 1.09764
R22887 VSS.n9309 VSS.n9307 1.09764
R22888 VSS.n809 VSS.n808 1.09764
R22889 VSS.n9331 VSS.n32 1.09764
R22890 VSS.n8418 VSS.n8417 1.09764
R22891 VSS.n8357 VSS.n7293 1.09764
R22892 VSS.n7378 VSS.n7376 1.04225
R22893 VSS.n7792 VSS.n7790 1.04225
R22894 VSS.n8819 VSS.n8817 1.04225
R22895 VSS.n1509 VSS.n1507 1.04225
R22896 VSS.n2082 VSS.n2080 1.04225
R22897 VSS.n3402 VSS.n3400 1.04225
R22898 VSS.n3994 VSS.n3992 1.04225
R22899 VSS.n4586 VSS.n4584 1.04225
R22900 VSS.n5178 VSS.n5176 1.04225
R22901 VSS.n5770 VSS.n5768 1.04225
R22902 VSS.n6362 VSS.n6360 1.04225
R22903 VSS.n2680 VSS.n2678 1.04225
R22904 VSS.n2809 VSS.n2807 1.04225
R22905 VSS.n76 VSS.n74 1.04225
R22906 VSS.n672 VSS.n670 1.04225
R22907 VSS.n7248 VSS.n7246 1.04225
R22908 VSS.n7122 VSS.n7059 1.00621
R22909 VSS.n7185 VSS.n7098 1.00621
R22910 VSS.n1072 VSS.n1007 1.00621
R22911 VSS.n1134 VSS.n1047 1.00621
R22912 VSS.n7629 VSS.n7401 1.00621
R22913 VSS.n7631 VSS.n7630 1.00621
R22914 VSS.n7679 VSS.n7678 1.00621
R22915 VSS.n7484 VSS.n7479 1.00621
R22916 VSS.n7580 VSS.n7415 1.00621
R22917 VSS.n7979 VSS.n7973 1.00621
R22918 VSS.n7915 VSS.n7904 1.00621
R22919 VSS.n8221 VSS.n7815 1.00621
R22920 VSS.n8223 VSS.n8222 1.00621
R22921 VSS.n8271 VSS.n8270 1.00621
R22922 VSS.n7898 VSS.n7893 1.00621
R22923 VSS.n8172 VSS.n7829 1.00621
R22924 VSS.n8701 VSS.n195 1.00621
R22925 VSS.n8764 VSS.n8677 1.00621
R22926 VSS.n8990 VSS.n8776 1.00621
R22927 VSS.n8828 VSS.n8827 1.00621
R22928 VSS.n8868 VSS.n8867 1.00621
R22929 VSS.n8540 VSS.n270 1.00621
R22930 VSS.n212 VSS.n201 1.00621
R22931 VSS.n1383 VSS.n1141 1.00621
R22932 VSS.n1446 VSS.n1359 1.00621
R22933 VSS.n1653 VSS.n1458 1.00621
R22934 VSS.n1646 VSS.n1645 1.00621
R22935 VSS.n1572 VSS.n1571 1.00621
R22936 VSS.n1222 VSS.n1216 1.00621
R22937 VSS.n1158 VSS.n1147 1.00621
R22938 VSS.n1956 VSS.n1714 1.00621
R22939 VSS.n2019 VSS.n1932 1.00621
R22940 VSS.n2245 VSS.n2031 1.00621
R22941 VSS.n2238 VSS.n2237 1.00621
R22942 VSS.n2132 VSS.n2131 1.00621
R22943 VSS.n1795 VSS.n1789 1.00621
R22944 VSS.n1731 VSS.n1720 1.00621
R22945 VSS.n3508 VSS.n3503 1.00621
R22946 VSS.n3782 VSS.n3439 1.00621
R22947 VSS.n3831 VSS.n3425 1.00621
R22948 VSS.n3833 VSS.n3832 1.00621
R22949 VSS.n3881 VSS.n3880 1.00621
R22950 VSS.n3589 VSS.n3583 1.00621
R22951 VSS.n3525 VSS.n3514 1.00621
R22952 VSS.n4100 VSS.n4095 1.00621
R22953 VSS.n4374 VSS.n4031 1.00621
R22954 VSS.n4423 VSS.n4017 1.00621
R22955 VSS.n4425 VSS.n4424 1.00621
R22956 VSS.n4473 VSS.n4472 1.00621
R22957 VSS.n4181 VSS.n4175 1.00621
R22958 VSS.n4117 VSS.n4106 1.00621
R22959 VSS.n4692 VSS.n4687 1.00621
R22960 VSS.n4966 VSS.n4623 1.00621
R22961 VSS.n5015 VSS.n4609 1.00621
R22962 VSS.n5017 VSS.n5016 1.00621
R22963 VSS.n5065 VSS.n5064 1.00621
R22964 VSS.n4773 VSS.n4767 1.00621
R22965 VSS.n4709 VSS.n4698 1.00621
R22966 VSS.n5284 VSS.n5279 1.00621
R22967 VSS.n5558 VSS.n5215 1.00621
R22968 VSS.n5607 VSS.n5201 1.00621
R22969 VSS.n5609 VSS.n5608 1.00621
R22970 VSS.n5657 VSS.n5656 1.00621
R22971 VSS.n5365 VSS.n5359 1.00621
R22972 VSS.n5301 VSS.n5290 1.00621
R22973 VSS.n5876 VSS.n5871 1.00621
R22974 VSS.n6150 VSS.n5807 1.00621
R22975 VSS.n6199 VSS.n5793 1.00621
R22976 VSS.n6201 VSS.n6200 1.00621
R22977 VSS.n6249 VSS.n6248 1.00621
R22978 VSS.n5957 VSS.n5951 1.00621
R22979 VSS.n5893 VSS.n5882 1.00621
R22980 VSS.n6468 VSS.n6463 1.00621
R22981 VSS.n6742 VSS.n6399 1.00621
R22982 VSS.n6791 VSS.n6385 1.00621
R22983 VSS.n6793 VSS.n6792 1.00621
R22984 VSS.n6841 VSS.n6840 1.00621
R22985 VSS.n6549 VSS.n6543 1.00621
R22986 VSS.n6485 VSS.n6474 1.00621
R22987 VSS.n2554 VSS.n2312 1.00621
R22988 VSS.n2617 VSS.n2530 1.00621
R22989 VSS.n6989 VSS.n2629 1.00621
R22990 VSS.n6982 VSS.n6981 1.00621
R22991 VSS.n2730 VSS.n2729 1.00621
R22992 VSS.n2393 VSS.n2387 1.00621
R22993 VSS.n2329 VSS.n2318 1.00621
R22994 VSS.n2915 VSS.n2910 1.00621
R22995 VSS.n3190 VSS.n2846 1.00621
R22996 VSS.n3239 VSS.n2832 1.00621
R22997 VSS.n3241 VSS.n3240 1.00621
R22998 VSS.n3289 VSS.n3288 1.00621
R22999 VSS.n2990 VSS.n2985 1.00621
R23000 VSS.n3086 VSS.n2921 1.00621
R23001 VSS.n187 VSS.n186 1.00621
R23002 VSS.n9150 VSS.n113 1.00621
R23003 VSS.n9199 VSS.n99 1.00621
R23004 VSS.n9201 VSS.n9200 1.00621
R23005 VSS.n9249 VSS.n9248 1.00621
R23006 VSS.n341 VSS.n274 1.00621
R23007 VSS.n387 VSS.n181 1.00621
R23008 VSS.n548 VSS.n541 1.00621
R23009 VSS.n609 VSS.n519 1.00621
R23010 VSS.n808 VSS.n621 1.00621
R23011 VSS.n801 VSS.n800 1.00621
R23012 VSS.n731 VSS.n730 1.00621
R23013 VSS.n891 VSS.n440 1.00621
R23014 VSS.n953 VSS.n866 1.00621
R23015 VSS.n8417 VSS.n7197 1.00621
R23016 VSS.n8410 VSS.n8409 1.00621
R23017 VSS.n7298 VSS.n7297 1.00621
R23018 VSS.n7601 VSS.n7586 0.914786
R23019 VSS.n7663 VSS.n7662 0.914786
R23020 VSS.n7664 VSS.n7374 0.914786
R23021 VSS.n7720 VSS.n7719 0.914786
R23022 VSS.n7736 VSS.n7349 0.914786
R23023 VSS.n7746 VSS.n7745 0.914786
R23024 VSS.n8193 VSS.n8178 0.914786
R23025 VSS.n8255 VSS.n8254 0.914786
R23026 VSS.n8256 VSS.n7788 0.914786
R23027 VSS.n8312 VSS.n8311 0.914786
R23028 VSS.n8328 VSS.n7763 0.914786
R23029 VSS.n8338 VSS.n8337 0.914786
R23030 VSS.n8997 VSS.n8770 0.914786
R23031 VSS.n8838 VSS.n8837 0.914786
R23032 VSS.n8962 VSS.n8820 0.914786
R23033 VSS.n8944 VSS.n8943 0.914786
R23034 VSS.n8942 VSS.n8884 0.914786
R23035 VSS.n8926 VSS.n8925 0.914786
R23036 VSS.n1660 VSS.n1452 0.914786
R23037 VSS.n1524 VSS.n1523 0.914786
R23038 VSS.n1525 VSS.n1505 0.914786
R23039 VSS.n1585 VSS.n1565 0.914786
R23040 VSS.n1594 VSS.n1593 0.914786
R23041 VSS.n9346 VSS.n9345 0.914786
R23042 VSS.n2252 VSS.n2025 0.914786
R23043 VSS.n2097 VSS.n2096 0.914786
R23044 VSS.n2098 VSS.n2078 0.914786
R23045 VSS.n2145 VSS.n2126 0.914786
R23046 VSS.n2186 VSS.n2185 0.914786
R23047 VSS.n2159 VSS.n2152 0.914786
R23048 VSS.n3803 VSS.n3788 0.914786
R23049 VSS.n3865 VSS.n3864 0.914786
R23050 VSS.n3866 VSS.n3398 0.914786
R23051 VSS.n3922 VSS.n3921 0.914786
R23052 VSS.n3939 VSS.n3374 0.914786
R23053 VSS.n3949 VSS.n3948 0.914786
R23054 VSS.n4395 VSS.n4380 0.914786
R23055 VSS.n4457 VSS.n4456 0.914786
R23056 VSS.n4458 VSS.n3990 0.914786
R23057 VSS.n4514 VSS.n4513 0.914786
R23058 VSS.n4531 VSS.n3966 0.914786
R23059 VSS.n4541 VSS.n4540 0.914786
R23060 VSS.n4987 VSS.n4972 0.914786
R23061 VSS.n5049 VSS.n5048 0.914786
R23062 VSS.n5050 VSS.n4582 0.914786
R23063 VSS.n5106 VSS.n5105 0.914786
R23064 VSS.n5123 VSS.n4558 0.914786
R23065 VSS.n5133 VSS.n5132 0.914786
R23066 VSS.n5579 VSS.n5564 0.914786
R23067 VSS.n5641 VSS.n5640 0.914786
R23068 VSS.n5642 VSS.n5174 0.914786
R23069 VSS.n5698 VSS.n5697 0.914786
R23070 VSS.n5715 VSS.n5150 0.914786
R23071 VSS.n5725 VSS.n5724 0.914786
R23072 VSS.n6171 VSS.n6156 0.914786
R23073 VSS.n6233 VSS.n6232 0.914786
R23074 VSS.n6234 VSS.n5766 0.914786
R23075 VSS.n6290 VSS.n6289 0.914786
R23076 VSS.n6307 VSS.n5742 0.914786
R23077 VSS.n6317 VSS.n6316 0.914786
R23078 VSS.n6763 VSS.n6748 0.914786
R23079 VSS.n6825 VSS.n6824 0.914786
R23080 VSS.n6826 VSS.n6358 0.914786
R23081 VSS.n6882 VSS.n6881 0.914786
R23082 VSS.n6899 VSS.n6334 0.914786
R23083 VSS.n6909 VSS.n6908 0.914786
R23084 VSS.n6996 VSS.n2623 0.914786
R23085 VSS.n2695 VSS.n2694 0.914786
R23086 VSS.n2696 VSS.n2676 0.914786
R23087 VSS.n2743 VSS.n2724 0.914786
R23088 VSS.n6930 VSS.n6929 0.914786
R23089 VSS.n2757 VSS.n2750 0.914786
R23090 VSS.n3211 VSS.n3196 0.914786
R23091 VSS.n3273 VSS.n3272 0.914786
R23092 VSS.n3274 VSS.n2805 0.914786
R23093 VSS.n3330 VSS.n3329 0.914786
R23094 VSS.n3347 VSS.n2781 0.914786
R23095 VSS.n3357 VSS.n3356 0.914786
R23096 VSS.n9171 VSS.n9156 0.914786
R23097 VSS.n9233 VSS.n9232 0.914786
R23098 VSS.n9234 VSS.n72 0.914786
R23099 VSS.n9290 VSS.n9289 0.914786
R23100 VSS.n9307 VSS.n48 0.914786
R23101 VSS.n9317 VSS.n9316 0.914786
R23102 VSS.n815 VSS.n615 0.914786
R23103 VSS.n687 VSS.n686 0.914786
R23104 VSS.n688 VSS.n668 0.914786
R23105 VSS.n748 VSS.n747 0.914786
R23106 VSS.n749 VSS.n32 0.914786
R23107 VSS.n9337 VSS.n27 0.914786
R23108 VSS.n8424 VSS.n7191 0.914786
R23109 VSS.n7263 VSS.n7262 0.914786
R23110 VSS.n7264 VSS.n7244 0.914786
R23111 VSS.n7311 VSS.n7292 0.914786
R23112 VSS.n8358 VSS.n8357 0.914786
R23113 VSS.n7325 VSS.n7318 0.914786
R23114 VSS.n7749 VSS.n7341 0.908949
R23115 VSS.n8341 VSS.n7755 0.908949
R23116 VSS.n8929 VSS.n8895 0.908949
R23117 VSS.n9349 VSS.n3 0.908949
R23118 VSS.n2175 VSS.n2160 0.908949
R23119 VSS.n3952 VSS.n3366 0.908949
R23120 VSS.n4544 VSS.n3958 0.908949
R23121 VSS.n5136 VSS.n4550 0.908949
R23122 VSS.n5728 VSS.n5142 0.908949
R23123 VSS.n6320 VSS.n5734 0.908949
R23124 VSS.n6912 VSS.n6326 0.908949
R23125 VSS.n6919 VSS.n2758 0.908949
R23126 VSS.n3360 VSS.n2773 0.908949
R23127 VSS.n9320 VSS.n40 0.908949
R23128 VSS.n9326 VSS.n28 0.908949
R23129 VSS.n8347 VSS.n7326 0.908949
R23130 VSS.n7589 VSS.n7410 0.908879
R23131 VSS.n8181 VSS.n7824 0.908879
R23132 VSS.n8789 VSS.n8771 0.908879
R23133 VSS.n1470 VSS.n1453 0.908879
R23134 VSS.n2043 VSS.n2026 0.908879
R23135 VSS.n3791 VSS.n3434 0.908879
R23136 VSS.n4383 VSS.n4026 0.908879
R23137 VSS.n4975 VSS.n4618 0.908879
R23138 VSS.n5567 VSS.n5210 0.908879
R23139 VSS.n6159 VSS.n5802 0.908879
R23140 VSS.n6751 VSS.n6394 0.908879
R23141 VSS.n2641 VSS.n2624 0.908879
R23142 VSS.n3199 VSS.n2841 0.908879
R23143 VSS.n9159 VSS.n108 0.908879
R23144 VSS.n633 VSS.n616 0.908879
R23145 VSS.n7209 VSS.n7192 0.908879
R23146 VSS.n7624 VSS.n7405 0.853
R23147 VSS.n7670 VSS.n7378 0.853
R23148 VSS.n7355 VSS.n7354 0.853
R23149 VSS.n8216 VSS.n7819 0.853
R23150 VSS.n8262 VSS.n7792 0.853
R23151 VSS.n7769 VSS.n7768 0.853
R23152 VSS.n8984 VSS.n8780 0.853
R23153 VSS.n8817 VSS.n8815 0.853
R23154 VSS.n8880 VSS.n8878 0.853
R23155 VSS.n1492 VSS.n1462 0.853
R23156 VSS.n1531 VSS.n1509 0.853
R23157 VSS.n1599 VSS.n1544 0.853
R23158 VSS.n2065 VSS.n2035 0.853
R23159 VSS.n2104 VSS.n2082 0.853
R23160 VSS.n2191 VSS.n2117 0.853
R23161 VSS.n3826 VSS.n3429 0.853
R23162 VSS.n3872 VSS.n3402 0.853
R23163 VSS.n3380 VSS.n3379 0.853
R23164 VSS.n4418 VSS.n4021 0.853
R23165 VSS.n4464 VSS.n3994 0.853
R23166 VSS.n3972 VSS.n3971 0.853
R23167 VSS.n5010 VSS.n4613 0.853
R23168 VSS.n5056 VSS.n4586 0.853
R23169 VSS.n4564 VSS.n4563 0.853
R23170 VSS.n5602 VSS.n5205 0.853
R23171 VSS.n5648 VSS.n5178 0.853
R23172 VSS.n5156 VSS.n5155 0.853
R23173 VSS.n6194 VSS.n5797 0.853
R23174 VSS.n6240 VSS.n5770 0.853
R23175 VSS.n5748 VSS.n5747 0.853
R23176 VSS.n6786 VSS.n6389 0.853
R23177 VSS.n6832 VSS.n6362 0.853
R23178 VSS.n6340 VSS.n6339 0.853
R23179 VSS.n2663 VSS.n2633 0.853
R23180 VSS.n2702 VSS.n2680 0.853
R23181 VSS.n6935 VSS.n2715 0.853
R23182 VSS.n3234 VSS.n2836 0.853
R23183 VSS.n3280 VSS.n2809 0.853
R23184 VSS.n2787 VSS.n2786 0.853
R23185 VSS.n9194 VSS.n103 0.853
R23186 VSS.n9240 VSS.n76 0.853
R23187 VSS.n54 VSS.n53 0.853
R23188 VSS.n655 VSS.n625 0.853
R23189 VSS.n694 VSS.n672 0.853
R23190 VSS.n754 VSS.n707 0.853
R23191 VSS.n7231 VSS.n7201 0.853
R23192 VSS.n7270 VSS.n7248 0.853
R23193 VSS.n8363 VSS.n7283 0.853
R23194 VSS.n7640 VSS.n7397 0.823357
R23195 VSS.n7649 VSS.n7389 0.823357
R23196 VSS.n7691 VSS.n7375 0.823357
R23197 VSS.n7701 VSS.n7362 0.823357
R23198 VSS.n8232 VSS.n7811 0.823357
R23199 VSS.n8241 VSS.n7803 0.823357
R23200 VSS.n8283 VSS.n7789 0.823357
R23201 VSS.n8293 VSS.n7776 0.823357
R23202 VSS.n8974 VSS.n8806 0.823357
R23203 VSS.n8973 VSS.n8972 0.823357
R23204 VSS.n8859 VSS.n8821 0.823357
R23205 VSS.n8904 VSS.n8850 0.823357
R23206 VSS.n1638 VSS.n1487 0.823357
R23207 VSS.n1630 VSS.n1499 0.823357
R23208 VSS.n1621 VSS.n1506 0.823357
R23209 VSS.n1610 VSS.n1609 0.823357
R23210 VSS.n2230 VSS.n2060 0.823357
R23211 VSS.n2222 VSS.n2072 0.823357
R23212 VSS.n2213 VSS.n2079 0.823357
R23213 VSS.n2202 VSS.n2201 0.823357
R23214 VSS.n3842 VSS.n3421 0.823357
R23215 VSS.n3851 VSS.n3413 0.823357
R23216 VSS.n3893 VSS.n3399 0.823357
R23217 VSS.n3903 VSS.n3386 0.823357
R23218 VSS.n4434 VSS.n4013 0.823357
R23219 VSS.n4443 VSS.n4005 0.823357
R23220 VSS.n4485 VSS.n3991 0.823357
R23221 VSS.n4495 VSS.n3978 0.823357
R23222 VSS.n5026 VSS.n4605 0.823357
R23223 VSS.n5035 VSS.n4597 0.823357
R23224 VSS.n5077 VSS.n4583 0.823357
R23225 VSS.n5087 VSS.n4570 0.823357
R23226 VSS.n5618 VSS.n5197 0.823357
R23227 VSS.n5627 VSS.n5189 0.823357
R23228 VSS.n5669 VSS.n5175 0.823357
R23229 VSS.n5679 VSS.n5162 0.823357
R23230 VSS.n6210 VSS.n5789 0.823357
R23231 VSS.n6219 VSS.n5781 0.823357
R23232 VSS.n6261 VSS.n5767 0.823357
R23233 VSS.n6271 VSS.n5754 0.823357
R23234 VSS.n6802 VSS.n6381 0.823357
R23235 VSS.n6811 VSS.n6373 0.823357
R23236 VSS.n6853 VSS.n6359 0.823357
R23237 VSS.n6863 VSS.n6346 0.823357
R23238 VSS.n6974 VSS.n2658 0.823357
R23239 VSS.n6966 VSS.n2670 0.823357
R23240 VSS.n6957 VSS.n2677 0.823357
R23241 VSS.n6946 VSS.n6945 0.823357
R23242 VSS.n3250 VSS.n2828 0.823357
R23243 VSS.n3259 VSS.n2820 0.823357
R23244 VSS.n3301 VSS.n2806 0.823357
R23245 VSS.n3311 VSS.n2793 0.823357
R23246 VSS.n9210 VSS.n95 0.823357
R23247 VSS.n9219 VSS.n87 0.823357
R23248 VSS.n9261 VSS.n73 0.823357
R23249 VSS.n9271 VSS.n60 0.823357
R23250 VSS.n793 VSS.n650 0.823357
R23251 VSS.n785 VSS.n662 0.823357
R23252 VSS.n776 VSS.n669 0.823357
R23253 VSS.n765 VSS.n764 0.823357
R23254 VSS.n8402 VSS.n7226 0.823357
R23255 VSS.n8394 VSS.n7238 0.823357
R23256 VSS.n8385 VSS.n7245 0.823357
R23257 VSS.n8374 VSS.n8373 0.823357
R23258 VSS.n7397 VSS.n7389 0.731929
R23259 VSS.n7701 VSS.n7700 0.731929
R23260 VSS.n7713 VSS.n7362 0.731929
R23261 VSS.n7811 VSS.n7803 0.731929
R23262 VSS.n8293 VSS.n8292 0.731929
R23263 VSS.n8305 VSS.n7776 0.731929
R23264 VSS.n8974 VSS.n8973 0.731929
R23265 VSS.n8953 VSS.n8850 0.731929
R23266 VSS.n8911 VSS.n8904 0.731929
R23267 VSS.n1499 VSS.n1487 0.731929
R23268 VSS.n1611 VSS.n1610 0.731929
R23269 VSS.n1609 VSS.n1538 0.731929
R23270 VSS.n2072 VSS.n2060 0.731929
R23271 VSS.n2203 VSS.n2202 0.731929
R23272 VSS.n2201 VSS.n2111 0.731929
R23273 VSS.n3421 VSS.n3413 0.731929
R23274 VSS.n3903 VSS.n3902 0.731929
R23275 VSS.n3915 VSS.n3386 0.731929
R23276 VSS.n4013 VSS.n4005 0.731929
R23277 VSS.n4495 VSS.n4494 0.731929
R23278 VSS.n4507 VSS.n3978 0.731929
R23279 VSS.n4605 VSS.n4597 0.731929
R23280 VSS.n5087 VSS.n5086 0.731929
R23281 VSS.n5099 VSS.n4570 0.731929
R23282 VSS.n5197 VSS.n5189 0.731929
R23283 VSS.n5679 VSS.n5678 0.731929
R23284 VSS.n5691 VSS.n5162 0.731929
R23285 VSS.n5789 VSS.n5781 0.731929
R23286 VSS.n6271 VSS.n6270 0.731929
R23287 VSS.n6283 VSS.n5754 0.731929
R23288 VSS.n6381 VSS.n6373 0.731929
R23289 VSS.n6863 VSS.n6862 0.731929
R23290 VSS.n6875 VSS.n6346 0.731929
R23291 VSS.n2670 VSS.n2658 0.731929
R23292 VSS.n6947 VSS.n6946 0.731929
R23293 VSS.n6945 VSS.n2709 0.731929
R23294 VSS.n2828 VSS.n2820 0.731929
R23295 VSS.n3311 VSS.n3310 0.731929
R23296 VSS.n3323 VSS.n2793 0.731929
R23297 VSS.n95 VSS.n87 0.731929
R23298 VSS.n9271 VSS.n9270 0.731929
R23299 VSS.n9283 VSS.n60 0.731929
R23300 VSS.n662 VSS.n650 0.731929
R23301 VSS.n766 VSS.n765 0.731929
R23302 VSS.n764 VSS.n701 0.731929
R23303 VSS.n7238 VSS.n7226 0.731929
R23304 VSS.n8375 VSS.n8374 0.731929
R23305 VSS.n8373 VSS.n7277 0.731929
R23306 VSS VSS.n3363 0.680647
R23307 VSS VSS.n0 0.680647
R23308 VSS.n7593 VSS.n7586 0.6405
R23309 VSS.n7662 VSS.n7383 0.6405
R23310 VSS.n7720 VSS.n7349 0.6405
R23311 VSS.n7746 VSS.n7343 0.6405
R23312 VSS.n8185 VSS.n8178 0.6405
R23313 VSS.n8254 VSS.n7797 0.6405
R23314 VSS.n8312 VSS.n7763 0.6405
R23315 VSS.n8338 VSS.n7757 0.6405
R23316 VSS.n8785 VSS.n8770 0.6405
R23317 VSS.n8842 VSS.n8837 0.6405
R23318 VSS.n8943 VSS.n8942 0.6405
R23319 VSS.n8926 VSS.n8898 0.6405
R23320 VSS.n1466 VSS.n1452 0.6405
R23321 VSS.n1523 VSS.n1501 0.6405
R23322 VSS.n1594 VSS.n1565 0.6405
R23323 VSS.n9346 VSS.n5 0.6405
R23324 VSS.n2039 VSS.n2025 0.6405
R23325 VSS.n2096 VSS.n2074 0.6405
R23326 VSS.n2186 VSS.n2126 0.6405
R23327 VSS.n2178 VSS.n2152 0.6405
R23328 VSS.n3795 VSS.n3788 0.6405
R23329 VSS.n3864 VSS.n3407 0.6405
R23330 VSS.n3922 VSS.n3374 0.6405
R23331 VSS.n3949 VSS.n3368 0.6405
R23332 VSS.n4387 VSS.n4380 0.6405
R23333 VSS.n4456 VSS.n3999 0.6405
R23334 VSS.n4514 VSS.n3966 0.6405
R23335 VSS.n4541 VSS.n3960 0.6405
R23336 VSS.n4979 VSS.n4972 0.6405
R23337 VSS.n5048 VSS.n4591 0.6405
R23338 VSS.n5106 VSS.n4558 0.6405
R23339 VSS.n5133 VSS.n4552 0.6405
R23340 VSS.n5571 VSS.n5564 0.6405
R23341 VSS.n5640 VSS.n5183 0.6405
R23342 VSS.n5698 VSS.n5150 0.6405
R23343 VSS.n5725 VSS.n5144 0.6405
R23344 VSS.n6163 VSS.n6156 0.6405
R23345 VSS.n6232 VSS.n5775 0.6405
R23346 VSS.n6290 VSS.n5742 0.6405
R23347 VSS.n6317 VSS.n5736 0.6405
R23348 VSS.n6755 VSS.n6748 0.6405
R23349 VSS.n6824 VSS.n6367 0.6405
R23350 VSS.n6882 VSS.n6334 0.6405
R23351 VSS.n6909 VSS.n6328 0.6405
R23352 VSS.n2637 VSS.n2623 0.6405
R23353 VSS.n2694 VSS.n2672 0.6405
R23354 VSS.n6930 VSS.n2724 0.6405
R23355 VSS.n6922 VSS.n2750 0.6405
R23356 VSS.n3203 VSS.n3196 0.6405
R23357 VSS.n3272 VSS.n2814 0.6405
R23358 VSS.n3330 VSS.n2781 0.6405
R23359 VSS.n3357 VSS.n2775 0.6405
R23360 VSS.n9163 VSS.n9156 0.6405
R23361 VSS.n9232 VSS.n81 0.6405
R23362 VSS.n9290 VSS.n48 0.6405
R23363 VSS.n9317 VSS.n42 0.6405
R23364 VSS.n629 VSS.n615 0.6405
R23365 VSS.n686 VSS.n664 0.6405
R23366 VSS.n749 VSS.n748 0.6405
R23367 VSS.n9329 VSS.n27 0.6405
R23368 VSS.n7205 VSS.n7191 0.6405
R23369 VSS.n7262 VSS.n7240 0.6405
R23370 VSS.n8358 VSS.n7292 0.6405
R23371 VSS.n8350 VSS.n7318 0.6405
R23372 VSS.n7630 VSS.n7629 0.549071
R23373 VSS.n7679 VSS.n7370 0.549071
R23374 VSS.n8222 VSS.n8221 0.549071
R23375 VSS.n8271 VSS.n7784 0.549071
R23376 VSS.n8827 VSS.n8776 0.549071
R23377 VSS.n8868 VSS.n8849 0.549071
R23378 VSS.n1646 VSS.n1458 0.549071
R23379 VSS.n1578 VSS.n1571 0.549071
R23380 VSS.n2238 VSS.n2031 0.549071
R23381 VSS.n2138 VSS.n2131 0.549071
R23382 VSS.n3832 VSS.n3831 0.549071
R23383 VSS.n3881 VSS.n3394 0.549071
R23384 VSS.n4424 VSS.n4423 0.549071
R23385 VSS.n4473 VSS.n3986 0.549071
R23386 VSS.n5016 VSS.n5015 0.549071
R23387 VSS.n5065 VSS.n4578 0.549071
R23388 VSS.n5608 VSS.n5607 0.549071
R23389 VSS.n5657 VSS.n5170 0.549071
R23390 VSS.n6200 VSS.n6199 0.549071
R23391 VSS.n6249 VSS.n5762 0.549071
R23392 VSS.n6792 VSS.n6791 0.549071
R23393 VSS.n6841 VSS.n6354 0.549071
R23394 VSS.n6982 VSS.n2629 0.549071
R23395 VSS.n2736 VSS.n2729 0.549071
R23396 VSS.n3240 VSS.n3239 0.549071
R23397 VSS.n3289 VSS.n2801 0.549071
R23398 VSS.n9200 VSS.n9199 0.549071
R23399 VSS.n9249 VSS.n68 0.549071
R23400 VSS.n801 VSS.n621 0.549071
R23401 VSS.n737 VSS.n730 0.549071
R23402 VSS.n8410 VSS.n7197 0.549071
R23403 VSS.n7304 VSS.n7297 0.549071
R23404 VSS.n7613 VSS 0.517836
R23405 VSS.n8205 VSS 0.517836
R23406 VSS.n8791 VSS 0.517836
R23407 VSS.n1472 VSS 0.517836
R23408 VSS.n2045 VSS 0.517836
R23409 VSS.n3815 VSS 0.517836
R23410 VSS.n4407 VSS 0.517836
R23411 VSS.n4999 VSS 0.517836
R23412 VSS.n5591 VSS 0.517836
R23413 VSS.n6183 VSS 0.517836
R23414 VSS.n6775 VSS 0.517836
R23415 VSS.n2643 VSS 0.517836
R23416 VSS.n3223 VSS 0.517836
R23417 VSS.n9183 VSS 0.517836
R23418 VSS.n635 VSS 0.517836
R23419 VSS.n7211 VSS 0.517836
R23420 VSS.n8472 VSS.n7059 0.465127
R23421 VSS.n8521 VSS.n1007 0.465127
R23422 VSS.n7485 VSS.n7484 0.465127
R23423 VSS.n7980 VSS.n7979 0.465127
R23424 VSS.n7899 VSS.n7898 0.465127
R23425 VSS.n9045 VSS.n195 0.465127
R23426 VSS.n8541 VSS.n8540 0.465127
R23427 VSS.n1708 VSS.n1141 0.465127
R23428 VSS.n1223 VSS.n1222 0.465127
R23429 VSS.n2300 VSS.n1714 0.465127
R23430 VSS.n1796 VSS.n1795 0.465127
R23431 VSS.n3509 VSS.n3508 0.465127
R23432 VSS.n3590 VSS.n3589 0.465127
R23433 VSS.n4101 VSS.n4100 0.465127
R23434 VSS.n4182 VSS.n4181 0.465127
R23435 VSS.n4693 VSS.n4692 0.465127
R23436 VSS.n4774 VSS.n4773 0.465127
R23437 VSS.n5285 VSS.n5284 0.465127
R23438 VSS.n5366 VSS.n5365 0.465127
R23439 VSS.n5877 VSS.n5876 0.465127
R23440 VSS.n5958 VSS.n5957 0.465127
R23441 VSS.n6469 VSS.n6468 0.465127
R23442 VSS.n6550 VSS.n6549 0.465127
R23443 VSS.n7044 VSS.n2312 0.465127
R23444 VSS.n2394 VSS.n2393 0.465127
R23445 VSS.n2916 VSS.n2915 0.465127
R23446 VSS.n2991 VSS.n2990 0.465127
R23447 VSS.n187 VSS.n176 0.465127
R23448 VSS.n435 VSS.n274 0.465127
R23449 VSS.n541 VSS.n481 0.465127
R23450 VSS.n1000 VSS.n440 0.465127
R23451 VSS.n8432 VSS.n7098 0.457643
R23452 VSS.n8481 VSS.n1047 0.457643
R23453 VSS.n7595 VSS.n7594 0.457643
R23454 VSS.n7738 VSS.n7737 0.457643
R23455 VSS.n7609 VSS.n7415 0.457643
R23456 VSS.n8075 VSS.n7904 0.457643
R23457 VSS.n8187 VSS.n8186 0.457643
R23458 VSS.n8330 VSS.n8329 0.457643
R23459 VSS.n8201 VSS.n7829 0.457643
R23460 VSS.n9005 VSS.n8677 0.457643
R23461 VSS.n8991 VSS.n8775 0.457643
R23462 VSS.n8918 VSS.n8917 0.457643
R23463 VSS.n8636 VSS.n201 0.457643
R23464 VSS.n1668 VSS.n1359 0.457643
R23465 VSS.n1654 VSS.n1457 0.457643
R23466 VSS.n1567 VSS.n1566 0.457643
R23467 VSS.n1318 VSS.n1147 0.457643
R23468 VSS.n2260 VSS.n1932 0.457643
R23469 VSS.n2246 VSS.n2030 0.457643
R23470 VSS.n2179 VSS.n2127 0.457643
R23471 VSS.n1891 VSS.n1720 0.457643
R23472 VSS.n3811 VSS.n3439 0.457643
R23473 VSS.n3797 VSS.n3796 0.457643
R23474 VSS.n3941 VSS.n3940 0.457643
R23475 VSS.n3685 VSS.n3514 0.457643
R23476 VSS.n4403 VSS.n4031 0.457643
R23477 VSS.n4389 VSS.n4388 0.457643
R23478 VSS.n4533 VSS.n4532 0.457643
R23479 VSS.n4277 VSS.n4106 0.457643
R23480 VSS.n4995 VSS.n4623 0.457643
R23481 VSS.n4981 VSS.n4980 0.457643
R23482 VSS.n5125 VSS.n5124 0.457643
R23483 VSS.n4869 VSS.n4698 0.457643
R23484 VSS.n5587 VSS.n5215 0.457643
R23485 VSS.n5573 VSS.n5572 0.457643
R23486 VSS.n5717 VSS.n5716 0.457643
R23487 VSS.n5461 VSS.n5290 0.457643
R23488 VSS.n6179 VSS.n5807 0.457643
R23489 VSS.n6165 VSS.n6164 0.457643
R23490 VSS.n6309 VSS.n6308 0.457643
R23491 VSS.n6053 VSS.n5882 0.457643
R23492 VSS.n6771 VSS.n6399 0.457643
R23493 VSS.n6757 VSS.n6756 0.457643
R23494 VSS.n6901 VSS.n6900 0.457643
R23495 VSS.n6645 VSS.n6474 0.457643
R23496 VSS.n7004 VSS.n2530 0.457643
R23497 VSS.n6990 VSS.n2628 0.457643
R23498 VSS.n6923 VSS.n2725 0.457643
R23499 VSS.n2489 VSS.n2318 0.457643
R23500 VSS.n3219 VSS.n2846 0.457643
R23501 VSS.n3205 VSS.n3204 0.457643
R23502 VSS.n3349 VSS.n3348 0.457643
R23503 VSS.n3093 VSS.n2921 0.457643
R23504 VSS.n9179 VSS.n113 0.457643
R23505 VSS.n9165 VSS.n9164 0.457643
R23506 VSS.n9309 VSS.n9308 0.457643
R23507 VSS.n9053 VSS.n181 0.457643
R23508 VSS.n823 VSS.n519 0.457643
R23509 VSS.n809 VSS.n620 0.457643
R23510 VSS.n9331 VSS.n9330 0.457643
R23511 VSS.n960 VSS.n866 0.457643
R23512 VSS.n8418 VSS.n7196 0.457643
R23513 VSS.n8351 VSS.n7293 0.457643
R23514 VSS.n9324 VSS 0.415989
R23515 VSS.n6916 VSS 0.415941
R23516 VSS.n5139 VSS 0.415941
R23517 VSS.n9352 VSS 0.415941
R23518 VSS.n5731 VSS 0.382853
R23519 VSS.n7144 VSS.n7135 0.366214
R23520 VSS.n7175 VSS.n7174 0.366214
R23521 VSS.n1092 VSS.n1085 0.366214
R23522 VSS.n1124 VSS.n1123 0.366214
R23523 VSS.n7505 VSS.n7466 0.366214
R23524 VSS.n7565 VSS.n7563 0.366214
R23525 VSS.n8001 VSS.n7999 0.366214
R23526 VSS.n8067 VSS.n7907 0.366214
R23527 VSS.n8097 VSS.n7880 0.366214
R23528 VSS.n8157 VSS.n8155 0.366214
R23529 VSS.n8723 VSS.n8714 0.366214
R23530 VSS.n8754 VSS.n8753 0.366214
R23531 VSS.n8562 VSS.n8560 0.366214
R23532 VSS.n8628 VSS.n204 0.366214
R23533 VSS.n1405 VSS.n1396 0.366214
R23534 VSS.n1436 VSS.n1435 0.366214
R23535 VSS.n1244 VSS.n1242 0.366214
R23536 VSS.n1310 VSS.n1150 0.366214
R23537 VSS.n1978 VSS.n1969 0.366214
R23538 VSS.n2009 VSS.n2008 0.366214
R23539 VSS.n1817 VSS.n1815 0.366214
R23540 VSS.n1883 VSS.n1723 0.366214
R23541 VSS.n3707 VSS.n3490 0.366214
R23542 VSS.n3767 VSS.n3765 0.366214
R23543 VSS.n3611 VSS.n3609 0.366214
R23544 VSS.n3677 VSS.n3517 0.366214
R23545 VSS.n4299 VSS.n4082 0.366214
R23546 VSS.n4359 VSS.n4357 0.366214
R23547 VSS.n4203 VSS.n4201 0.366214
R23548 VSS.n4269 VSS.n4109 0.366214
R23549 VSS.n4891 VSS.n4674 0.366214
R23550 VSS.n4951 VSS.n4949 0.366214
R23551 VSS.n4795 VSS.n4793 0.366214
R23552 VSS.n4861 VSS.n4701 0.366214
R23553 VSS.n5483 VSS.n5266 0.366214
R23554 VSS.n5543 VSS.n5541 0.366214
R23555 VSS.n5387 VSS.n5385 0.366214
R23556 VSS.n5453 VSS.n5293 0.366214
R23557 VSS.n6075 VSS.n5858 0.366214
R23558 VSS.n6135 VSS.n6133 0.366214
R23559 VSS.n5979 VSS.n5977 0.366214
R23560 VSS.n6045 VSS.n5885 0.366214
R23561 VSS.n6667 VSS.n6450 0.366214
R23562 VSS.n6727 VSS.n6725 0.366214
R23563 VSS.n6571 VSS.n6569 0.366214
R23564 VSS.n6637 VSS.n6477 0.366214
R23565 VSS.n2576 VSS.n2567 0.366214
R23566 VSS.n2607 VSS.n2606 0.366214
R23567 VSS.n2415 VSS.n2413 0.366214
R23568 VSS.n2481 VSS.n2321 0.366214
R23569 VSS.n3115 VSS.n2897 0.366214
R23570 VSS.n3175 VSS.n3173 0.366214
R23571 VSS.n3010 VSS.n2972 0.366214
R23572 VSS.n3071 VSS.n3069 0.366214
R23573 VSS.n9075 VSS.n164 0.366214
R23574 VSS.n9135 VSS.n9133 0.366214
R23575 VSS.n347 VSS.n327 0.366214
R23576 VSS.n381 VSS.n380 0.366214
R23577 VSS.n568 VSS.n559 0.366214
R23578 VSS.n599 VSS.n598 0.366214
R23579 VSS.n911 VSS.n904 0.366214
R23580 VSS.n943 VSS.n942 0.366214
R23581 VSS.n1009 VSS 0.301636
R23582 VSS.n7981 VSS 0.301636
R23583 VSS.n8542 VSS 0.301636
R23584 VSS.n1224 VSS 0.301636
R23585 VSS.n1797 VSS 0.301636
R23586 VSS.n3591 VSS 0.301636
R23587 VSS.n4183 VSS 0.301636
R23588 VSS.n4775 VSS 0.301636
R23589 VSS.n5367 VSS 0.301636
R23590 VSS.n5959 VSS 0.301636
R23591 VSS.n6551 VSS 0.301636
R23592 VSS.n2395 VSS 0.301636
R23593 VSS.n2992 VSS 0.301636
R23594 VSS.n276 VSS 0.301636
R23595 VSS.n442 VSS 0.301636
R23596 VSS.n7061 VSS 0.301636
R23597 VSS VSS.n7750 0.300964
R23598 VSS VSS.n8342 0.300964
R23599 VSS.n8893 VSS 0.300964
R23600 VSS VSS.n9350 0.300964
R23601 VSS.n2174 VSS 0.300964
R23602 VSS VSS.n3953 0.300964
R23603 VSS VSS.n4545 0.300964
R23604 VSS VSS.n5137 0.300964
R23605 VSS VSS.n5729 0.300964
R23606 VSS VSS.n6321 0.300964
R23607 VSS VSS.n6913 0.300964
R23608 VSS.n6918 VSS 0.300964
R23609 VSS VSS.n3361 0.300964
R23610 VSS VSS.n9321 0.300964
R23611 VSS.n9325 VSS 0.300964
R23612 VSS.n8346 VSS 0.300964
R23613 VSS.n7487 VSS 0.29425
R23614 VSS.n8079 VSS 0.29425
R23615 VSS.n8640 VSS 0.29425
R23616 VSS.n1322 VSS 0.29425
R23617 VSS.n1895 VSS 0.29425
R23618 VSS.n3689 VSS 0.29425
R23619 VSS.n4281 VSS 0.29425
R23620 VSS.n4873 VSS 0.29425
R23621 VSS.n5465 VSS 0.29425
R23622 VSS.n6057 VSS 0.29425
R23623 VSS.n6649 VSS 0.29425
R23624 VSS.n2493 VSS 0.29425
R23625 VSS.n3097 VSS 0.29425
R23626 VSS.n9057 VSS 0.29425
R23627 VSS VSS.n863 0.29425
R23628 VSS.n7641 VSS.n7396 0.274786
R23629 VSS.n7664 VSS.n7663 0.274786
R23630 VSS.n7678 VSS.n7375 0.274786
R23631 VSS.n7718 VSS.n7358 0.274786
R23632 VSS.n8233 VSS.n7810 0.274786
R23633 VSS.n8256 VSS.n8255 0.274786
R23634 VSS.n8270 VSS.n7789 0.274786
R23635 VSS.n8310 VSS.n7772 0.274786
R23636 VSS.n8830 VSS.n8829 0.274786
R23637 VSS.n8838 VSS.n8820 0.274786
R23638 VSS.n8867 VSS.n8859 0.274786
R23639 VSS.n8905 VSS.n8883 0.274786
R23640 VSS.n1644 VSS.n1483 0.274786
R23641 VSS.n1525 VSS.n1524 0.274786
R23642 VSS.n1572 VSS.n1506 0.274786
R23643 VSS.n1587 VSS.n1586 0.274786
R23644 VSS.n2236 VSS.n2056 0.274786
R23645 VSS.n2098 VSS.n2097 0.274786
R23646 VSS.n2132 VSS.n2079 0.274786
R23647 VSS.n2147 VSS.n2146 0.274786
R23648 VSS.n3843 VSS.n3420 0.274786
R23649 VSS.n3866 VSS.n3865 0.274786
R23650 VSS.n3880 VSS.n3399 0.274786
R23651 VSS.n3920 VSS.n3382 0.274786
R23652 VSS.n4435 VSS.n4012 0.274786
R23653 VSS.n4458 VSS.n4457 0.274786
R23654 VSS.n4472 VSS.n3991 0.274786
R23655 VSS.n4512 VSS.n3974 0.274786
R23656 VSS.n5027 VSS.n4604 0.274786
R23657 VSS.n5050 VSS.n5049 0.274786
R23658 VSS.n5064 VSS.n4583 0.274786
R23659 VSS.n5104 VSS.n4566 0.274786
R23660 VSS.n5619 VSS.n5196 0.274786
R23661 VSS.n5642 VSS.n5641 0.274786
R23662 VSS.n5656 VSS.n5175 0.274786
R23663 VSS.n5696 VSS.n5158 0.274786
R23664 VSS.n6211 VSS.n5788 0.274786
R23665 VSS.n6234 VSS.n6233 0.274786
R23666 VSS.n6248 VSS.n5767 0.274786
R23667 VSS.n6288 VSS.n5750 0.274786
R23668 VSS.n6803 VSS.n6380 0.274786
R23669 VSS.n6826 VSS.n6825 0.274786
R23670 VSS.n6840 VSS.n6359 0.274786
R23671 VSS.n6880 VSS.n6342 0.274786
R23672 VSS.n6980 VSS.n2654 0.274786
R23673 VSS.n2696 VSS.n2695 0.274786
R23674 VSS.n2730 VSS.n2677 0.274786
R23675 VSS.n2745 VSS.n2744 0.274786
R23676 VSS.n3251 VSS.n2827 0.274786
R23677 VSS.n3274 VSS.n3273 0.274786
R23678 VSS.n3288 VSS.n2806 0.274786
R23679 VSS.n3328 VSS.n2789 0.274786
R23680 VSS.n9211 VSS.n94 0.274786
R23681 VSS.n9234 VSS.n9233 0.274786
R23682 VSS.n9248 VSS.n73 0.274786
R23683 VSS.n9288 VSS.n56 0.274786
R23684 VSS.n799 VSS.n646 0.274786
R23685 VSS.n688 VSS.n687 0.274786
R23686 VSS.n731 VSS.n669 0.274786
R23687 VSS.n746 VSS.n727 0.274786
R23688 VSS.n8408 VSS.n7222 0.274786
R23689 VSS.n7264 VSS.n7263 0.274786
R23690 VSS.n7298 VSS.n7245 0.274786
R23691 VSS.n7313 VSS.n7312 0.274786
R23692 VSS VSS.n7486 0.206964
R23693 VSS VSS.n8078 0.206964
R23694 VSS VSS.n8639 0.206964
R23695 VSS VSS.n1321 0.206964
R23696 VSS VSS.n1894 0.206964
R23697 VSS VSS.n3688 0.206964
R23698 VSS VSS.n4280 0.206964
R23699 VSS VSS.n4872 0.206964
R23700 VSS VSS.n5464 0.206964
R23701 VSS VSS.n6056 0.206964
R23702 VSS VSS.n6648 0.206964
R23703 VSS VSS.n2492 0.206964
R23704 VSS VSS.n3096 0.206964
R23705 VSS VSS.n9056 0.206964
R23706 VSS.n864 VSS 0.206964
R23707 VSS.n7150 VSS.n7115 0.183357
R23708 VSS.n7151 VSS.n7150 0.183357
R23709 VSS.n7169 VSS.n7159 0.183357
R23710 VSS.n7169 VSS.n7160 0.183357
R23711 VSS.n1098 VSS.n1065 0.183357
R23712 VSS.n1099 VSS.n1098 0.183357
R23713 VSS.n1117 VSS.n1107 0.183357
R23714 VSS.n1117 VSS.n1108 0.183357
R23715 VSS.n7526 VSS.n7455 0.183357
R23716 VSS.n7527 VSS.n7526 0.183357
R23717 VSS.n7558 VSS.n7434 0.183357
R23718 VSS.n7558 VSS.n7435 0.183357
R23719 VSS.n8011 VSS.n8010 0.183357
R23720 VSS.n8010 VSS.n7957 0.183357
R23721 VSS.n8043 VSS.n7927 0.183357
R23722 VSS.n8043 VSS.n7928 0.183357
R23723 VSS.n8118 VSS.n7869 0.183357
R23724 VSS.n8119 VSS.n8118 0.183357
R23725 VSS.n8150 VSS.n7848 0.183357
R23726 VSS.n8150 VSS.n7849 0.183357
R23727 VSS.n8729 VSS.n8694 0.183357
R23728 VSS.n8730 VSS.n8729 0.183357
R23729 VSS.n8748 VSS.n8738 0.183357
R23730 VSS.n8748 VSS.n8739 0.183357
R23731 VSS.n8572 VSS.n8571 0.183357
R23732 VSS.n8571 VSS.n254 0.183357
R23733 VSS.n8604 VSS.n224 0.183357
R23734 VSS.n8604 VSS.n225 0.183357
R23735 VSS.n1411 VSS.n1376 0.183357
R23736 VSS.n1412 VSS.n1411 0.183357
R23737 VSS.n1430 VSS.n1420 0.183357
R23738 VSS.n1430 VSS.n1421 0.183357
R23739 VSS.n1254 VSS.n1253 0.183357
R23740 VSS.n1253 VSS.n1200 0.183357
R23741 VSS.n1286 VSS.n1170 0.183357
R23742 VSS.n1286 VSS.n1171 0.183357
R23743 VSS.n1984 VSS.n1949 0.183357
R23744 VSS.n1985 VSS.n1984 0.183357
R23745 VSS.n2003 VSS.n1993 0.183357
R23746 VSS.n2003 VSS.n1994 0.183357
R23747 VSS.n1827 VSS.n1826 0.183357
R23748 VSS.n1826 VSS.n1773 0.183357
R23749 VSS.n1859 VSS.n1743 0.183357
R23750 VSS.n1859 VSS.n1744 0.183357
R23751 VSS.n3728 VSS.n3479 0.183357
R23752 VSS.n3729 VSS.n3728 0.183357
R23753 VSS.n3760 VSS.n3458 0.183357
R23754 VSS.n3760 VSS.n3459 0.183357
R23755 VSS.n3621 VSS.n3620 0.183357
R23756 VSS.n3620 VSS.n3567 0.183357
R23757 VSS.n3653 VSS.n3537 0.183357
R23758 VSS.n3653 VSS.n3538 0.183357
R23759 VSS.n4320 VSS.n4071 0.183357
R23760 VSS.n4321 VSS.n4320 0.183357
R23761 VSS.n4352 VSS.n4050 0.183357
R23762 VSS.n4352 VSS.n4051 0.183357
R23763 VSS.n4213 VSS.n4212 0.183357
R23764 VSS.n4212 VSS.n4159 0.183357
R23765 VSS.n4245 VSS.n4129 0.183357
R23766 VSS.n4245 VSS.n4130 0.183357
R23767 VSS.n4912 VSS.n4663 0.183357
R23768 VSS.n4913 VSS.n4912 0.183357
R23769 VSS.n4944 VSS.n4642 0.183357
R23770 VSS.n4944 VSS.n4643 0.183357
R23771 VSS.n4805 VSS.n4804 0.183357
R23772 VSS.n4804 VSS.n4751 0.183357
R23773 VSS.n4837 VSS.n4721 0.183357
R23774 VSS.n4837 VSS.n4722 0.183357
R23775 VSS.n5504 VSS.n5255 0.183357
R23776 VSS.n5505 VSS.n5504 0.183357
R23777 VSS.n5536 VSS.n5234 0.183357
R23778 VSS.n5536 VSS.n5235 0.183357
R23779 VSS.n5397 VSS.n5396 0.183357
R23780 VSS.n5396 VSS.n5343 0.183357
R23781 VSS.n5429 VSS.n5313 0.183357
R23782 VSS.n5429 VSS.n5314 0.183357
R23783 VSS.n6096 VSS.n5847 0.183357
R23784 VSS.n6097 VSS.n6096 0.183357
R23785 VSS.n6128 VSS.n5826 0.183357
R23786 VSS.n6128 VSS.n5827 0.183357
R23787 VSS.n5989 VSS.n5988 0.183357
R23788 VSS.n5988 VSS.n5935 0.183357
R23789 VSS.n6021 VSS.n5905 0.183357
R23790 VSS.n6021 VSS.n5906 0.183357
R23791 VSS.n6688 VSS.n6439 0.183357
R23792 VSS.n6689 VSS.n6688 0.183357
R23793 VSS.n6720 VSS.n6418 0.183357
R23794 VSS.n6720 VSS.n6419 0.183357
R23795 VSS.n6581 VSS.n6580 0.183357
R23796 VSS.n6580 VSS.n6527 0.183357
R23797 VSS.n6613 VSS.n6497 0.183357
R23798 VSS.n6613 VSS.n6498 0.183357
R23799 VSS.n2582 VSS.n2547 0.183357
R23800 VSS.n2583 VSS.n2582 0.183357
R23801 VSS.n2601 VSS.n2591 0.183357
R23802 VSS.n2601 VSS.n2592 0.183357
R23803 VSS.n2425 VSS.n2424 0.183357
R23804 VSS.n2424 VSS.n2371 0.183357
R23805 VSS.n2457 VSS.n2341 0.183357
R23806 VSS.n2457 VSS.n2342 0.183357
R23807 VSS.n3136 VSS.n2886 0.183357
R23808 VSS.n3137 VSS.n3136 0.183357
R23809 VSS.n3168 VSS.n2865 0.183357
R23810 VSS.n3168 VSS.n2866 0.183357
R23811 VSS.n3031 VSS.n2963 0.183357
R23812 VSS.n3032 VSS.n3031 0.183357
R23813 VSS.n3063 VSS.n2940 0.183357
R23814 VSS.n3063 VSS.n2941 0.183357
R23815 VSS.n9096 VSS.n153 0.183357
R23816 VSS.n9097 VSS.n9096 0.183357
R23817 VSS.n9128 VSS.n132 0.183357
R23818 VSS.n9128 VSS.n133 0.183357
R23819 VSS.n355 VSS.n326 0.183357
R23820 VSS.n355 VSS.n322 0.183357
R23821 VSS.n370 VSS.n318 0.183357
R23822 VSS.n370 VSS.n316 0.183357
R23823 VSS.n574 VSS.n536 0.183357
R23824 VSS.n575 VSS.n574 0.183357
R23825 VSS.n593 VSS.n583 0.183357
R23826 VSS.n593 VSS.n584 0.183357
R23827 VSS.n917 VSS.n884 0.183357
R23828 VSS.n918 VSS.n917 0.183357
R23829 VSS.n936 VSS.n926 0.183357
R23830 VSS.n936 VSS.n927 0.183357
R23831 VSS.n7751 VSS 0.107929
R23832 VSS.n8343 VSS 0.107929
R23833 VSS VSS.n8892 0.107929
R23834 VSS.n9351 VSS 0.107929
R23835 VSS VSS.n2173 0.107929
R23836 VSS.n3954 VSS 0.107929
R23837 VSS.n4546 VSS 0.107929
R23838 VSS.n5138 VSS 0.107929
R23839 VSS.n5730 VSS 0.107929
R23840 VSS.n6322 VSS 0.107929
R23841 VSS.n6914 VSS 0.107929
R23842 VSS VSS.n6917 0.107929
R23843 VSS.n3362 VSS 0.107929
R23844 VSS.n9322 VSS 0.107929
R23845 VSS VSS.n9324 0.107929
R23846 VSS VSS.n8345 0.107929
R23847 VSS VSS.n7612 0.107593
R23848 VSS VSS.n8204 0.107593
R23849 VSS VSS.n8790 0.107593
R23850 VSS VSS.n1471 0.107593
R23851 VSS VSS.n2044 0.107593
R23852 VSS VSS.n3814 0.107593
R23853 VSS VSS.n4406 0.107593
R23854 VSS VSS.n4998 0.107593
R23855 VSS VSS.n5590 0.107593
R23856 VSS VSS.n6182 0.107593
R23857 VSS VSS.n6774 0.107593
R23858 VSS VSS.n2642 0.107593
R23859 VSS VSS.n3222 0.107593
R23860 VSS VSS.n9182 0.107593
R23861 VSS VSS.n634 0.107593
R23862 VSS VSS.n7210 0.107593
R23863 VSS.n7176 VSS.n7175 0.0919286
R23864 VSS.n7184 VSS.n7102 0.0919286
R23865 VSS.n8432 VSS.n8431 0.0919286
R23866 VSS.n1125 VSS.n1124 0.0919286
R23867 VSS.n1133 VSS.n1051 0.0919286
R23868 VSS.n8481 VSS.n8480 0.0919286
R23869 VSS.n7648 VSS.n7391 0.0919286
R23870 VSS.n7699 VSS.n7698 0.0919286
R23871 VSS.n7565 VSS.n7564 0.0919286
R23872 VSS.n7579 VSS.n7419 0.0919286
R23873 VSS.n7609 VSS.n7608 0.0919286
R23874 VSS.n8067 VSS.n7908 0.0919286
R23875 VSS.n7916 VSS.n7914 0.0919286
R23876 VSS.n8075 VSS.n8074 0.0919286
R23877 VSS.n8240 VSS.n7805 0.0919286
R23878 VSS.n8291 VSS.n8290 0.0919286
R23879 VSS.n8157 VSS.n8156 0.0919286
R23880 VSS.n8171 VSS.n7833 0.0919286
R23881 VSS.n8201 VSS.n8200 0.0919286
R23882 VSS.n8755 VSS.n8754 0.0919286
R23883 VSS.n8763 VSS.n8681 0.0919286
R23884 VSS.n9005 VSS.n9004 0.0919286
R23885 VSS.n8843 VSS.n8807 0.0919286
R23886 VSS.n8955 VSS.n8954 0.0919286
R23887 VSS.n8628 VSS.n205 0.0919286
R23888 VSS.n213 VSS.n211 0.0919286
R23889 VSS.n8636 VSS.n8635 0.0919286
R23890 VSS.n1437 VSS.n1436 0.0919286
R23891 VSS.n1445 VSS.n1363 0.0919286
R23892 VSS.n1668 VSS.n1667 0.0919286
R23893 VSS.n1629 VSS.n1628 0.0919286
R23894 VSS.n1579 VSS.n1537 0.0919286
R23895 VSS.n1310 VSS.n1151 0.0919286
R23896 VSS.n1159 VSS.n1157 0.0919286
R23897 VSS.n1318 VSS.n1317 0.0919286
R23898 VSS.n2010 VSS.n2009 0.0919286
R23899 VSS.n2018 VSS.n1936 0.0919286
R23900 VSS.n2260 VSS.n2259 0.0919286
R23901 VSS.n2221 VSS.n2220 0.0919286
R23902 VSS.n2139 VSS.n2110 0.0919286
R23903 VSS.n1883 VSS.n1724 0.0919286
R23904 VSS.n1732 VSS.n1730 0.0919286
R23905 VSS.n1891 VSS.n1890 0.0919286
R23906 VSS.n3767 VSS.n3766 0.0919286
R23907 VSS.n3781 VSS.n3443 0.0919286
R23908 VSS.n3811 VSS.n3810 0.0919286
R23909 VSS.n3850 VSS.n3415 0.0919286
R23910 VSS.n3901 VSS.n3900 0.0919286
R23911 VSS.n3677 VSS.n3518 0.0919286
R23912 VSS.n3526 VSS.n3524 0.0919286
R23913 VSS.n3685 VSS.n3684 0.0919286
R23914 VSS.n4359 VSS.n4358 0.0919286
R23915 VSS.n4373 VSS.n4035 0.0919286
R23916 VSS.n4403 VSS.n4402 0.0919286
R23917 VSS.n4442 VSS.n4007 0.0919286
R23918 VSS.n4493 VSS.n4492 0.0919286
R23919 VSS.n4269 VSS.n4110 0.0919286
R23920 VSS.n4118 VSS.n4116 0.0919286
R23921 VSS.n4277 VSS.n4276 0.0919286
R23922 VSS.n4951 VSS.n4950 0.0919286
R23923 VSS.n4965 VSS.n4627 0.0919286
R23924 VSS.n4995 VSS.n4994 0.0919286
R23925 VSS.n5034 VSS.n4599 0.0919286
R23926 VSS.n5085 VSS.n5084 0.0919286
R23927 VSS.n4861 VSS.n4702 0.0919286
R23928 VSS.n4710 VSS.n4708 0.0919286
R23929 VSS.n4869 VSS.n4868 0.0919286
R23930 VSS.n5543 VSS.n5542 0.0919286
R23931 VSS.n5557 VSS.n5219 0.0919286
R23932 VSS.n5587 VSS.n5586 0.0919286
R23933 VSS.n5626 VSS.n5191 0.0919286
R23934 VSS.n5677 VSS.n5676 0.0919286
R23935 VSS.n5453 VSS.n5294 0.0919286
R23936 VSS.n5302 VSS.n5300 0.0919286
R23937 VSS.n5461 VSS.n5460 0.0919286
R23938 VSS.n6135 VSS.n6134 0.0919286
R23939 VSS.n6149 VSS.n5811 0.0919286
R23940 VSS.n6179 VSS.n6178 0.0919286
R23941 VSS.n6218 VSS.n5783 0.0919286
R23942 VSS.n6269 VSS.n6268 0.0919286
R23943 VSS.n6045 VSS.n5886 0.0919286
R23944 VSS.n5894 VSS.n5892 0.0919286
R23945 VSS.n6053 VSS.n6052 0.0919286
R23946 VSS.n6727 VSS.n6726 0.0919286
R23947 VSS.n6741 VSS.n6403 0.0919286
R23948 VSS.n6771 VSS.n6770 0.0919286
R23949 VSS.n6810 VSS.n6375 0.0919286
R23950 VSS.n6861 VSS.n6860 0.0919286
R23951 VSS.n6637 VSS.n6478 0.0919286
R23952 VSS.n6486 VSS.n6484 0.0919286
R23953 VSS.n6645 VSS.n6644 0.0919286
R23954 VSS.n2608 VSS.n2607 0.0919286
R23955 VSS.n2616 VSS.n2534 0.0919286
R23956 VSS.n7004 VSS.n7003 0.0919286
R23957 VSS.n6965 VSS.n6964 0.0919286
R23958 VSS.n2737 VSS.n2708 0.0919286
R23959 VSS.n2481 VSS.n2322 0.0919286
R23960 VSS.n2330 VSS.n2328 0.0919286
R23961 VSS.n2489 VSS.n2488 0.0919286
R23962 VSS.n3175 VSS.n3174 0.0919286
R23963 VSS.n3189 VSS.n2850 0.0919286
R23964 VSS.n3219 VSS.n3218 0.0919286
R23965 VSS.n3258 VSS.n2822 0.0919286
R23966 VSS.n3309 VSS.n3308 0.0919286
R23967 VSS.n3071 VSS.n3070 0.0919286
R23968 VSS.n3085 VSS.n2925 0.0919286
R23969 VSS.n3093 VSS.n3092 0.0919286
R23970 VSS.n9135 VSS.n9134 0.0919286
R23971 VSS.n9149 VSS.n117 0.0919286
R23972 VSS.n9179 VSS.n9178 0.0919286
R23973 VSS.n9218 VSS.n89 0.0919286
R23974 VSS.n9269 VSS.n9268 0.0919286
R23975 VSS.n380 VSS.n312 0.0919286
R23976 VSS.n389 VSS.n388 0.0919286
R23977 VSS.n9053 VSS.n9052 0.0919286
R23978 VSS.n600 VSS.n599 0.0919286
R23979 VSS.n608 VSS.n523 0.0919286
R23980 VSS.n823 VSS.n822 0.0919286
R23981 VSS.n784 VSS.n783 0.0919286
R23982 VSS.n738 VSS.n700 0.0919286
R23983 VSS.n944 VSS.n943 0.0919286
R23984 VSS.n952 VSS.n870 0.0919286
R23985 VSS.n960 VSS.n959 0.0919286
R23986 VSS.n8393 VSS.n8392 0.0919286
R23987 VSS.n7305 VSS.n7276 0.0919286
R23988 VSS.n8516 VSS.n8515 0.024
R23989 VSS.n8486 VSS.n8485 0.024
R23990 VSS.n7500 VSS.n7499 0.024
R23991 VSS.n7571 VSS.n7570 0.024
R23992 VSS.n7994 VSS.n7993 0.024
R23993 VSS.n8056 VSS.n8055 0.024
R23994 VSS.n8092 VSS.n8091 0.024
R23995 VSS.n8163 VSS.n8162 0.024
R23996 VSS.n8555 VSS.n8554 0.024
R23997 VSS.n8617 VSS.n8616 0.024
R23998 VSS.n9040 VSS.n9039 0.024
R23999 VSS.n9010 VSS.n9009 0.024
R24000 VSS.n1237 VSS.n1236 0.024
R24001 VSS.n1299 VSS.n1298 0.024
R24002 VSS.n1703 VSS.n1702 0.024
R24003 VSS.n1673 VSS.n1672 0.024
R24004 VSS.n1810 VSS.n1809 0.024
R24005 VSS.n1872 VSS.n1871 0.024
R24006 VSS.n2295 VSS.n2294 0.024
R24007 VSS.n2265 VSS.n2264 0.024
R24008 VSS.n3604 VSS.n3603 0.024
R24009 VSS.n3666 VSS.n3665 0.024
R24010 VSS.n3702 VSS.n3701 0.024
R24011 VSS.n3773 VSS.n3772 0.024
R24012 VSS.n4196 VSS.n4195 0.024
R24013 VSS.n4258 VSS.n4257 0.024
R24014 VSS.n4294 VSS.n4293 0.024
R24015 VSS.n4365 VSS.n4364 0.024
R24016 VSS.n4788 VSS.n4787 0.024
R24017 VSS.n4850 VSS.n4849 0.024
R24018 VSS.n4886 VSS.n4885 0.024
R24019 VSS.n4957 VSS.n4956 0.024
R24020 VSS.n5380 VSS.n5379 0.024
R24021 VSS.n5442 VSS.n5441 0.024
R24022 VSS.n5478 VSS.n5477 0.024
R24023 VSS.n5549 VSS.n5548 0.024
R24024 VSS.n5972 VSS.n5971 0.024
R24025 VSS.n6034 VSS.n6033 0.024
R24026 VSS.n6070 VSS.n6069 0.024
R24027 VSS.n6141 VSS.n6140 0.024
R24028 VSS.n6564 VSS.n6563 0.024
R24029 VSS.n6626 VSS.n6625 0.024
R24030 VSS.n6662 VSS.n6661 0.024
R24031 VSS.n6733 VSS.n6732 0.024
R24032 VSS.n2408 VSS.n2407 0.024
R24033 VSS.n2470 VSS.n2469 0.024
R24034 VSS.n7039 VSS.n7038 0.024
R24035 VSS.n7009 VSS.n7008 0.024
R24036 VSS.n3005 VSS.n3004 0.024
R24037 VSS.n3077 VSS.n3076 0.024
R24038 VSS.n3110 VSS.n3109 0.024
R24039 VSS.n3181 VSS.n3180 0.024
R24040 VSS.n430 VSS.n429 0.024
R24041 VSS.n400 VSS.n399 0.024
R24042 VSS.n9070 VSS.n9069 0.024
R24043 VSS.n9141 VSS.n9140 0.024
R24044 VSS.n995 VSS.n994 0.024
R24045 VSS.n965 VSS.n964 0.024
R24046 VSS.n858 VSS.n857 0.024
R24047 VSS.n828 VSS.n827 0.024
R24048 VSS.n8467 VSS.n8466 0.024
R24049 VSS.n8437 VSS.n8436 0.024
R24050 VSS.n8456 VSS.n8455 0.0228214
R24051 VSS.n8448 VSS.n8447 0.0228214
R24052 VSS.n8440 VSS.n7089 0.0228214
R24053 VSS.n984 VSS.n983 0.0228214
R24054 VSS.n976 VSS.n975 0.0228214
R24055 VSS.n968 VSS.n471 0.0228214
R24056 VSS.n7459 VSS.n7448 0.0228214
R24057 VSS.n7544 VSS.n7543 0.0228214
R24058 VSS.n7552 VSS.n7426 0.0228214
R24059 VSS.n8505 VSS.n8504 0.0228214
R24060 VSS.n8497 VSS.n8496 0.0228214
R24061 VSS.n8489 VSS.n1038 0.0228214
R24062 VSS.n7683 VSS.n7369 0.0228214
R24063 VSS.n7873 VSS.n7862 0.0228214
R24064 VSS.n8136 VSS.n8135 0.0228214
R24065 VSS.n8144 VSS.n7840 0.0228214
R24066 VSS.n8022 VSS.n8021 0.0228214
R24067 VSS.n7943 VSS.n7925 0.0228214
R24068 VSS.n8052 VSS.n7920 0.0228214
R24069 VSS.n8275 VSS.n7783 0.0228214
R24070 VSS.n8583 VSS.n8582 0.0228214
R24071 VSS.n240 VSS.n222 0.0228214
R24072 VSS.n8613 VSS.n217 0.0228214
R24073 VSS.n9029 VSS.n9028 0.0228214
R24074 VSS.n9021 VSS.n9020 0.0228214
R24075 VSS.n9013 VSS.n8668 0.0228214
R24076 VSS.n8952 VSS.n8851 0.0228214
R24077 VSS.n1265 VSS.n1264 0.0228214
R24078 VSS.n1186 VSS.n1168 0.0228214
R24079 VSS.n1295 VSS.n1163 0.0228214
R24080 VSS.n1692 VSS.n1691 0.0228214
R24081 VSS.n1684 VSS.n1683 0.0228214
R24082 VSS.n1676 VSS.n1350 0.0228214
R24083 VSS.n1613 VSS.n1612 0.0228214
R24084 VSS.n1838 VSS.n1837 0.0228214
R24085 VSS.n1759 VSS.n1741 0.0228214
R24086 VSS.n1868 VSS.n1736 0.0228214
R24087 VSS.n2284 VSS.n2283 0.0228214
R24088 VSS.n2276 VSS.n2275 0.0228214
R24089 VSS.n2268 VSS.n1923 0.0228214
R24090 VSS.n2205 VSS.n2204 0.0228214
R24091 VSS.n3632 VSS.n3631 0.0228214
R24092 VSS.n3553 VSS.n3535 0.0228214
R24093 VSS.n3662 VSS.n3530 0.0228214
R24094 VSS.n3483 VSS.n3472 0.0228214
R24095 VSS.n3746 VSS.n3745 0.0228214
R24096 VSS.n3754 VSS.n3450 0.0228214
R24097 VSS.n3885 VSS.n3393 0.0228214
R24098 VSS.n4224 VSS.n4223 0.0228214
R24099 VSS.n4145 VSS.n4127 0.0228214
R24100 VSS.n4254 VSS.n4122 0.0228214
R24101 VSS.n4075 VSS.n4064 0.0228214
R24102 VSS.n4338 VSS.n4337 0.0228214
R24103 VSS.n4346 VSS.n4042 0.0228214
R24104 VSS.n4477 VSS.n3985 0.0228214
R24105 VSS.n4816 VSS.n4815 0.0228214
R24106 VSS.n4737 VSS.n4719 0.0228214
R24107 VSS.n4846 VSS.n4714 0.0228214
R24108 VSS.n4667 VSS.n4656 0.0228214
R24109 VSS.n4930 VSS.n4929 0.0228214
R24110 VSS.n4938 VSS.n4634 0.0228214
R24111 VSS.n5069 VSS.n4577 0.0228214
R24112 VSS.n5408 VSS.n5407 0.0228214
R24113 VSS.n5329 VSS.n5311 0.0228214
R24114 VSS.n5438 VSS.n5306 0.0228214
R24115 VSS.n5259 VSS.n5248 0.0228214
R24116 VSS.n5522 VSS.n5521 0.0228214
R24117 VSS.n5530 VSS.n5226 0.0228214
R24118 VSS.n5661 VSS.n5169 0.0228214
R24119 VSS.n6000 VSS.n5999 0.0228214
R24120 VSS.n5921 VSS.n5903 0.0228214
R24121 VSS.n6030 VSS.n5898 0.0228214
R24122 VSS.n5851 VSS.n5840 0.0228214
R24123 VSS.n6114 VSS.n6113 0.0228214
R24124 VSS.n6122 VSS.n5818 0.0228214
R24125 VSS.n6253 VSS.n5761 0.0228214
R24126 VSS.n6592 VSS.n6591 0.0228214
R24127 VSS.n6513 VSS.n6495 0.0228214
R24128 VSS.n6622 VSS.n6490 0.0228214
R24129 VSS.n6443 VSS.n6432 0.0228214
R24130 VSS.n6706 VSS.n6705 0.0228214
R24131 VSS.n6714 VSS.n6410 0.0228214
R24132 VSS.n6845 VSS.n6353 0.0228214
R24133 VSS.n2436 VSS.n2435 0.0228214
R24134 VSS.n2357 VSS.n2339 0.0228214
R24135 VSS.n2466 VSS.n2334 0.0228214
R24136 VSS.n7028 VSS.n7027 0.0228214
R24137 VSS.n7020 VSS.n7019 0.0228214
R24138 VSS.n7012 VSS.n2521 0.0228214
R24139 VSS.n6949 VSS.n6948 0.0228214
R24140 VSS.n2967 VSS.n2954 0.0228214
R24141 VSS.n3049 VSS.n3048 0.0228214
R24142 VSS.n3057 VSS.n2932 0.0228214
R24143 VSS.n2890 VSS.n2879 0.0228214
R24144 VSS.n3154 VSS.n3153 0.0228214
R24145 VSS.n3162 VSS.n2857 0.0228214
R24146 VSS.n3293 VSS.n2800 0.0228214
R24147 VSS.n419 VSS.n418 0.0228214
R24148 VSS.n411 VSS.n410 0.0228214
R24149 VSS.n403 VSS.n305 0.0228214
R24150 VSS.n157 VSS.n146 0.0228214
R24151 VSS.n9114 VSS.n9113 0.0228214
R24152 VSS.n9122 VSS.n124 0.0228214
R24153 VSS.n9253 VSS.n67 0.0228214
R24154 VSS.n847 VSS.n846 0.0228214
R24155 VSS.n839 VSS.n838 0.0228214
R24156 VSS.n831 VSS.n510 0.0228214
R24157 VSS.n768 VSS.n767 0.0228214
R24158 VSS.n8377 VSS.n8376 0.0228214
R24159 VSS.n8463 VSS.n7067 0.0210357
R24160 VSS.n991 VSS.n448 0.0210357
R24161 VSS.n7472 VSS.n7464 0.0210357
R24162 VSS.n8512 VSS.n1015 0.0210357
R24163 VSS.n7650 VSS.n7390 0.0210357
R24164 VSS.n7690 VSS.n7376 0.0210357
R24165 VSS.n7689 VSS.n7378 0.0210357
R24166 VSS.n7886 VSS.n7878 0.0210357
R24167 VSS.n7966 VSS.n7965 0.0210357
R24168 VSS.n8242 VSS.n7804 0.0210357
R24169 VSS.n8282 VSS.n7790 0.0210357
R24170 VSS.n8281 VSS.n7792 0.0210357
R24171 VSS.n263 VSS.n262 0.0210357
R24172 VSS.n9036 VSS.n8646 0.0210357
R24173 VSS.n8971 VSS.n8970 0.0210357
R24174 VSS.n8864 VSS.n8819 0.0210357
R24175 VSS.n8863 VSS.n8817 0.0210357
R24176 VSS.n1209 VSS.n1208 0.0210357
R24177 VSS.n1699 VSS.n1328 0.0210357
R24178 VSS.n1631 VSS.n1500 0.0210357
R24179 VSS.n1620 VSS.n1507 0.0210357
R24180 VSS.n1619 VSS.n1509 0.0210357
R24181 VSS.n1782 VSS.n1781 0.0210357
R24182 VSS.n2291 VSS.n1901 0.0210357
R24183 VSS.n2223 VSS.n2073 0.0210357
R24184 VSS.n2212 VSS.n2080 0.0210357
R24185 VSS.n2211 VSS.n2082 0.0210357
R24186 VSS.n3576 VSS.n3575 0.0210357
R24187 VSS.n3496 VSS.n3488 0.0210357
R24188 VSS.n3852 VSS.n3414 0.0210357
R24189 VSS.n3892 VSS.n3400 0.0210357
R24190 VSS.n3891 VSS.n3402 0.0210357
R24191 VSS.n4168 VSS.n4167 0.0210357
R24192 VSS.n4088 VSS.n4080 0.0210357
R24193 VSS.n4444 VSS.n4006 0.0210357
R24194 VSS.n4484 VSS.n3992 0.0210357
R24195 VSS.n4483 VSS.n3994 0.0210357
R24196 VSS.n4760 VSS.n4759 0.0210357
R24197 VSS.n4680 VSS.n4672 0.0210357
R24198 VSS.n5036 VSS.n4598 0.0210357
R24199 VSS.n5076 VSS.n4584 0.0210357
R24200 VSS.n5075 VSS.n4586 0.0210357
R24201 VSS.n5352 VSS.n5351 0.0210357
R24202 VSS.n5272 VSS.n5264 0.0210357
R24203 VSS.n5628 VSS.n5190 0.0210357
R24204 VSS.n5668 VSS.n5176 0.0210357
R24205 VSS.n5667 VSS.n5178 0.0210357
R24206 VSS.n5944 VSS.n5943 0.0210357
R24207 VSS.n5864 VSS.n5856 0.0210357
R24208 VSS.n6220 VSS.n5782 0.0210357
R24209 VSS.n6260 VSS.n5768 0.0210357
R24210 VSS.n6259 VSS.n5770 0.0210357
R24211 VSS.n6536 VSS.n6535 0.0210357
R24212 VSS.n6456 VSS.n6448 0.0210357
R24213 VSS.n6812 VSS.n6374 0.0210357
R24214 VSS.n6852 VSS.n6360 0.0210357
R24215 VSS.n6851 VSS.n6362 0.0210357
R24216 VSS.n2380 VSS.n2379 0.0210357
R24217 VSS.n7035 VSS.n2499 0.0210357
R24218 VSS.n6967 VSS.n2671 0.0210357
R24219 VSS.n6956 VSS.n2678 0.0210357
R24220 VSS.n6955 VSS.n2680 0.0210357
R24221 VSS.n2978 VSS.n2971 0.0210357
R24222 VSS.n2903 VSS.n2895 0.0210357
R24223 VSS.n3260 VSS.n2821 0.0210357
R24224 VSS.n3300 VSS.n2807 0.0210357
R24225 VSS.n3299 VSS.n2809 0.0210357
R24226 VSS.n426 VSS.n282 0.0210357
R24227 VSS.n170 VSS.n162 0.0210357
R24228 VSS.n9220 VSS.n88 0.0210357
R24229 VSS.n9260 VSS.n74 0.0210357
R24230 VSS.n9259 VSS.n76 0.0210357
R24231 VSS.n854 VSS.n488 0.0210357
R24232 VSS.n786 VSS.n663 0.0210357
R24233 VSS.n775 VSS.n670 0.0210357
R24234 VSS.n774 VSS.n672 0.0210357
R24235 VSS.n8395 VSS.n7239 0.0210357
R24236 VSS.n8384 VSS.n7246 0.0210357
R24237 VSS.n8383 VSS.n7248 0.0210357
R24238 VSS.n7666 VSS.n7376 0.0201429
R24239 VSS.n7707 VSS.n7357 0.0201429
R24240 VSS.n7667 VSS.n7378 0.0201429
R24241 VSS.n8258 VSS.n7790 0.0201429
R24242 VSS.n8299 VSS.n7771 0.0201429
R24243 VSS.n8259 VSS.n7792 0.0201429
R24244 VSS.n8963 VSS.n8819 0.0201429
R24245 VSS.n8946 VSS.n8945 0.0201429
R24246 VSS.n8964 VSS.n8817 0.0201429
R24247 VSS.n1527 VSS.n1507 0.0201429
R24248 VSS.n1602 VSS.n1543 0.0201429
R24249 VSS.n1528 VSS.n1509 0.0201429
R24250 VSS.n2100 VSS.n2080 0.0201429
R24251 VSS.n2194 VSS.n2116 0.0201429
R24252 VSS.n2101 VSS.n2082 0.0201429
R24253 VSS.n3868 VSS.n3400 0.0201429
R24254 VSS.n3909 VSS.n3381 0.0201429
R24255 VSS.n3869 VSS.n3402 0.0201429
R24256 VSS.n4460 VSS.n3992 0.0201429
R24257 VSS.n4501 VSS.n3973 0.0201429
R24258 VSS.n4461 VSS.n3994 0.0201429
R24259 VSS.n5052 VSS.n4584 0.0201429
R24260 VSS.n5093 VSS.n4565 0.0201429
R24261 VSS.n5053 VSS.n4586 0.0201429
R24262 VSS.n5644 VSS.n5176 0.0201429
R24263 VSS.n5685 VSS.n5157 0.0201429
R24264 VSS.n5645 VSS.n5178 0.0201429
R24265 VSS.n6236 VSS.n5768 0.0201429
R24266 VSS.n6277 VSS.n5749 0.0201429
R24267 VSS.n6237 VSS.n5770 0.0201429
R24268 VSS.n6828 VSS.n6360 0.0201429
R24269 VSS.n6869 VSS.n6341 0.0201429
R24270 VSS.n6829 VSS.n6362 0.0201429
R24271 VSS.n2698 VSS.n2678 0.0201429
R24272 VSS.n6938 VSS.n2714 0.0201429
R24273 VSS.n2699 VSS.n2680 0.0201429
R24274 VSS.n3276 VSS.n2807 0.0201429
R24275 VSS.n3317 VSS.n2788 0.0201429
R24276 VSS.n3277 VSS.n2809 0.0201429
R24277 VSS.n9236 VSS.n74 0.0201429
R24278 VSS.n9277 VSS.n55 0.0201429
R24279 VSS.n9237 VSS.n76 0.0201429
R24280 VSS.n690 VSS.n670 0.0201429
R24281 VSS.n757 VSS.n706 0.0201429
R24282 VSS.n691 VSS.n672 0.0201429
R24283 VSS.n7266 VSS.n7246 0.0201429
R24284 VSS.n8366 VSS.n7282 0.0201429
R24285 VSS.n7267 VSS.n7248 0.0201429
R24286 VSS.n7633 VSS.n7632 0.01925
R24287 VSS.n8225 VSS.n8224 0.01925
R24288 VSS.n8981 VSS.n8802 0.01925
R24289 VSS.n1495 VSS.n1482 0.01925
R24290 VSS.n2068 VSS.n2055 0.01925
R24291 VSS.n3835 VSS.n3834 0.01925
R24292 VSS.n4427 VSS.n4426 0.01925
R24293 VSS.n5019 VSS.n5018 0.01925
R24294 VSS.n5611 VSS.n5610 0.01925
R24295 VSS.n6203 VSS.n6202 0.01925
R24296 VSS.n6795 VSS.n6794 0.01925
R24297 VSS.n2666 VSS.n2653 0.01925
R24298 VSS.n3243 VSS.n3242 0.01925
R24299 VSS.n9203 VSS.n9202 0.01925
R24300 VSS.n658 VSS.n645 0.01925
R24301 VSS.n7234 VSS.n7221 0.01925
R24302 VSS.n7080 VSS.n7073 0.0174643
R24303 VSS.n8449 VSS.n7080 0.0174643
R24304 VSS.n8453 VSS.n7076 0.0174643
R24305 VSS.n8450 VSS.n7076 0.0174643
R24306 VSS.n977 VSS.n462 0.0174643
R24307 VSS.n7536 VSS.n7535 0.0174643
R24308 VSS.n7535 VSS.n7442 0.0174643
R24309 VSS.n8498 VSS.n1029 0.0174643
R24310 VSS.n8499 VSS.n1027 0.0174643
R24311 VSS.n7658 VSS.n7381 0.0174643
R24312 VSS.n7537 VSS.n7447 0.0174643
R24313 VSS.n7447 VSS.n7443 0.0174643
R24314 VSS.n8128 VSS.n8127 0.0174643
R24315 VSS.n8127 VSS.n7856 0.0174643
R24316 VSS.n8032 VSS.n7942 0.0174643
R24317 VSS.n8031 VSS.n8030 0.0174643
R24318 VSS.n8250 VSS.n7795 0.0174643
R24319 VSS.n8129 VSS.n7861 0.0174643
R24320 VSS.n7861 VSS.n7857 0.0174643
R24321 VSS.n8593 VSS.n239 0.0174643
R24322 VSS.n8659 VSS.n8652 0.0174643
R24323 VSS.n9022 VSS.n8659 0.0174643
R24324 VSS.n9026 VSS.n8655 0.0174643
R24325 VSS.n9023 VSS.n8655 0.0174643
R24326 VSS.n8816 VSS.n8810 0.0174643
R24327 VSS.n8592 VSS.n8591 0.0174643
R24328 VSS.n1275 VSS.n1185 0.0174643
R24329 VSS.n1341 VSS.n1334 0.0174643
R24330 VSS.n1685 VSS.n1341 0.0174643
R24331 VSS.n1689 VSS.n1337 0.0174643
R24332 VSS.n1686 VSS.n1337 0.0174643
R24333 VSS.n1519 VSS.n1512 0.0174643
R24334 VSS.n1274 VSS.n1273 0.0174643
R24335 VSS.n1848 VSS.n1758 0.0174643
R24336 VSS.n1914 VSS.n1907 0.0174643
R24337 VSS.n2277 VSS.n1914 0.0174643
R24338 VSS.n2281 VSS.n1910 0.0174643
R24339 VSS.n2278 VSS.n1910 0.0174643
R24340 VSS.n2092 VSS.n2085 0.0174643
R24341 VSS.n1847 VSS.n1846 0.0174643
R24342 VSS.n3642 VSS.n3552 0.0174643
R24343 VSS.n3738 VSS.n3737 0.0174643
R24344 VSS.n3737 VSS.n3466 0.0174643
R24345 VSS.n3739 VSS.n3471 0.0174643
R24346 VSS.n3471 VSS.n3467 0.0174643
R24347 VSS.n3860 VSS.n3405 0.0174643
R24348 VSS.n3641 VSS.n3640 0.0174643
R24349 VSS.n4234 VSS.n4144 0.0174643
R24350 VSS.n4330 VSS.n4329 0.0174643
R24351 VSS.n4329 VSS.n4058 0.0174643
R24352 VSS.n4331 VSS.n4063 0.0174643
R24353 VSS.n4063 VSS.n4059 0.0174643
R24354 VSS.n4452 VSS.n3997 0.0174643
R24355 VSS.n4233 VSS.n4232 0.0174643
R24356 VSS.n4826 VSS.n4736 0.0174643
R24357 VSS.n4922 VSS.n4921 0.0174643
R24358 VSS.n4921 VSS.n4650 0.0174643
R24359 VSS.n4923 VSS.n4655 0.0174643
R24360 VSS.n4655 VSS.n4651 0.0174643
R24361 VSS.n5044 VSS.n4589 0.0174643
R24362 VSS.n4825 VSS.n4824 0.0174643
R24363 VSS.n5418 VSS.n5328 0.0174643
R24364 VSS.n5514 VSS.n5513 0.0174643
R24365 VSS.n5513 VSS.n5242 0.0174643
R24366 VSS.n5515 VSS.n5247 0.0174643
R24367 VSS.n5247 VSS.n5243 0.0174643
R24368 VSS.n5636 VSS.n5181 0.0174643
R24369 VSS.n5417 VSS.n5416 0.0174643
R24370 VSS.n6010 VSS.n5920 0.0174643
R24371 VSS.n6106 VSS.n6105 0.0174643
R24372 VSS.n6105 VSS.n5834 0.0174643
R24373 VSS.n6107 VSS.n5839 0.0174643
R24374 VSS.n5839 VSS.n5835 0.0174643
R24375 VSS.n6228 VSS.n5773 0.0174643
R24376 VSS.n6009 VSS.n6008 0.0174643
R24377 VSS.n6602 VSS.n6512 0.0174643
R24378 VSS.n6698 VSS.n6697 0.0174643
R24379 VSS.n6697 VSS.n6426 0.0174643
R24380 VSS.n6699 VSS.n6431 0.0174643
R24381 VSS.n6431 VSS.n6427 0.0174643
R24382 VSS.n6820 VSS.n6365 0.0174643
R24383 VSS.n6601 VSS.n6600 0.0174643
R24384 VSS.n2446 VSS.n2356 0.0174643
R24385 VSS.n2512 VSS.n2505 0.0174643
R24386 VSS.n7021 VSS.n2512 0.0174643
R24387 VSS.n7025 VSS.n2508 0.0174643
R24388 VSS.n7022 VSS.n2508 0.0174643
R24389 VSS.n2690 VSS.n2683 0.0174643
R24390 VSS.n2445 VSS.n2444 0.0174643
R24391 VSS.n2956 VSS.n2948 0.0174643
R24392 VSS.n3146 VSS.n3145 0.0174643
R24393 VSS.n3145 VSS.n2873 0.0174643
R24394 VSS.n3147 VSS.n2878 0.0174643
R24395 VSS.n2878 VSS.n2874 0.0174643
R24396 VSS.n3268 VSS.n2812 0.0174643
R24397 VSS.n2955 VSS.n2949 0.0174643
R24398 VSS.n412 VSS.n296 0.0174643
R24399 VSS.n9106 VSS.n9105 0.0174643
R24400 VSS.n9105 VSS.n140 0.0174643
R24401 VSS.n9107 VSS.n145 0.0174643
R24402 VSS.n145 VSS.n141 0.0174643
R24403 VSS.n9228 VSS.n79 0.0174643
R24404 VSS.n413 VSS.n294 0.0174643
R24405 VSS.n501 VSS.n494 0.0174643
R24406 VSS.n840 VSS.n501 0.0174643
R24407 VSS.n844 VSS.n497 0.0174643
R24408 VSS.n841 VSS.n497 0.0174643
R24409 VSS.n682 VSS.n675 0.0174643
R24410 VSS.n978 VSS.n460 0.0174643
R24411 VSS.n7258 VSS.n7251 0.0174643
R24412 VSS.n7132 VSS.n7131 0.0165714
R24413 VSS.n8442 VSS.n8441 0.0165714
R24414 VSS.n7181 VSS.n7179 0.0165714
R24415 VSS.n879 VSS.n454 0.0165714
R24416 VSS.n1060 VSS.n1021 0.0165714
R24417 VSS.n1082 VSS.n1081 0.0165714
R24418 VSS.n8511 VSS.n8510 0.0165714
R24419 VSS.n8510 VSS.n1016 0.0165714
R24420 VSS.n8502 VSS.n1024 0.0165714
R24421 VSS.n1130 VSS.n1128 0.0165714
R24422 VSS.n7668 VSS.n7381 0.0165714
R24423 VSS.n7688 VSS.n7379 0.0165714
R24424 VSS.n7676 VSS.n7672 0.0165714
R24425 VSS.n7493 VSS.n7492 0.0165714
R24426 VSS.n7549 VSS.n7439 0.0165714
R24427 VSS.n7576 VSS.n7422 0.0165714
R24428 VSS.n8033 VSS.n7940 0.0165714
R24429 VSS.n7987 VSS.n7986 0.0165714
R24430 VSS.n8015 VSS.n7950 0.0165714
R24431 VSS.n8015 VSS.n8014 0.0165714
R24432 VSS.n8024 VSS.n7941 0.0165714
R24433 VSS.n8063 VSS.n8062 0.0165714
R24434 VSS.n8260 VSS.n7795 0.0165714
R24435 VSS.n8280 VSS.n7793 0.0165714
R24436 VSS.n8268 VSS.n8264 0.0165714
R24437 VSS.n8085 VSS.n8084 0.0165714
R24438 VSS.n8141 VSS.n7853 0.0165714
R24439 VSS.n8168 VSS.n7836 0.0165714
R24440 VSS.n8594 VSS.n237 0.0165714
R24441 VSS.n8711 VSS.n8710 0.0165714
R24442 VSS.n9015 VSS.n9014 0.0165714
R24443 VSS.n8760 VSS.n8758 0.0165714
R24444 VSS.n8965 VSS.n8816 0.0165714
R24445 VSS.n8862 VSS.n8860 0.0165714
R24446 VSS.n8858 VSS.n8856 0.0165714
R24447 VSS.n8548 VSS.n8547 0.0165714
R24448 VSS.n8576 VSS.n247 0.0165714
R24449 VSS.n8576 VSS.n8575 0.0165714
R24450 VSS.n8585 VSS.n238 0.0165714
R24451 VSS.n8624 VSS.n8623 0.0165714
R24452 VSS.n1276 VSS.n1183 0.0165714
R24453 VSS.n1393 VSS.n1392 0.0165714
R24454 VSS.n1678 VSS.n1677 0.0165714
R24455 VSS.n1442 VSS.n1440 0.0165714
R24456 VSS.n1529 VSS.n1512 0.0165714
R24457 VSS.n1618 VSS.n1510 0.0165714
R24458 VSS.n1575 VSS.n1533 0.0165714
R24459 VSS.n1230 VSS.n1229 0.0165714
R24460 VSS.n1258 VSS.n1193 0.0165714
R24461 VSS.n1258 VSS.n1257 0.0165714
R24462 VSS.n1267 VSS.n1184 0.0165714
R24463 VSS.n1306 VSS.n1305 0.0165714
R24464 VSS.n1849 VSS.n1756 0.0165714
R24465 VSS.n1966 VSS.n1965 0.0165714
R24466 VSS.n2270 VSS.n2269 0.0165714
R24467 VSS.n2015 VSS.n2013 0.0165714
R24468 VSS.n2102 VSS.n2085 0.0165714
R24469 VSS.n2210 VSS.n2083 0.0165714
R24470 VSS.n2135 VSS.n2106 0.0165714
R24471 VSS.n1803 VSS.n1802 0.0165714
R24472 VSS.n1831 VSS.n1766 0.0165714
R24473 VSS.n1831 VSS.n1830 0.0165714
R24474 VSS.n1840 VSS.n1757 0.0165714
R24475 VSS.n1879 VSS.n1878 0.0165714
R24476 VSS.n3643 VSS.n3550 0.0165714
R24477 VSS.n3695 VSS.n3694 0.0165714
R24478 VSS.n3751 VSS.n3463 0.0165714
R24479 VSS.n3778 VSS.n3446 0.0165714
R24480 VSS.n3870 VSS.n3405 0.0165714
R24481 VSS.n3890 VSS.n3403 0.0165714
R24482 VSS.n3878 VSS.n3874 0.0165714
R24483 VSS.n3597 VSS.n3596 0.0165714
R24484 VSS.n3625 VSS.n3560 0.0165714
R24485 VSS.n3625 VSS.n3624 0.0165714
R24486 VSS.n3634 VSS.n3551 0.0165714
R24487 VSS.n3673 VSS.n3672 0.0165714
R24488 VSS.n4235 VSS.n4142 0.0165714
R24489 VSS.n4287 VSS.n4286 0.0165714
R24490 VSS.n4343 VSS.n4055 0.0165714
R24491 VSS.n4370 VSS.n4038 0.0165714
R24492 VSS.n4462 VSS.n3997 0.0165714
R24493 VSS.n4482 VSS.n3995 0.0165714
R24494 VSS.n4470 VSS.n4466 0.0165714
R24495 VSS.n4189 VSS.n4188 0.0165714
R24496 VSS.n4217 VSS.n4152 0.0165714
R24497 VSS.n4217 VSS.n4216 0.0165714
R24498 VSS.n4226 VSS.n4143 0.0165714
R24499 VSS.n4265 VSS.n4264 0.0165714
R24500 VSS.n4827 VSS.n4734 0.0165714
R24501 VSS.n4879 VSS.n4878 0.0165714
R24502 VSS.n4935 VSS.n4647 0.0165714
R24503 VSS.n4962 VSS.n4630 0.0165714
R24504 VSS.n5054 VSS.n4589 0.0165714
R24505 VSS.n5074 VSS.n4587 0.0165714
R24506 VSS.n5062 VSS.n5058 0.0165714
R24507 VSS.n4781 VSS.n4780 0.0165714
R24508 VSS.n4809 VSS.n4744 0.0165714
R24509 VSS.n4809 VSS.n4808 0.0165714
R24510 VSS.n4818 VSS.n4735 0.0165714
R24511 VSS.n4857 VSS.n4856 0.0165714
R24512 VSS.n5419 VSS.n5326 0.0165714
R24513 VSS.n5471 VSS.n5470 0.0165714
R24514 VSS.n5527 VSS.n5239 0.0165714
R24515 VSS.n5554 VSS.n5222 0.0165714
R24516 VSS.n5646 VSS.n5181 0.0165714
R24517 VSS.n5666 VSS.n5179 0.0165714
R24518 VSS.n5654 VSS.n5650 0.0165714
R24519 VSS.n5373 VSS.n5372 0.0165714
R24520 VSS.n5401 VSS.n5336 0.0165714
R24521 VSS.n5401 VSS.n5400 0.0165714
R24522 VSS.n5410 VSS.n5327 0.0165714
R24523 VSS.n5449 VSS.n5448 0.0165714
R24524 VSS.n6011 VSS.n5918 0.0165714
R24525 VSS.n6063 VSS.n6062 0.0165714
R24526 VSS.n6119 VSS.n5831 0.0165714
R24527 VSS.n6146 VSS.n5814 0.0165714
R24528 VSS.n6238 VSS.n5773 0.0165714
R24529 VSS.n6258 VSS.n5771 0.0165714
R24530 VSS.n6246 VSS.n6242 0.0165714
R24531 VSS.n5965 VSS.n5964 0.0165714
R24532 VSS.n5993 VSS.n5928 0.0165714
R24533 VSS.n5993 VSS.n5992 0.0165714
R24534 VSS.n6002 VSS.n5919 0.0165714
R24535 VSS.n6041 VSS.n6040 0.0165714
R24536 VSS.n6603 VSS.n6510 0.0165714
R24537 VSS.n6655 VSS.n6654 0.0165714
R24538 VSS.n6711 VSS.n6423 0.0165714
R24539 VSS.n6738 VSS.n6406 0.0165714
R24540 VSS.n6830 VSS.n6365 0.0165714
R24541 VSS.n6850 VSS.n6363 0.0165714
R24542 VSS.n6838 VSS.n6834 0.0165714
R24543 VSS.n6557 VSS.n6556 0.0165714
R24544 VSS.n6585 VSS.n6520 0.0165714
R24545 VSS.n6585 VSS.n6584 0.0165714
R24546 VSS.n6594 VSS.n6511 0.0165714
R24547 VSS.n6633 VSS.n6632 0.0165714
R24548 VSS.n2447 VSS.n2354 0.0165714
R24549 VSS.n2564 VSS.n2563 0.0165714
R24550 VSS.n7014 VSS.n7013 0.0165714
R24551 VSS.n2613 VSS.n2611 0.0165714
R24552 VSS.n2700 VSS.n2683 0.0165714
R24553 VSS.n6954 VSS.n2681 0.0165714
R24554 VSS.n2733 VSS.n2704 0.0165714
R24555 VSS.n2401 VSS.n2400 0.0165714
R24556 VSS.n2429 VSS.n2364 0.0165714
R24557 VSS.n2429 VSS.n2428 0.0165714
R24558 VSS.n2438 VSS.n2355 0.0165714
R24559 VSS.n2477 VSS.n2476 0.0165714
R24560 VSS.n3041 VSS.n3040 0.0165714
R24561 VSS.n3103 VSS.n3102 0.0165714
R24562 VSS.n3159 VSS.n2870 0.0165714
R24563 VSS.n3186 VSS.n2853 0.0165714
R24564 VSS.n3278 VSS.n2812 0.0165714
R24565 VSS.n3298 VSS.n2810 0.0165714
R24566 VSS.n3286 VSS.n3282 0.0165714
R24567 VSS.n2998 VSS.n2997 0.0165714
R24568 VSS.n3021 VSS.n2970 0.0165714
R24569 VSS.n3021 VSS.n3020 0.0165714
R24570 VSS.n3042 VSS.n2953 0.0165714
R24571 VSS.n3082 VSS.n2928 0.0165714
R24572 VSS.n362 VSS.n288 0.0165714
R24573 VSS.n9063 VSS.n9062 0.0165714
R24574 VSS.n9119 VSS.n137 0.0165714
R24575 VSS.n9146 VSS.n120 0.0165714
R24576 VSS.n9238 VSS.n79 0.0165714
R24577 VSS.n9258 VSS.n77 0.0165714
R24578 VSS.n9246 VSS.n9242 0.0165714
R24579 VSS.n337 VSS.n335 0.0165714
R24580 VSS.n425 VSS.n424 0.0165714
R24581 VSS.n424 VSS.n283 0.0165714
R24582 VSS.n416 VSS.n291 0.0165714
R24583 VSS.n393 VSS.n392 0.0165714
R24584 VSS.n556 VSS.n555 0.0165714
R24585 VSS.n833 VSS.n832 0.0165714
R24586 VSS.n605 VSS.n603 0.0165714
R24587 VSS.n692 VSS.n675 0.0165714
R24588 VSS.n773 VSS.n673 0.0165714
R24589 VSS.n734 VSS.n696 0.0165714
R24590 VSS.n901 VSS.n900 0.0165714
R24591 VSS.n990 VSS.n989 0.0165714
R24592 VSS.n989 VSS.n449 0.0165714
R24593 VSS.n981 VSS.n457 0.0165714
R24594 VSS.n949 VSS.n947 0.0165714
R24595 VSS.n7268 VSS.n7251 0.0165714
R24596 VSS.n8382 VSS.n7249 0.0165714
R24597 VSS.n7301 VSS.n7272 0.0165714
R24598 VSS.n8462 VSS.n8461 0.0156786
R24599 VSS.n8491 VSS.n8490 0.0156786
R24600 VSS.n7621 VSS.n7617 0.0156786
R24601 VSS.n7626 VSS.n7405 0.0156786
R24602 VSS.n7405 VSS.n7399 0.0156786
R24603 VSS.n7708 VSS.n7355 0.0156786
R24604 VSS.n7723 VSS.n7355 0.0156786
R24605 VSS.n7516 VSS.n7462 0.0156786
R24606 VSS.n8051 VSS.n8050 0.0156786
R24607 VSS.n8213 VSS.n8209 0.0156786
R24608 VSS.n8218 VSS.n7819 0.0156786
R24609 VSS.n7819 VSS.n7813 0.0156786
R24610 VSS.n8300 VSS.n7769 0.0156786
R24611 VSS.n8315 VSS.n7769 0.0156786
R24612 VSS.n8108 VSS.n7876 0.0156786
R24613 VSS.n9035 VSS.n9034 0.0156786
R24614 VSS.n8797 VSS.n8795 0.0156786
R24615 VSS.n8986 VSS.n8780 0.0156786
R24616 VSS.n8982 VSS.n8780 0.0156786
R24617 VSS.n8947 VSS.n8880 0.0156786
R24618 VSS.n8887 VSS.n8880 0.0156786
R24619 VSS.n8612 VSS.n8611 0.0156786
R24620 VSS.n1698 VSS.n1697 0.0156786
R24621 VSS.n1478 VSS.n1476 0.0156786
R24622 VSS.n1649 VSS.n1462 0.0156786
R24623 VSS.n1496 VSS.n1462 0.0156786
R24624 VSS.n1601 VSS.n1544 0.0156786
R24625 VSS.n1597 VSS.n1544 0.0156786
R24626 VSS.n1294 VSS.n1293 0.0156786
R24627 VSS.n2290 VSS.n2289 0.0156786
R24628 VSS.n2051 VSS.n2049 0.0156786
R24629 VSS.n2241 VSS.n2035 0.0156786
R24630 VSS.n2069 VSS.n2035 0.0156786
R24631 VSS.n2193 VSS.n2117 0.0156786
R24632 VSS.n2189 VSS.n2117 0.0156786
R24633 VSS.n1867 VSS.n1866 0.0156786
R24634 VSS.n3718 VSS.n3486 0.0156786
R24635 VSS.n3823 VSS.n3819 0.0156786
R24636 VSS.n3828 VSS.n3429 0.0156786
R24637 VSS.n3429 VSS.n3423 0.0156786
R24638 VSS.n3910 VSS.n3380 0.0156786
R24639 VSS.n3925 VSS.n3380 0.0156786
R24640 VSS.n3661 VSS.n3660 0.0156786
R24641 VSS.n4310 VSS.n4078 0.0156786
R24642 VSS.n4415 VSS.n4411 0.0156786
R24643 VSS.n4420 VSS.n4021 0.0156786
R24644 VSS.n4021 VSS.n4015 0.0156786
R24645 VSS.n4502 VSS.n3972 0.0156786
R24646 VSS.n4517 VSS.n3972 0.0156786
R24647 VSS.n4253 VSS.n4252 0.0156786
R24648 VSS.n4902 VSS.n4670 0.0156786
R24649 VSS.n5007 VSS.n5003 0.0156786
R24650 VSS.n5012 VSS.n4613 0.0156786
R24651 VSS.n4613 VSS.n4607 0.0156786
R24652 VSS.n5094 VSS.n4564 0.0156786
R24653 VSS.n5109 VSS.n4564 0.0156786
R24654 VSS.n4845 VSS.n4844 0.0156786
R24655 VSS.n5494 VSS.n5262 0.0156786
R24656 VSS.n5599 VSS.n5595 0.0156786
R24657 VSS.n5604 VSS.n5205 0.0156786
R24658 VSS.n5205 VSS.n5199 0.0156786
R24659 VSS.n5686 VSS.n5156 0.0156786
R24660 VSS.n5701 VSS.n5156 0.0156786
R24661 VSS.n5437 VSS.n5436 0.0156786
R24662 VSS.n6086 VSS.n5854 0.0156786
R24663 VSS.n6191 VSS.n6187 0.0156786
R24664 VSS.n6196 VSS.n5797 0.0156786
R24665 VSS.n5797 VSS.n5791 0.0156786
R24666 VSS.n6278 VSS.n5748 0.0156786
R24667 VSS.n6293 VSS.n5748 0.0156786
R24668 VSS.n6029 VSS.n6028 0.0156786
R24669 VSS.n6678 VSS.n6446 0.0156786
R24670 VSS.n6783 VSS.n6779 0.0156786
R24671 VSS.n6788 VSS.n6389 0.0156786
R24672 VSS.n6389 VSS.n6383 0.0156786
R24673 VSS.n6870 VSS.n6340 0.0156786
R24674 VSS.n6885 VSS.n6340 0.0156786
R24675 VSS.n6621 VSS.n6620 0.0156786
R24676 VSS.n7034 VSS.n7033 0.0156786
R24677 VSS.n2649 VSS.n2647 0.0156786
R24678 VSS.n6985 VSS.n2633 0.0156786
R24679 VSS.n2667 VSS.n2633 0.0156786
R24680 VSS.n6937 VSS.n2715 0.0156786
R24681 VSS.n6933 VSS.n2715 0.0156786
R24682 VSS.n2465 VSS.n2464 0.0156786
R24683 VSS.n3126 VSS.n2893 0.0156786
R24684 VSS.n3231 VSS.n3227 0.0156786
R24685 VSS.n3236 VSS.n2836 0.0156786
R24686 VSS.n2836 VSS.n2830 0.0156786
R24687 VSS.n3318 VSS.n2787 0.0156786
R24688 VSS.n3333 VSS.n2787 0.0156786
R24689 VSS.n3054 VSS.n2945 0.0156786
R24690 VSS.n9086 VSS.n160 0.0156786
R24691 VSS.n9191 VSS.n9187 0.0156786
R24692 VSS.n9196 VSS.n103 0.0156786
R24693 VSS.n103 VSS.n97 0.0156786
R24694 VSS.n9278 VSS.n54 0.0156786
R24695 VSS.n9293 VSS.n54 0.0156786
R24696 VSS.n405 VSS.n404 0.0156786
R24697 VSS.n853 VSS.n852 0.0156786
R24698 VSS.n641 VSS.n639 0.0156786
R24699 VSS.n804 VSS.n625 0.0156786
R24700 VSS.n659 VSS.n625 0.0156786
R24701 VSS.n756 VSS.n707 0.0156786
R24702 VSS.n752 VSS.n707 0.0156786
R24703 VSS.n970 VSS.n969 0.0156786
R24704 VSS.n7217 VSS.n7215 0.0156786
R24705 VSS.n8413 VSS.n7201 0.0156786
R24706 VSS.n7235 VSS.n7201 0.0156786
R24707 VSS.n8365 VSS.n7283 0.0156786
R24708 VSS.n8361 VSS.n7283 0.0156786
R24709 VSS.n8509 VSS.n8508 0.0152714
R24710 VSS.n8493 VSS.n8492 0.0152714
R24711 VSS.n7521 VSS.n7517 0.0152714
R24712 VSS.n7548 VSS.n7547 0.0152714
R24713 VSS.n7669 VSS.n7380 0.0152714
R24714 VSS.n7687 VSS.n7686 0.0152714
R24715 VSS.n8017 VSS.n8016 0.0152714
R24716 VSS.n8049 VSS.n8048 0.0152714
R24717 VSS.n8113 VSS.n8109 0.0152714
R24718 VSS.n8140 VSS.n8139 0.0152714
R24719 VSS.n8261 VSS.n7794 0.0152714
R24720 VSS.n8279 VSS.n8278 0.0152714
R24721 VSS.n8578 VSS.n8577 0.0152714
R24722 VSS.n8610 VSS.n8609 0.0152714
R24723 VSS.n9033 VSS.n9032 0.0152714
R24724 VSS.n9017 VSS.n9016 0.0152714
R24725 VSS.n8967 VSS.n8966 0.0152714
R24726 VSS.n8861 VSS.n8855 0.0152714
R24727 VSS.n1260 VSS.n1259 0.0152714
R24728 VSS.n1292 VSS.n1291 0.0152714
R24729 VSS.n1696 VSS.n1695 0.0152714
R24730 VSS.n1680 VSS.n1679 0.0152714
R24731 VSS.n1530 VSS.n1511 0.0152714
R24732 VSS.n1617 VSS.n1616 0.0152714
R24733 VSS.n1833 VSS.n1832 0.0152714
R24734 VSS.n1865 VSS.n1864 0.0152714
R24735 VSS.n2288 VSS.n2287 0.0152714
R24736 VSS.n2272 VSS.n2271 0.0152714
R24737 VSS.n2103 VSS.n2084 0.0152714
R24738 VSS.n2209 VSS.n2208 0.0152714
R24739 VSS.n3627 VSS.n3626 0.0152714
R24740 VSS.n3659 VSS.n3658 0.0152714
R24741 VSS.n3723 VSS.n3719 0.0152714
R24742 VSS.n3750 VSS.n3749 0.0152714
R24743 VSS.n3871 VSS.n3404 0.0152714
R24744 VSS.n3889 VSS.n3888 0.0152714
R24745 VSS.n4219 VSS.n4218 0.0152714
R24746 VSS.n4251 VSS.n4250 0.0152714
R24747 VSS.n4315 VSS.n4311 0.0152714
R24748 VSS.n4342 VSS.n4341 0.0152714
R24749 VSS.n4463 VSS.n3996 0.0152714
R24750 VSS.n4481 VSS.n4480 0.0152714
R24751 VSS.n4811 VSS.n4810 0.0152714
R24752 VSS.n4843 VSS.n4842 0.0152714
R24753 VSS.n4907 VSS.n4903 0.0152714
R24754 VSS.n4934 VSS.n4933 0.0152714
R24755 VSS.n5055 VSS.n4588 0.0152714
R24756 VSS.n5073 VSS.n5072 0.0152714
R24757 VSS.n5403 VSS.n5402 0.0152714
R24758 VSS.n5435 VSS.n5434 0.0152714
R24759 VSS.n5499 VSS.n5495 0.0152714
R24760 VSS.n5526 VSS.n5525 0.0152714
R24761 VSS.n5647 VSS.n5180 0.0152714
R24762 VSS.n5665 VSS.n5664 0.0152714
R24763 VSS.n5995 VSS.n5994 0.0152714
R24764 VSS.n6027 VSS.n6026 0.0152714
R24765 VSS.n6091 VSS.n6087 0.0152714
R24766 VSS.n6118 VSS.n6117 0.0152714
R24767 VSS.n6239 VSS.n5772 0.0152714
R24768 VSS.n6257 VSS.n6256 0.0152714
R24769 VSS.n6587 VSS.n6586 0.0152714
R24770 VSS.n6619 VSS.n6618 0.0152714
R24771 VSS.n6683 VSS.n6679 0.0152714
R24772 VSS.n6710 VSS.n6709 0.0152714
R24773 VSS.n6831 VSS.n6364 0.0152714
R24774 VSS.n6849 VSS.n6848 0.0152714
R24775 VSS.n2431 VSS.n2430 0.0152714
R24776 VSS.n2463 VSS.n2462 0.0152714
R24777 VSS.n7032 VSS.n7031 0.0152714
R24778 VSS.n7016 VSS.n7015 0.0152714
R24779 VSS.n2701 VSS.n2682 0.0152714
R24780 VSS.n6953 VSS.n6952 0.0152714
R24781 VSS.n3026 VSS.n3022 0.0152714
R24782 VSS.n3053 VSS.n3052 0.0152714
R24783 VSS.n3131 VSS.n3127 0.0152714
R24784 VSS.n3158 VSS.n3157 0.0152714
R24785 VSS.n3279 VSS.n2811 0.0152714
R24786 VSS.n3297 VSS.n3296 0.0152714
R24787 VSS.n423 VSS.n422 0.0152714
R24788 VSS.n407 VSS.n406 0.0152714
R24789 VSS.n9091 VSS.n9087 0.0152714
R24790 VSS.n9118 VSS.n9117 0.0152714
R24791 VSS.n9239 VSS.n78 0.0152714
R24792 VSS.n9257 VSS.n9256 0.0152714
R24793 VSS.n988 VSS.n987 0.0152714
R24794 VSS.n972 VSS.n971 0.0152714
R24795 VSS.n851 VSS.n850 0.0152714
R24796 VSS.n835 VSS.n834 0.0152714
R24797 VSS.n693 VSS.n674 0.0152714
R24798 VSS.n772 VSS.n771 0.0152714
R24799 VSS.n8460 VSS.n8459 0.0152714
R24800 VSS.n8444 VSS.n8443 0.0152714
R24801 VSS.n7269 VSS.n7250 0.0152714
R24802 VSS.n8381 VSS.n8380 0.0152714
R24803 VSS.n7656 VSS.n7385 0.0147857
R24804 VSS.n7673 VSS.n7367 0.0147857
R24805 VSS.n8248 VSS.n7799 0.0147857
R24806 VSS.n8265 VSS.n7781 0.0147857
R24807 VSS.n8812 VSS.n8809 0.0147857
R24808 VSS.n8875 VSS.n8853 0.0147857
R24809 VSS.n1517 VSS.n1491 0.0147857
R24810 VSS.n1546 VSS.n1545 0.0147857
R24811 VSS.n2090 VSS.n2064 0.0147857
R24812 VSS.n2119 VSS.n2118 0.0147857
R24813 VSS.n3858 VSS.n3409 0.0147857
R24814 VSS.n3875 VSS.n3391 0.0147857
R24815 VSS.n4450 VSS.n4001 0.0147857
R24816 VSS.n4467 VSS.n3983 0.0147857
R24817 VSS.n5042 VSS.n4593 0.0147857
R24818 VSS.n5059 VSS.n4575 0.0147857
R24819 VSS.n5634 VSS.n5185 0.0147857
R24820 VSS.n5651 VSS.n5167 0.0147857
R24821 VSS.n6226 VSS.n5777 0.0147857
R24822 VSS.n6243 VSS.n5759 0.0147857
R24823 VSS.n6818 VSS.n6369 0.0147857
R24824 VSS.n6835 VSS.n6351 0.0147857
R24825 VSS.n2688 VSS.n2662 0.0147857
R24826 VSS.n2717 VSS.n2716 0.0147857
R24827 VSS.n3266 VSS.n2816 0.0147857
R24828 VSS.n3283 VSS.n2798 0.0147857
R24829 VSS.n9226 VSS.n83 0.0147857
R24830 VSS.n9243 VSS.n65 0.0147857
R24831 VSS.n680 VSS.n654 0.0147857
R24832 VSS.n709 VSS.n708 0.0147857
R24833 VSS.n7256 VSS.n7230 0.0147857
R24834 VSS.n7285 VSS.n7284 0.0147857
R24835 VSS.n7729 VSS.n7728 0.0138929
R24836 VSS.n8321 VSS.n8320 0.0138929
R24837 VSS.n8896 VSS.n8889 0.0138929
R24838 VSS.n1558 VSS.n1557 0.0138929
R24839 VSS.n2166 VSS.n2153 0.0138929
R24840 VSS.n3932 VSS.n3931 0.0138929
R24841 VSS.n4524 VSS.n4523 0.0138929
R24842 VSS.n5116 VSS.n5115 0.0138929
R24843 VSS.n5708 VSS.n5707 0.0138929
R24844 VSS.n6300 VSS.n6299 0.0138929
R24845 VSS.n6892 VSS.n6891 0.0138929
R24846 VSS.n2764 VSS.n2751 0.0138929
R24847 VSS.n3340 VSS.n3339 0.0138929
R24848 VSS.n9300 VSS.n9299 0.0138929
R24849 VSS.n720 VSS.n33 0.0138929
R24850 VSS.n7332 VSS.n7319 0.0138929
R24851 VSS.n8501 VSS.n8500 0.0132571
R24852 VSS.n7539 VSS.n7538 0.0132571
R24853 VSS.n7625 VSS.n7623 0.0132571
R24854 VSS.n7653 VSS.n7386 0.0132571
R24855 VSS.n7706 VSS.n7705 0.0132571
R24856 VSS.n7726 VSS.n7724 0.0132571
R24857 VSS.n8029 VSS.n8025 0.0132571
R24858 VSS.n8131 VSS.n8130 0.0132571
R24859 VSS.n8217 VSS.n8215 0.0132571
R24860 VSS.n8245 VSS.n7800 0.0132571
R24861 VSS.n8298 VSS.n8297 0.0132571
R24862 VSS.n8318 VSS.n8316 0.0132571
R24863 VSS.n8590 VSS.n8586 0.0132571
R24864 VSS.n9025 VSS.n9024 0.0132571
R24865 VSS.n8985 VSS.n8799 0.0132571
R24866 VSS.n8983 VSS.n8800 0.0132571
R24867 VSS.n8949 VSS.n8948 0.0132571
R24868 VSS.n8933 VSS.n8891 0.0132571
R24869 VSS.n1272 VSS.n1268 0.0132571
R24870 VSS.n1688 VSS.n1687 0.0132571
R24871 VSS.n1481 VSS.n1480 0.0132571
R24872 VSS.n1498 VSS.n1497 0.0132571
R24873 VSS.n1600 VSS.n1548 0.0132571
R24874 VSS.n1598 VSS.n1549 0.0132571
R24875 VSS.n1845 VSS.n1841 0.0132571
R24876 VSS.n2280 VSS.n2279 0.0132571
R24877 VSS.n2054 VSS.n2053 0.0132571
R24878 VSS.n2071 VSS.n2070 0.0132571
R24879 VSS.n2192 VSS.n2121 0.0132571
R24880 VSS.n2190 VSS.n2122 0.0132571
R24881 VSS.n3639 VSS.n3635 0.0132571
R24882 VSS.n3741 VSS.n3740 0.0132571
R24883 VSS.n3827 VSS.n3825 0.0132571
R24884 VSS.n3855 VSS.n3410 0.0132571
R24885 VSS.n3908 VSS.n3907 0.0132571
R24886 VSS.n3927 VSS.n3926 0.0132571
R24887 VSS.n4231 VSS.n4227 0.0132571
R24888 VSS.n4333 VSS.n4332 0.0132571
R24889 VSS.n4419 VSS.n4417 0.0132571
R24890 VSS.n4447 VSS.n4002 0.0132571
R24891 VSS.n4500 VSS.n4499 0.0132571
R24892 VSS.n4519 VSS.n4518 0.0132571
R24893 VSS.n4823 VSS.n4819 0.0132571
R24894 VSS.n4925 VSS.n4924 0.0132571
R24895 VSS.n5011 VSS.n5009 0.0132571
R24896 VSS.n5039 VSS.n4594 0.0132571
R24897 VSS.n5092 VSS.n5091 0.0132571
R24898 VSS.n5111 VSS.n5110 0.0132571
R24899 VSS.n5415 VSS.n5411 0.0132571
R24900 VSS.n5517 VSS.n5516 0.0132571
R24901 VSS.n5603 VSS.n5601 0.0132571
R24902 VSS.n5631 VSS.n5186 0.0132571
R24903 VSS.n5684 VSS.n5683 0.0132571
R24904 VSS.n5703 VSS.n5702 0.0132571
R24905 VSS.n6007 VSS.n6003 0.0132571
R24906 VSS.n6109 VSS.n6108 0.0132571
R24907 VSS.n6195 VSS.n6193 0.0132571
R24908 VSS.n6223 VSS.n5778 0.0132571
R24909 VSS.n6276 VSS.n6275 0.0132571
R24910 VSS.n6295 VSS.n6294 0.0132571
R24911 VSS.n6599 VSS.n6595 0.0132571
R24912 VSS.n6701 VSS.n6700 0.0132571
R24913 VSS.n6787 VSS.n6785 0.0132571
R24914 VSS.n6815 VSS.n6370 0.0132571
R24915 VSS.n6868 VSS.n6867 0.0132571
R24916 VSS.n6887 VSS.n6886 0.0132571
R24917 VSS.n2443 VSS.n2439 0.0132571
R24918 VSS.n7024 VSS.n7023 0.0132571
R24919 VSS.n2652 VSS.n2651 0.0132571
R24920 VSS.n2669 VSS.n2668 0.0132571
R24921 VSS.n6936 VSS.n2719 0.0132571
R24922 VSS.n6934 VSS.n2720 0.0132571
R24923 VSS.n3044 VSS.n3043 0.0132571
R24924 VSS.n3149 VSS.n3148 0.0132571
R24925 VSS.n3235 VSS.n3233 0.0132571
R24926 VSS.n3263 VSS.n2817 0.0132571
R24927 VSS.n3316 VSS.n3315 0.0132571
R24928 VSS.n3335 VSS.n3334 0.0132571
R24929 VSS.n415 VSS.n414 0.0132571
R24930 VSS.n9109 VSS.n9108 0.0132571
R24931 VSS.n9195 VSS.n9193 0.0132571
R24932 VSS.n9223 VSS.n84 0.0132571
R24933 VSS.n9276 VSS.n9275 0.0132571
R24934 VSS.n9295 VSS.n9294 0.0132571
R24935 VSS.n980 VSS.n979 0.0132571
R24936 VSS.n843 VSS.n842 0.0132571
R24937 VSS.n644 VSS.n643 0.0132571
R24938 VSS.n661 VSS.n660 0.0132571
R24939 VSS.n755 VSS.n711 0.0132571
R24940 VSS.n753 VSS.n712 0.0132571
R24941 VSS.n8452 VSS.n8451 0.0132571
R24942 VSS.n7220 VSS.n7219 0.0132571
R24943 VSS.n7237 VSS.n7236 0.0132571
R24944 VSS.n8364 VSS.n7287 0.0132571
R24945 VSS.n8362 VSS.n7288 0.0132571
R24946 VSS.n7182 VSS.n7104 0.013
R24947 VSS.n8434 VSS.n8433 0.013
R24948 VSS.n7181 VSS.n7180 0.013
R24949 VSS.n999 VSS.n441 0.013
R24950 VSS.n899 VSS.n897 0.013
R24951 VSS.n7577 VSS.n7421 0.013
R24952 VSS.n7610 VSS.n7413 0.013
R24953 VSS.n8520 VSS.n1008 0.013
R24954 VSS.n1080 VSS.n1078 0.013
R24955 VSS.n1081 VSS.n1075 0.013
R24956 VSS.n7576 VSS.n7575 0.013
R24957 VSS.n8169 VSS.n7835 0.013
R24958 VSS.n8202 VSS.n7827 0.013
R24959 VSS.n7991 VSS.n7983 0.013
R24960 VSS.n7989 VSS.n7985 0.013
R24961 VSS.n7988 VSS.n7987 0.013
R24962 VSS.n8168 VSS.n8167 0.013
R24963 VSS.n8552 VSS.n8544 0.013
R24964 VSS.n8550 VSS.n8546 0.013
R24965 VSS.n8761 VSS.n8683 0.013
R24966 VSS.n9007 VSS.n9006 0.013
R24967 VSS.n8760 VSS.n8759 0.013
R24968 VSS.n8549 VSS.n8548 0.013
R24969 VSS.n1234 VSS.n1226 0.013
R24970 VSS.n1232 VSS.n1228 0.013
R24971 VSS.n1443 VSS.n1365 0.013
R24972 VSS.n1670 VSS.n1669 0.013
R24973 VSS.n1442 VSS.n1441 0.013
R24974 VSS.n1231 VSS.n1230 0.013
R24975 VSS.n1807 VSS.n1799 0.013
R24976 VSS.n1805 VSS.n1801 0.013
R24977 VSS.n2016 VSS.n1938 0.013
R24978 VSS.n2262 VSS.n2261 0.013
R24979 VSS.n2015 VSS.n2014 0.013
R24980 VSS.n1804 VSS.n1803 0.013
R24981 VSS.n3601 VSS.n3593 0.013
R24982 VSS.n3599 VSS.n3595 0.013
R24983 VSS.n3779 VSS.n3445 0.013
R24984 VSS.n3812 VSS.n3437 0.013
R24985 VSS.n3778 VSS.n3777 0.013
R24986 VSS.n3598 VSS.n3597 0.013
R24987 VSS.n4193 VSS.n4185 0.013
R24988 VSS.n4191 VSS.n4187 0.013
R24989 VSS.n4371 VSS.n4037 0.013
R24990 VSS.n4404 VSS.n4029 0.013
R24991 VSS.n4370 VSS.n4369 0.013
R24992 VSS.n4190 VSS.n4189 0.013
R24993 VSS.n4785 VSS.n4777 0.013
R24994 VSS.n4783 VSS.n4779 0.013
R24995 VSS.n4963 VSS.n4629 0.013
R24996 VSS.n4996 VSS.n4621 0.013
R24997 VSS.n4962 VSS.n4961 0.013
R24998 VSS.n4782 VSS.n4781 0.013
R24999 VSS.n5377 VSS.n5369 0.013
R25000 VSS.n5375 VSS.n5371 0.013
R25001 VSS.n5555 VSS.n5221 0.013
R25002 VSS.n5588 VSS.n5213 0.013
R25003 VSS.n5554 VSS.n5553 0.013
R25004 VSS.n5374 VSS.n5373 0.013
R25005 VSS.n5969 VSS.n5961 0.013
R25006 VSS.n5967 VSS.n5963 0.013
R25007 VSS.n6147 VSS.n5813 0.013
R25008 VSS.n6180 VSS.n5805 0.013
R25009 VSS.n6146 VSS.n6145 0.013
R25010 VSS.n5966 VSS.n5965 0.013
R25011 VSS.n6561 VSS.n6553 0.013
R25012 VSS.n6559 VSS.n6555 0.013
R25013 VSS.n6739 VSS.n6405 0.013
R25014 VSS.n6772 VSS.n6397 0.013
R25015 VSS.n6738 VSS.n6737 0.013
R25016 VSS.n6558 VSS.n6557 0.013
R25017 VSS.n2405 VSS.n2397 0.013
R25018 VSS.n2403 VSS.n2399 0.013
R25019 VSS.n2614 VSS.n2536 0.013
R25020 VSS.n7006 VSS.n7005 0.013
R25021 VSS.n2613 VSS.n2612 0.013
R25022 VSS.n2402 VSS.n2401 0.013
R25023 VSS.n3002 VSS.n2994 0.013
R25024 VSS.n3000 VSS.n2996 0.013
R25025 VSS.n3187 VSS.n2852 0.013
R25026 VSS.n3220 VSS.n2844 0.013
R25027 VSS.n3186 VSS.n3185 0.013
R25028 VSS.n2999 VSS.n2998 0.013
R25029 VSS.n434 VSS.n275 0.013
R25030 VSS.n333 VSS.n329 0.013
R25031 VSS.n9147 VSS.n119 0.013
R25032 VSS.n9180 VSS.n111 0.013
R25033 VSS.n9146 VSS.n9145 0.013
R25034 VSS.n335 VSS.n334 0.013
R25035 VSS.n606 VSS.n525 0.013
R25036 VSS.n825 VSS.n824 0.013
R25037 VSS.n605 VSS.n604 0.013
R25038 VSS.n900 VSS.n894 0.013
R25039 VSS.n8471 VSS.n7060 0.0121071
R25040 VSS.n7130 VSS.n7128 0.0121071
R25041 VSS.n7131 VSS.n7125 0.0121071
R25042 VSS.n7105 VSS.n7091 0.0121071
R25043 VSS.n903 VSS.n447 0.0121071
R25044 VSS.n950 VSS.n872 0.0121071
R25045 VSS.n962 VSS.n961 0.0121071
R25046 VSS.n7497 VSS.n7489 0.0121071
R25047 VSS.n7495 VSS.n7491 0.0121071
R25048 VSS.n1084 VSS.n1014 0.0121071
R25049 VSS.n1131 VSS.n1053 0.0121071
R25050 VSS.n8483 VSS.n8482 0.0121071
R25051 VSS.n1083 VSS.n1012 0.0121071
R25052 VSS.n1130 VSS.n1129 0.0121071
R25053 VSS.n7617 VSS.n7409 0.0121071
R25054 VSS.n7494 VSS.n7493 0.0121071
R25055 VSS.n7428 VSS.n7425 0.0121071
R25056 VSS.n8089 VSS.n8081 0.0121071
R25057 VSS.n8087 VSS.n8083 0.0121071
R25058 VSS.n7998 VSS.n7997 0.0121071
R25059 VSS.n8061 VSS.n8060 0.0121071
R25060 VSS.n8076 VSS.n7902 0.0121071
R25061 VSS.n7996 VSS.n7964 0.0121071
R25062 VSS.n8062 VSS.n7912 0.0121071
R25063 VSS.n8209 VSS.n7823 0.0121071
R25064 VSS.n8086 VSS.n8085 0.0121071
R25065 VSS.n7842 VSS.n7839 0.0121071
R25066 VSS.n8559 VSS.n8558 0.0121071
R25067 VSS.n8622 VSS.n8621 0.0121071
R25068 VSS.n8637 VSS.n199 0.0121071
R25069 VSS.n9044 VSS.n196 0.0121071
R25070 VSS.n8709 VSS.n8707 0.0121071
R25071 VSS.n8710 VSS.n8704 0.0121071
R25072 VSS.n8684 VSS.n8670 0.0121071
R25073 VSS.n8795 VSS.n8786 0.0121071
R25074 VSS.n8557 VSS.n261 0.0121071
R25075 VSS.n8623 VSS.n209 0.0121071
R25076 VSS.n1241 VSS.n1240 0.0121071
R25077 VSS.n1304 VSS.n1303 0.0121071
R25078 VSS.n1319 VSS.n1145 0.0121071
R25079 VSS.n1707 VSS.n1142 0.0121071
R25080 VSS.n1391 VSS.n1389 0.0121071
R25081 VSS.n1392 VSS.n1386 0.0121071
R25082 VSS.n1366 VSS.n1352 0.0121071
R25083 VSS.n1476 VSS.n1467 0.0121071
R25084 VSS.n1239 VSS.n1207 0.0121071
R25085 VSS.n1305 VSS.n1155 0.0121071
R25086 VSS.n1814 VSS.n1813 0.0121071
R25087 VSS.n1877 VSS.n1876 0.0121071
R25088 VSS.n1892 VSS.n1718 0.0121071
R25089 VSS.n2299 VSS.n1715 0.0121071
R25090 VSS.n1964 VSS.n1962 0.0121071
R25091 VSS.n1965 VSS.n1959 0.0121071
R25092 VSS.n1939 VSS.n1925 0.0121071
R25093 VSS.n2049 VSS.n2040 0.0121071
R25094 VSS.n1812 VSS.n1780 0.0121071
R25095 VSS.n1878 VSS.n1728 0.0121071
R25096 VSS.n3608 VSS.n3607 0.0121071
R25097 VSS.n3671 VSS.n3670 0.0121071
R25098 VSS.n3686 VSS.n3512 0.0121071
R25099 VSS.n3699 VSS.n3691 0.0121071
R25100 VSS.n3697 VSS.n3693 0.0121071
R25101 VSS.n3696 VSS.n3695 0.0121071
R25102 VSS.n3452 VSS.n3449 0.0121071
R25103 VSS.n3819 VSS.n3433 0.0121071
R25104 VSS.n3606 VSS.n3574 0.0121071
R25105 VSS.n3672 VSS.n3522 0.0121071
R25106 VSS.n4200 VSS.n4199 0.0121071
R25107 VSS.n4263 VSS.n4262 0.0121071
R25108 VSS.n4278 VSS.n4104 0.0121071
R25109 VSS.n4291 VSS.n4283 0.0121071
R25110 VSS.n4289 VSS.n4285 0.0121071
R25111 VSS.n4288 VSS.n4287 0.0121071
R25112 VSS.n4044 VSS.n4041 0.0121071
R25113 VSS.n4411 VSS.n4025 0.0121071
R25114 VSS.n4198 VSS.n4166 0.0121071
R25115 VSS.n4264 VSS.n4114 0.0121071
R25116 VSS.n4792 VSS.n4791 0.0121071
R25117 VSS.n4855 VSS.n4854 0.0121071
R25118 VSS.n4870 VSS.n4696 0.0121071
R25119 VSS.n4883 VSS.n4875 0.0121071
R25120 VSS.n4881 VSS.n4877 0.0121071
R25121 VSS.n4880 VSS.n4879 0.0121071
R25122 VSS.n4636 VSS.n4633 0.0121071
R25123 VSS.n5003 VSS.n4617 0.0121071
R25124 VSS.n4790 VSS.n4758 0.0121071
R25125 VSS.n4856 VSS.n4706 0.0121071
R25126 VSS.n5384 VSS.n5383 0.0121071
R25127 VSS.n5447 VSS.n5446 0.0121071
R25128 VSS.n5462 VSS.n5288 0.0121071
R25129 VSS.n5475 VSS.n5467 0.0121071
R25130 VSS.n5473 VSS.n5469 0.0121071
R25131 VSS.n5472 VSS.n5471 0.0121071
R25132 VSS.n5228 VSS.n5225 0.0121071
R25133 VSS.n5595 VSS.n5209 0.0121071
R25134 VSS.n5382 VSS.n5350 0.0121071
R25135 VSS.n5448 VSS.n5298 0.0121071
R25136 VSS.n5976 VSS.n5975 0.0121071
R25137 VSS.n6039 VSS.n6038 0.0121071
R25138 VSS.n6054 VSS.n5880 0.0121071
R25139 VSS.n6067 VSS.n6059 0.0121071
R25140 VSS.n6065 VSS.n6061 0.0121071
R25141 VSS.n6064 VSS.n6063 0.0121071
R25142 VSS.n5820 VSS.n5817 0.0121071
R25143 VSS.n6187 VSS.n5801 0.0121071
R25144 VSS.n5974 VSS.n5942 0.0121071
R25145 VSS.n6040 VSS.n5890 0.0121071
R25146 VSS.n6568 VSS.n6567 0.0121071
R25147 VSS.n6631 VSS.n6630 0.0121071
R25148 VSS.n6646 VSS.n6472 0.0121071
R25149 VSS.n6659 VSS.n6651 0.0121071
R25150 VSS.n6657 VSS.n6653 0.0121071
R25151 VSS.n6656 VSS.n6655 0.0121071
R25152 VSS.n6412 VSS.n6409 0.0121071
R25153 VSS.n6779 VSS.n6393 0.0121071
R25154 VSS.n6566 VSS.n6534 0.0121071
R25155 VSS.n6632 VSS.n6482 0.0121071
R25156 VSS.n2412 VSS.n2411 0.0121071
R25157 VSS.n2475 VSS.n2474 0.0121071
R25158 VSS.n2490 VSS.n2316 0.0121071
R25159 VSS.n7043 VSS.n2313 0.0121071
R25160 VSS.n2562 VSS.n2560 0.0121071
R25161 VSS.n2563 VSS.n2557 0.0121071
R25162 VSS.n2537 VSS.n2523 0.0121071
R25163 VSS.n2647 VSS.n2638 0.0121071
R25164 VSS.n2410 VSS.n2378 0.0121071
R25165 VSS.n2476 VSS.n2326 0.0121071
R25166 VSS.n3009 VSS.n3008 0.0121071
R25167 VSS.n3083 VSS.n2927 0.0121071
R25168 VSS.n3094 VSS.n2919 0.0121071
R25169 VSS.n3107 VSS.n3099 0.0121071
R25170 VSS.n3105 VSS.n3101 0.0121071
R25171 VSS.n3104 VSS.n3103 0.0121071
R25172 VSS.n2859 VSS.n2856 0.0121071
R25173 VSS.n3227 VSS.n2840 0.0121071
R25174 VSS.n3007 VSS.n2977 0.0121071
R25175 VSS.n3082 VSS.n3081 0.0121071
R25176 VSS.n330 VSS.n281 0.0121071
R25177 VSS.n395 VSS.n394 0.0121071
R25178 VSS.n9054 VSS.n179 0.0121071
R25179 VSS.n9067 VSS.n9059 0.0121071
R25180 VSS.n9065 VSS.n9061 0.0121071
R25181 VSS.n9064 VSS.n9063 0.0121071
R25182 VSS.n126 VSS.n123 0.0121071
R25183 VSS.n9187 VSS.n107 0.0121071
R25184 VSS.n336 VSS.n279 0.0121071
R25185 VSS.n393 VSS.n308 0.0121071
R25186 VSS.n861 VSS.n860 0.0121071
R25187 VSS.n554 VSS.n552 0.0121071
R25188 VSS.n555 VSS.n551 0.0121071
R25189 VSS.n526 VSS.n512 0.0121071
R25190 VSS.n639 VSS.n630 0.0121071
R25191 VSS.n902 VSS.n445 0.0121071
R25192 VSS.n949 VSS.n948 0.0121071
R25193 VSS.n7215 VSS.n7206 0.0121071
R25194 VSS.n7130 VSS.n7129 0.0112143
R25195 VSS.n7134 VSS.n7066 0.0112143
R25196 VSS.n7106 VSS.n7090 0.0112143
R25197 VSS.n7133 VSS.n7064 0.0112143
R25198 VSS.n951 VSS.n950 0.0112143
R25199 VSS.n7491 VSS.n7490 0.0112143
R25200 VSS.n7504 VSS.n7503 0.0112143
R25201 VSS.n7567 VSS.n7566 0.0112143
R25202 VSS.n1132 VSS.n1131 0.0112143
R25203 VSS.n1054 VSS.n1040 0.0112143
R25204 VSS.n7660 VSS.n7659 0.0112143
R25205 VSS.n7682 VSS.n7681 0.0112143
R25206 VSS.n7711 VSS.n7364 0.0112143
R25207 VSS.n7728 VSS.n7342 0.0112143
R25208 VSS.n7710 VSS.n7709 0.0112143
R25209 VSS.n7502 VSS.n7471 0.0112143
R25210 VSS.n8083 VSS.n8082 0.0112143
R25211 VSS.n8096 VSS.n8095 0.0112143
R25212 VSS.n8159 VSS.n8158 0.0112143
R25213 VSS.n8061 VSS.n7917 0.0112143
R25214 VSS.n8064 VSS.n7911 0.0112143
R25215 VSS.n8252 VSS.n8251 0.0112143
R25216 VSS.n8274 VSS.n8273 0.0112143
R25217 VSS.n8303 VSS.n7778 0.0112143
R25218 VSS.n8320 VSS.n7756 0.0112143
R25219 VSS.n8302 VSS.n8301 0.0112143
R25220 VSS.n8094 VSS.n7885 0.0112143
R25221 VSS.n8622 VSS.n214 0.0112143
R25222 VSS.n8709 VSS.n8708 0.0112143
R25223 VSS.n8713 VSS.n8645 0.0112143
R25224 VSS.n8685 VSS.n8669 0.0112143
R25225 VSS.n8712 VSS.n8643 0.0112143
R25226 VSS.n8841 VSS.n8808 0.0112143
R25227 VSS.n8871 VSS.n8870 0.0112143
R25228 VSS.n8909 VSS.n8881 0.0112143
R25229 VSS.n8897 VSS.n8896 0.0112143
R25230 VSS.n8908 VSS.n8879 0.0112143
R25231 VSS.n8625 VSS.n208 0.0112143
R25232 VSS.n1304 VSS.n1160 0.0112143
R25233 VSS.n1391 VSS.n1390 0.0112143
R25234 VSS.n1395 VSS.n1327 0.0112143
R25235 VSS.n1367 VSS.n1351 0.0112143
R25236 VSS.n1394 VSS.n1325 0.0112143
R25237 VSS.n1521 VSS.n1520 0.0112143
R25238 VSS.n1577 VSS.n1535 0.0112143
R25239 VSS.n1604 VSS.n1603 0.0112143
R25240 VSS.n1557 VSS.n4 0.0112143
R25241 VSS.n1605 VSS.n1541 0.0112143
R25242 VSS.n1307 VSS.n1154 0.0112143
R25243 VSS.n1877 VSS.n1733 0.0112143
R25244 VSS.n1964 VSS.n1963 0.0112143
R25245 VSS.n1968 VSS.n1900 0.0112143
R25246 VSS.n1940 VSS.n1924 0.0112143
R25247 VSS.n1967 VSS.n1898 0.0112143
R25248 VSS.n2094 VSS.n2093 0.0112143
R25249 VSS.n2137 VSS.n2108 0.0112143
R25250 VSS.n2196 VSS.n2195 0.0112143
R25251 VSS.n2177 VSS.n2153 0.0112143
R25252 VSS.n2197 VSS.n2114 0.0112143
R25253 VSS.n1880 VSS.n1727 0.0112143
R25254 VSS.n3671 VSS.n3527 0.0112143
R25255 VSS.n3693 VSS.n3692 0.0112143
R25256 VSS.n3706 VSS.n3705 0.0112143
R25257 VSS.n3769 VSS.n3768 0.0112143
R25258 VSS.n3704 VSS.n3495 0.0112143
R25259 VSS.n3862 VSS.n3861 0.0112143
R25260 VSS.n3884 VSS.n3883 0.0112143
R25261 VSS.n3913 VSS.n3388 0.0112143
R25262 VSS.n3931 VSS.n3367 0.0112143
R25263 VSS.n3912 VSS.n3911 0.0112143
R25264 VSS.n3674 VSS.n3521 0.0112143
R25265 VSS.n4263 VSS.n4119 0.0112143
R25266 VSS.n4285 VSS.n4284 0.0112143
R25267 VSS.n4298 VSS.n4297 0.0112143
R25268 VSS.n4361 VSS.n4360 0.0112143
R25269 VSS.n4296 VSS.n4087 0.0112143
R25270 VSS.n4454 VSS.n4453 0.0112143
R25271 VSS.n4476 VSS.n4475 0.0112143
R25272 VSS.n4505 VSS.n3980 0.0112143
R25273 VSS.n4523 VSS.n3959 0.0112143
R25274 VSS.n4504 VSS.n4503 0.0112143
R25275 VSS.n4266 VSS.n4113 0.0112143
R25276 VSS.n4855 VSS.n4711 0.0112143
R25277 VSS.n4877 VSS.n4876 0.0112143
R25278 VSS.n4890 VSS.n4889 0.0112143
R25279 VSS.n4953 VSS.n4952 0.0112143
R25280 VSS.n4888 VSS.n4679 0.0112143
R25281 VSS.n5046 VSS.n5045 0.0112143
R25282 VSS.n5068 VSS.n5067 0.0112143
R25283 VSS.n5097 VSS.n4572 0.0112143
R25284 VSS.n5115 VSS.n4551 0.0112143
R25285 VSS.n5096 VSS.n5095 0.0112143
R25286 VSS.n4858 VSS.n4705 0.0112143
R25287 VSS.n5447 VSS.n5303 0.0112143
R25288 VSS.n5469 VSS.n5468 0.0112143
R25289 VSS.n5482 VSS.n5481 0.0112143
R25290 VSS.n5545 VSS.n5544 0.0112143
R25291 VSS.n5480 VSS.n5271 0.0112143
R25292 VSS.n5638 VSS.n5637 0.0112143
R25293 VSS.n5660 VSS.n5659 0.0112143
R25294 VSS.n5689 VSS.n5164 0.0112143
R25295 VSS.n5707 VSS.n5143 0.0112143
R25296 VSS.n5688 VSS.n5687 0.0112143
R25297 VSS.n5450 VSS.n5297 0.0112143
R25298 VSS.n6039 VSS.n5895 0.0112143
R25299 VSS.n6061 VSS.n6060 0.0112143
R25300 VSS.n6074 VSS.n6073 0.0112143
R25301 VSS.n6137 VSS.n6136 0.0112143
R25302 VSS.n6072 VSS.n5863 0.0112143
R25303 VSS.n6230 VSS.n6229 0.0112143
R25304 VSS.n6252 VSS.n6251 0.0112143
R25305 VSS.n6281 VSS.n5756 0.0112143
R25306 VSS.n6299 VSS.n5735 0.0112143
R25307 VSS.n6280 VSS.n6279 0.0112143
R25308 VSS.n6042 VSS.n5889 0.0112143
R25309 VSS.n6631 VSS.n6487 0.0112143
R25310 VSS.n6653 VSS.n6652 0.0112143
R25311 VSS.n6666 VSS.n6665 0.0112143
R25312 VSS.n6729 VSS.n6728 0.0112143
R25313 VSS.n6664 VSS.n6455 0.0112143
R25314 VSS.n6822 VSS.n6821 0.0112143
R25315 VSS.n6844 VSS.n6843 0.0112143
R25316 VSS.n6873 VSS.n6348 0.0112143
R25317 VSS.n6891 VSS.n6327 0.0112143
R25318 VSS.n6872 VSS.n6871 0.0112143
R25319 VSS.n6634 VSS.n6481 0.0112143
R25320 VSS.n2475 VSS.n2331 0.0112143
R25321 VSS.n2562 VSS.n2561 0.0112143
R25322 VSS.n2566 VSS.n2498 0.0112143
R25323 VSS.n2538 VSS.n2522 0.0112143
R25324 VSS.n2565 VSS.n2496 0.0112143
R25325 VSS.n2692 VSS.n2691 0.0112143
R25326 VSS.n2735 VSS.n2706 0.0112143
R25327 VSS.n6940 VSS.n6939 0.0112143
R25328 VSS.n6921 VSS.n2751 0.0112143
R25329 VSS.n6941 VSS.n2712 0.0112143
R25330 VSS.n2478 VSS.n2325 0.0112143
R25331 VSS.n3084 VSS.n3083 0.0112143
R25332 VSS.n3101 VSS.n3100 0.0112143
R25333 VSS.n3114 VSS.n3113 0.0112143
R25334 VSS.n3177 VSS.n3176 0.0112143
R25335 VSS.n3112 VSS.n2902 0.0112143
R25336 VSS.n3270 VSS.n3269 0.0112143
R25337 VSS.n3292 VSS.n3291 0.0112143
R25338 VSS.n3321 VSS.n2795 0.0112143
R25339 VSS.n3339 VSS.n2774 0.0112143
R25340 VSS.n3320 VSS.n3319 0.0112143
R25341 VSS.n2934 VSS.n2931 0.0112143
R25342 VSS.n394 VSS.n309 0.0112143
R25343 VSS.n9061 VSS.n9060 0.0112143
R25344 VSS.n9074 VSS.n9073 0.0112143
R25345 VSS.n9137 VSS.n9136 0.0112143
R25346 VSS.n9072 VSS.n169 0.0112143
R25347 VSS.n9230 VSS.n9229 0.0112143
R25348 VSS.n9252 VSS.n9251 0.0112143
R25349 VSS.n9281 VSS.n62 0.0112143
R25350 VSS.n9299 VSS.n41 0.0112143
R25351 VSS.n9280 VSS.n9279 0.0112143
R25352 VSS.n310 VSS.n307 0.0112143
R25353 VSS.n554 VSS.n553 0.0112143
R25354 VSS.n558 VSS.n487 0.0112143
R25355 VSS.n527 VSS.n511 0.0112143
R25356 VSS.n557 VSS.n485 0.0112143
R25357 VSS.n684 VSS.n683 0.0112143
R25358 VSS.n736 VSS.n698 0.0112143
R25359 VSS.n759 VSS.n758 0.0112143
R25360 VSS.n9328 VSS.n33 0.0112143
R25361 VSS.n760 VSS.n704 0.0112143
R25362 VSS.n873 VSS.n473 0.0112143
R25363 VSS.n7260 VSS.n7259 0.0112143
R25364 VSS.n7303 VSS.n7274 0.0112143
R25365 VSS.n8368 VSS.n8367 0.0112143
R25366 VSS.n8349 VSS.n7319 0.0112143
R25367 VSS.n8369 VSS.n7280 0.0112143
R25368 VSS.n7134 VSS.n7124 0.0103214
R25369 VSS.n8464 VSS.n8463 0.0103214
R25370 VSS.n8457 VSS.n7072 0.0103214
R25371 VSS.n7161 VSS.n7081 0.0103214
R25372 VSS.n7183 VSS.n7182 0.0103214
R25373 VSS.n7133 VSS.n7132 0.0103214
R25374 VSS.n8458 VSS.n7070 0.0103214
R25375 VSS.n8454 VSS.n7075 0.0103214
R25376 VSS.n8445 VSS.n7084 0.0103214
R25377 VSS.n7165 VSS.n7087 0.0103214
R25378 VSS.n899 VSS.n898 0.0103214
R25379 VSS.n985 VSS.n453 0.0103214
R25380 VSS.n928 VSS.n463 0.0103214
R25381 VSS.n968 VSS.n967 0.0103214
R25382 VSS.n874 VSS.n472 0.0103214
R25383 VSS.n946 VSS.n945 0.0103214
R25384 VSS.n7504 VSS.n7470 0.0103214
R25385 VSS.n7473 VSS.n7472 0.0103214
R25386 VSS.n7524 VSS.n7457 0.0103214
R25387 VSS.n7545 VSS.n7436 0.0103214
R25388 VSS.n7578 VSS.n7577 0.0103214
R25389 VSS.n1080 VSS.n1079 0.0103214
R25390 VSS.n8506 VSS.n1020 0.0103214
R25391 VSS.n1109 VSS.n1030 0.0103214
R25392 VSS.n8489 VSS.n8488 0.0103214
R25393 VSS.n1055 VSS.n1039 0.0103214
R25394 VSS.n1127 VSS.n1126 0.0103214
R25395 VSS.n8507 VSS.n1018 0.0103214
R25396 VSS.n1031 VSS.n1028 0.0103214
R25397 VSS.n8494 VSS.n1033 0.0103214
R25398 VSS.n1128 VSS.n1054 0.0103214
R25399 VSS.n7628 VSS.n7402 0.0103214
R25400 VSS.n7632 VSS.n7400 0.0103214
R25401 VSS.n7634 VSS.n7398 0.0103214
R25402 VSS.n7627 VSS.n7404 0.0103214
R25403 VSS.n7636 VSS.n7635 0.0103214
R25404 VSS.n7492 VSS.n7471 0.0103214
R25405 VSS.n7523 VSS.n7522 0.0103214
R25406 VSS.n7518 VSS.n7446 0.0103214
R25407 VSS.n7546 VSS.n7438 0.0103214
R25408 VSS.n7554 VSS.n7553 0.0103214
R25409 VSS.n8096 VSS.n7884 0.0103214
R25410 VSS.n7887 VSS.n7886 0.0103214
R25411 VSS.n8116 VSS.n7871 0.0103214
R25412 VSS.n8137 VSS.n7850 0.0103214
R25413 VSS.n8170 VSS.n8169 0.0103214
R25414 VSS.n7985 VSS.n7984 0.0103214
R25415 VSS.n7954 VSS.n7947 0.0103214
R25416 VSS.n8046 VSS.n8045 0.0103214
R25417 VSS.n8053 VSS.n8052 0.0103214
R25418 VSS.n8066 VSS.n7909 0.0103214
R25419 VSS.n8065 VSS.n7910 0.0103214
R25420 VSS.n7953 VSS.n7948 0.0103214
R25421 VSS.n8027 VSS.n7944 0.0103214
R25422 VSS.n8047 VSS.n7924 0.0103214
R25423 VSS.n8064 VSS.n8063 0.0103214
R25424 VSS.n8220 VSS.n7816 0.0103214
R25425 VSS.n8224 VSS.n7814 0.0103214
R25426 VSS.n8226 VSS.n7812 0.0103214
R25427 VSS.n8219 VSS.n7818 0.0103214
R25428 VSS.n8228 VSS.n8227 0.0103214
R25429 VSS.n8084 VSS.n7885 0.0103214
R25430 VSS.n8115 VSS.n8114 0.0103214
R25431 VSS.n8110 VSS.n7860 0.0103214
R25432 VSS.n8138 VSS.n7852 0.0103214
R25433 VSS.n8146 VSS.n8145 0.0103214
R25434 VSS.n8546 VSS.n8545 0.0103214
R25435 VSS.n251 VSS.n244 0.0103214
R25436 VSS.n8607 VSS.n8606 0.0103214
R25437 VSS.n8614 VSS.n8613 0.0103214
R25438 VSS.n8627 VSS.n206 0.0103214
R25439 VSS.n8626 VSS.n207 0.0103214
R25440 VSS.n8713 VSS.n8703 0.0103214
R25441 VSS.n9037 VSS.n9036 0.0103214
R25442 VSS.n9030 VSS.n8651 0.0103214
R25443 VSS.n8740 VSS.n8660 0.0103214
R25444 VSS.n8762 VSS.n8761 0.0103214
R25445 VSS.n8712 VSS.n8711 0.0103214
R25446 VSS.n9031 VSS.n8649 0.0103214
R25447 VSS.n9027 VSS.n8654 0.0103214
R25448 VSS.n9018 VSS.n8663 0.0103214
R25449 VSS.n8744 VSS.n8666 0.0103214
R25450 VSS.n8989 VSS.n8988 0.0103214
R25451 VSS.n8826 VSS.n8802 0.0103214
R25452 VSS.n8980 VSS.n8979 0.0103214
R25453 VSS.n8987 VSS.n8778 0.0103214
R25454 VSS.n8978 VSS.n8801 0.0103214
R25455 VSS.n250 VSS.n245 0.0103214
R25456 VSS.n8588 VSS.n241 0.0103214
R25457 VSS.n8608 VSS.n221 0.0103214
R25458 VSS.n8625 VSS.n8624 0.0103214
R25459 VSS.n1228 VSS.n1227 0.0103214
R25460 VSS.n1197 VSS.n1190 0.0103214
R25461 VSS.n1289 VSS.n1288 0.0103214
R25462 VSS.n1296 VSS.n1295 0.0103214
R25463 VSS.n1309 VSS.n1152 0.0103214
R25464 VSS.n1308 VSS.n1153 0.0103214
R25465 VSS.n1395 VSS.n1385 0.0103214
R25466 VSS.n1700 VSS.n1699 0.0103214
R25467 VSS.n1693 VSS.n1333 0.0103214
R25468 VSS.n1422 VSS.n1342 0.0103214
R25469 VSS.n1444 VSS.n1443 0.0103214
R25470 VSS.n1394 VSS.n1393 0.0103214
R25471 VSS.n1694 VSS.n1331 0.0103214
R25472 VSS.n1690 VSS.n1336 0.0103214
R25473 VSS.n1681 VSS.n1345 0.0103214
R25474 VSS.n1426 VSS.n1348 0.0103214
R25475 VSS.n1652 VSS.n1460 0.0103214
R25476 VSS.n1647 VSS.n1482 0.0103214
R25477 VSS.n1494 VSS.n1488 0.0103214
R25478 VSS.n1651 VSS.n1650 0.0103214
R25479 VSS.n1493 VSS.n1490 0.0103214
R25480 VSS.n1196 VSS.n1191 0.0103214
R25481 VSS.n1270 VSS.n1187 0.0103214
R25482 VSS.n1290 VSS.n1167 0.0103214
R25483 VSS.n1307 VSS.n1306 0.0103214
R25484 VSS.n1801 VSS.n1800 0.0103214
R25485 VSS.n1770 VSS.n1763 0.0103214
R25486 VSS.n1862 VSS.n1861 0.0103214
R25487 VSS.n1869 VSS.n1868 0.0103214
R25488 VSS.n1882 VSS.n1725 0.0103214
R25489 VSS.n1881 VSS.n1726 0.0103214
R25490 VSS.n1968 VSS.n1958 0.0103214
R25491 VSS.n2292 VSS.n2291 0.0103214
R25492 VSS.n2285 VSS.n1906 0.0103214
R25493 VSS.n1995 VSS.n1915 0.0103214
R25494 VSS.n2017 VSS.n2016 0.0103214
R25495 VSS.n1967 VSS.n1966 0.0103214
R25496 VSS.n2286 VSS.n1904 0.0103214
R25497 VSS.n2282 VSS.n1909 0.0103214
R25498 VSS.n2273 VSS.n1918 0.0103214
R25499 VSS.n1999 VSS.n1921 0.0103214
R25500 VSS.n2244 VSS.n2033 0.0103214
R25501 VSS.n2239 VSS.n2055 0.0103214
R25502 VSS.n2067 VSS.n2061 0.0103214
R25503 VSS.n2243 VSS.n2242 0.0103214
R25504 VSS.n2066 VSS.n2063 0.0103214
R25505 VSS.n1769 VSS.n1764 0.0103214
R25506 VSS.n1843 VSS.n1760 0.0103214
R25507 VSS.n1863 VSS.n1740 0.0103214
R25508 VSS.n1880 VSS.n1879 0.0103214
R25509 VSS.n3595 VSS.n3594 0.0103214
R25510 VSS.n3564 VSS.n3557 0.0103214
R25511 VSS.n3656 VSS.n3655 0.0103214
R25512 VSS.n3663 VSS.n3662 0.0103214
R25513 VSS.n3676 VSS.n3519 0.0103214
R25514 VSS.n3675 VSS.n3520 0.0103214
R25515 VSS.n3706 VSS.n3494 0.0103214
R25516 VSS.n3497 VSS.n3496 0.0103214
R25517 VSS.n3726 VSS.n3481 0.0103214
R25518 VSS.n3747 VSS.n3460 0.0103214
R25519 VSS.n3780 VSS.n3779 0.0103214
R25520 VSS.n3694 VSS.n3495 0.0103214
R25521 VSS.n3725 VSS.n3724 0.0103214
R25522 VSS.n3720 VSS.n3470 0.0103214
R25523 VSS.n3748 VSS.n3462 0.0103214
R25524 VSS.n3756 VSS.n3755 0.0103214
R25525 VSS.n3830 VSS.n3426 0.0103214
R25526 VSS.n3834 VSS.n3424 0.0103214
R25527 VSS.n3836 VSS.n3422 0.0103214
R25528 VSS.n3829 VSS.n3428 0.0103214
R25529 VSS.n3838 VSS.n3837 0.0103214
R25530 VSS.n3563 VSS.n3558 0.0103214
R25531 VSS.n3637 VSS.n3554 0.0103214
R25532 VSS.n3657 VSS.n3534 0.0103214
R25533 VSS.n3674 VSS.n3673 0.0103214
R25534 VSS.n4187 VSS.n4186 0.0103214
R25535 VSS.n4156 VSS.n4149 0.0103214
R25536 VSS.n4248 VSS.n4247 0.0103214
R25537 VSS.n4255 VSS.n4254 0.0103214
R25538 VSS.n4268 VSS.n4111 0.0103214
R25539 VSS.n4267 VSS.n4112 0.0103214
R25540 VSS.n4298 VSS.n4086 0.0103214
R25541 VSS.n4089 VSS.n4088 0.0103214
R25542 VSS.n4318 VSS.n4073 0.0103214
R25543 VSS.n4339 VSS.n4052 0.0103214
R25544 VSS.n4372 VSS.n4371 0.0103214
R25545 VSS.n4286 VSS.n4087 0.0103214
R25546 VSS.n4317 VSS.n4316 0.0103214
R25547 VSS.n4312 VSS.n4062 0.0103214
R25548 VSS.n4340 VSS.n4054 0.0103214
R25549 VSS.n4348 VSS.n4347 0.0103214
R25550 VSS.n4422 VSS.n4018 0.0103214
R25551 VSS.n4426 VSS.n4016 0.0103214
R25552 VSS.n4428 VSS.n4014 0.0103214
R25553 VSS.n4421 VSS.n4020 0.0103214
R25554 VSS.n4430 VSS.n4429 0.0103214
R25555 VSS.n4155 VSS.n4150 0.0103214
R25556 VSS.n4229 VSS.n4146 0.0103214
R25557 VSS.n4249 VSS.n4126 0.0103214
R25558 VSS.n4266 VSS.n4265 0.0103214
R25559 VSS.n4779 VSS.n4778 0.0103214
R25560 VSS.n4748 VSS.n4741 0.0103214
R25561 VSS.n4840 VSS.n4839 0.0103214
R25562 VSS.n4847 VSS.n4846 0.0103214
R25563 VSS.n4860 VSS.n4703 0.0103214
R25564 VSS.n4859 VSS.n4704 0.0103214
R25565 VSS.n4890 VSS.n4678 0.0103214
R25566 VSS.n4681 VSS.n4680 0.0103214
R25567 VSS.n4910 VSS.n4665 0.0103214
R25568 VSS.n4931 VSS.n4644 0.0103214
R25569 VSS.n4964 VSS.n4963 0.0103214
R25570 VSS.n4878 VSS.n4679 0.0103214
R25571 VSS.n4909 VSS.n4908 0.0103214
R25572 VSS.n4904 VSS.n4654 0.0103214
R25573 VSS.n4932 VSS.n4646 0.0103214
R25574 VSS.n4940 VSS.n4939 0.0103214
R25575 VSS.n5014 VSS.n4610 0.0103214
R25576 VSS.n5018 VSS.n4608 0.0103214
R25577 VSS.n5020 VSS.n4606 0.0103214
R25578 VSS.n5013 VSS.n4612 0.0103214
R25579 VSS.n5022 VSS.n5021 0.0103214
R25580 VSS.n4747 VSS.n4742 0.0103214
R25581 VSS.n4821 VSS.n4738 0.0103214
R25582 VSS.n4841 VSS.n4718 0.0103214
R25583 VSS.n4858 VSS.n4857 0.0103214
R25584 VSS.n5371 VSS.n5370 0.0103214
R25585 VSS.n5340 VSS.n5333 0.0103214
R25586 VSS.n5432 VSS.n5431 0.0103214
R25587 VSS.n5439 VSS.n5438 0.0103214
R25588 VSS.n5452 VSS.n5295 0.0103214
R25589 VSS.n5451 VSS.n5296 0.0103214
R25590 VSS.n5482 VSS.n5270 0.0103214
R25591 VSS.n5273 VSS.n5272 0.0103214
R25592 VSS.n5502 VSS.n5257 0.0103214
R25593 VSS.n5523 VSS.n5236 0.0103214
R25594 VSS.n5556 VSS.n5555 0.0103214
R25595 VSS.n5470 VSS.n5271 0.0103214
R25596 VSS.n5501 VSS.n5500 0.0103214
R25597 VSS.n5496 VSS.n5246 0.0103214
R25598 VSS.n5524 VSS.n5238 0.0103214
R25599 VSS.n5532 VSS.n5531 0.0103214
R25600 VSS.n5606 VSS.n5202 0.0103214
R25601 VSS.n5610 VSS.n5200 0.0103214
R25602 VSS.n5612 VSS.n5198 0.0103214
R25603 VSS.n5605 VSS.n5204 0.0103214
R25604 VSS.n5614 VSS.n5613 0.0103214
R25605 VSS.n5339 VSS.n5334 0.0103214
R25606 VSS.n5413 VSS.n5330 0.0103214
R25607 VSS.n5433 VSS.n5310 0.0103214
R25608 VSS.n5450 VSS.n5449 0.0103214
R25609 VSS.n5963 VSS.n5962 0.0103214
R25610 VSS.n5932 VSS.n5925 0.0103214
R25611 VSS.n6024 VSS.n6023 0.0103214
R25612 VSS.n6031 VSS.n6030 0.0103214
R25613 VSS.n6044 VSS.n5887 0.0103214
R25614 VSS.n6043 VSS.n5888 0.0103214
R25615 VSS.n6074 VSS.n5862 0.0103214
R25616 VSS.n5865 VSS.n5864 0.0103214
R25617 VSS.n6094 VSS.n5849 0.0103214
R25618 VSS.n6115 VSS.n5828 0.0103214
R25619 VSS.n6148 VSS.n6147 0.0103214
R25620 VSS.n6062 VSS.n5863 0.0103214
R25621 VSS.n6093 VSS.n6092 0.0103214
R25622 VSS.n6088 VSS.n5838 0.0103214
R25623 VSS.n6116 VSS.n5830 0.0103214
R25624 VSS.n6124 VSS.n6123 0.0103214
R25625 VSS.n6198 VSS.n5794 0.0103214
R25626 VSS.n6202 VSS.n5792 0.0103214
R25627 VSS.n6204 VSS.n5790 0.0103214
R25628 VSS.n6197 VSS.n5796 0.0103214
R25629 VSS.n6206 VSS.n6205 0.0103214
R25630 VSS.n5931 VSS.n5926 0.0103214
R25631 VSS.n6005 VSS.n5922 0.0103214
R25632 VSS.n6025 VSS.n5902 0.0103214
R25633 VSS.n6042 VSS.n6041 0.0103214
R25634 VSS.n6555 VSS.n6554 0.0103214
R25635 VSS.n6524 VSS.n6517 0.0103214
R25636 VSS.n6616 VSS.n6615 0.0103214
R25637 VSS.n6623 VSS.n6622 0.0103214
R25638 VSS.n6636 VSS.n6479 0.0103214
R25639 VSS.n6635 VSS.n6480 0.0103214
R25640 VSS.n6666 VSS.n6454 0.0103214
R25641 VSS.n6457 VSS.n6456 0.0103214
R25642 VSS.n6686 VSS.n6441 0.0103214
R25643 VSS.n6707 VSS.n6420 0.0103214
R25644 VSS.n6740 VSS.n6739 0.0103214
R25645 VSS.n6654 VSS.n6455 0.0103214
R25646 VSS.n6685 VSS.n6684 0.0103214
R25647 VSS.n6680 VSS.n6430 0.0103214
R25648 VSS.n6708 VSS.n6422 0.0103214
R25649 VSS.n6716 VSS.n6715 0.0103214
R25650 VSS.n6790 VSS.n6386 0.0103214
R25651 VSS.n6794 VSS.n6384 0.0103214
R25652 VSS.n6796 VSS.n6382 0.0103214
R25653 VSS.n6789 VSS.n6388 0.0103214
R25654 VSS.n6798 VSS.n6797 0.0103214
R25655 VSS.n6523 VSS.n6518 0.0103214
R25656 VSS.n6597 VSS.n6514 0.0103214
R25657 VSS.n6617 VSS.n6494 0.0103214
R25658 VSS.n6634 VSS.n6633 0.0103214
R25659 VSS.n2399 VSS.n2398 0.0103214
R25660 VSS.n2368 VSS.n2361 0.0103214
R25661 VSS.n2460 VSS.n2459 0.0103214
R25662 VSS.n2467 VSS.n2466 0.0103214
R25663 VSS.n2480 VSS.n2323 0.0103214
R25664 VSS.n2479 VSS.n2324 0.0103214
R25665 VSS.n2566 VSS.n2556 0.0103214
R25666 VSS.n7036 VSS.n7035 0.0103214
R25667 VSS.n7029 VSS.n2504 0.0103214
R25668 VSS.n2593 VSS.n2513 0.0103214
R25669 VSS.n2615 VSS.n2614 0.0103214
R25670 VSS.n2565 VSS.n2564 0.0103214
R25671 VSS.n7030 VSS.n2502 0.0103214
R25672 VSS.n7026 VSS.n2507 0.0103214
R25673 VSS.n7017 VSS.n2516 0.0103214
R25674 VSS.n2597 VSS.n2519 0.0103214
R25675 VSS.n6988 VSS.n2631 0.0103214
R25676 VSS.n6983 VSS.n2653 0.0103214
R25677 VSS.n2665 VSS.n2659 0.0103214
R25678 VSS.n6987 VSS.n6986 0.0103214
R25679 VSS.n2664 VSS.n2661 0.0103214
R25680 VSS.n2367 VSS.n2362 0.0103214
R25681 VSS.n2441 VSS.n2358 0.0103214
R25682 VSS.n2461 VSS.n2338 0.0103214
R25683 VSS.n2478 VSS.n2477 0.0103214
R25684 VSS.n2996 VSS.n2995 0.0103214
R25685 VSS.n3029 VSS.n2965 0.0103214
R25686 VSS.n3050 VSS.n2942 0.0103214
R25687 VSS.n3074 VSS.n2932 0.0103214
R25688 VSS.n3073 VSS.n3072 0.0103214
R25689 VSS.n2935 VSS.n2933 0.0103214
R25690 VSS.n3114 VSS.n2901 0.0103214
R25691 VSS.n2904 VSS.n2903 0.0103214
R25692 VSS.n3134 VSS.n2888 0.0103214
R25693 VSS.n3155 VSS.n2867 0.0103214
R25694 VSS.n3188 VSS.n3187 0.0103214
R25695 VSS.n3102 VSS.n2902 0.0103214
R25696 VSS.n3133 VSS.n3132 0.0103214
R25697 VSS.n3128 VSS.n2877 0.0103214
R25698 VSS.n3156 VSS.n2869 0.0103214
R25699 VSS.n3164 VSS.n3163 0.0103214
R25700 VSS.n3238 VSS.n2833 0.0103214
R25701 VSS.n3242 VSS.n2831 0.0103214
R25702 VSS.n3244 VSS.n2829 0.0103214
R25703 VSS.n3237 VSS.n2835 0.0103214
R25704 VSS.n3246 VSS.n3245 0.0103214
R25705 VSS.n3028 VSS.n3027 0.0103214
R25706 VSS.n3047 VSS.n3046 0.0103214
R25707 VSS.n3051 VSS.n2944 0.0103214
R25708 VSS.n2934 VSS.n2928 0.0103214
R25709 VSS.n339 VSS.n329 0.0103214
R25710 VSS.n420 VSS.n287 0.0103214
R25711 VSS.n317 VSS.n297 0.0103214
R25712 VSS.n403 VSS.n402 0.0103214
R25713 VSS.n379 VSS.n306 0.0103214
R25714 VSS.n391 VSS.n311 0.0103214
R25715 VSS.n9074 VSS.n168 0.0103214
R25716 VSS.n171 VSS.n170 0.0103214
R25717 VSS.n9094 VSS.n155 0.0103214
R25718 VSS.n9115 VSS.n134 0.0103214
R25719 VSS.n9148 VSS.n9147 0.0103214
R25720 VSS.n9062 VSS.n169 0.0103214
R25721 VSS.n9093 VSS.n9092 0.0103214
R25722 VSS.n9088 VSS.n144 0.0103214
R25723 VSS.n9116 VSS.n136 0.0103214
R25724 VSS.n9124 VSS.n9123 0.0103214
R25725 VSS.n9198 VSS.n100 0.0103214
R25726 VSS.n9202 VSS.n98 0.0103214
R25727 VSS.n9204 VSS.n96 0.0103214
R25728 VSS.n9197 VSS.n102 0.0103214
R25729 VSS.n9206 VSS.n9205 0.0103214
R25730 VSS.n421 VSS.n285 0.0103214
R25731 VSS.n298 VSS.n295 0.0103214
R25732 VSS.n408 VSS.n300 0.0103214
R25733 VSS.n392 VSS.n310 0.0103214
R25734 VSS.n558 VSS.n550 0.0103214
R25735 VSS.n855 VSS.n854 0.0103214
R25736 VSS.n848 VSS.n493 0.0103214
R25737 VSS.n585 VSS.n502 0.0103214
R25738 VSS.n607 VSS.n606 0.0103214
R25739 VSS.n557 VSS.n556 0.0103214
R25740 VSS.n849 VSS.n491 0.0103214
R25741 VSS.n845 VSS.n496 0.0103214
R25742 VSS.n836 VSS.n505 0.0103214
R25743 VSS.n589 VSS.n508 0.0103214
R25744 VSS.n807 VSS.n623 0.0103214
R25745 VSS.n802 VSS.n645 0.0103214
R25746 VSS.n657 VSS.n651 0.0103214
R25747 VSS.n806 VSS.n805 0.0103214
R25748 VSS.n656 VSS.n653 0.0103214
R25749 VSS.n986 VSS.n451 0.0103214
R25750 VSS.n464 VSS.n461 0.0103214
R25751 VSS.n973 VSS.n466 0.0103214
R25752 VSS.n947 VSS.n873 0.0103214
R25753 VSS.n8416 VSS.n7199 0.0103214
R25754 VSS.n8411 VSS.n7221 0.0103214
R25755 VSS.n7233 VSS.n7227 0.0103214
R25756 VSS.n8415 VSS.n8414 0.0103214
R25757 VSS.n7232 VSS.n7229 0.0103214
R25758 VSS.n7670 VSS.n7669 0.00956429
R25759 VSS.n7687 VSS.n7670 0.00956429
R25760 VSS.n8262 VSS.n8261 0.00956429
R25761 VSS.n8279 VSS.n8262 0.00956429
R25762 VSS.n8966 VSS.n8815 0.00956429
R25763 VSS.n8861 VSS.n8815 0.00956429
R25764 VSS.n1531 VSS.n1530 0.00956429
R25765 VSS.n1617 VSS.n1531 0.00956429
R25766 VSS.n2104 VSS.n2103 0.00956429
R25767 VSS.n2209 VSS.n2104 0.00956429
R25768 VSS.n3872 VSS.n3871 0.00956429
R25769 VSS.n3889 VSS.n3872 0.00956429
R25770 VSS.n4464 VSS.n4463 0.00956429
R25771 VSS.n4481 VSS.n4464 0.00956429
R25772 VSS.n5056 VSS.n5055 0.00956429
R25773 VSS.n5073 VSS.n5056 0.00956429
R25774 VSS.n5648 VSS.n5647 0.00956429
R25775 VSS.n5665 VSS.n5648 0.00956429
R25776 VSS.n6240 VSS.n6239 0.00956429
R25777 VSS.n6257 VSS.n6240 0.00956429
R25778 VSS.n6832 VSS.n6831 0.00956429
R25779 VSS.n6849 VSS.n6832 0.00956429
R25780 VSS.n2702 VSS.n2701 0.00956429
R25781 VSS.n6953 VSS.n2702 0.00956429
R25782 VSS.n3280 VSS.n3279 0.00956429
R25783 VSS.n3297 VSS.n3280 0.00956429
R25784 VSS.n9240 VSS.n9239 0.00956429
R25785 VSS.n9257 VSS.n9240 0.00956429
R25786 VSS.n694 VSS.n693 0.00956429
R25787 VSS.n772 VSS.n694 0.00956429
R25788 VSS.n7270 VSS.n7269 0.00956429
R25789 VSS.n8381 VSS.n7270 0.00956429
R25790 VSS.n7128 VSS.n7127 0.00942857
R25791 VSS.n8440 VSS.n8439 0.00942857
R25792 VSS.n7178 VSS.n7177 0.00942857
R25793 VSS.n7126 VSS.n7125 0.00942857
R25794 VSS.n7139 VSS.n7068 0.00942857
R25795 VSS.n7082 VSS.n7079 0.00942857
R25796 VSS.n7179 VSS.n7105 0.00942857
R25797 VSS.n903 VSS.n893 0.00942857
R25798 VSS.n992 VSS.n991 0.00942857
R25799 VSS.n872 VSS.n477 0.00942857
R25800 VSS.n7496 VSS.n7495 0.00942857
R25801 VSS.n7568 VSS.n7426 0.00942857
R25802 VSS.n7429 VSS.n7427 0.00942857
R25803 VSS.n1084 VSS.n1074 0.00942857
R25804 VSS.n8513 VSS.n8512 0.00942857
R25805 VSS.n1053 VSS.n1044 0.00942857
R25806 VSS.n1083 VSS.n1082 0.00942857
R25807 VSS.n8503 VSS.n1023 0.00942857
R25808 VSS.n1113 VSS.n1036 0.00942857
R25809 VSS.n1129 VSS.n1042 0.00942857
R25810 VSS.n7661 VSS.n7382 0.00942857
R25811 VSS.n7666 VSS.n7665 0.00942857
R25812 VSS.n7677 VSS.n7675 0.00942857
R25813 VSS.n7721 VSS.n7357 0.00942857
R25814 VSS.n7735 VSS.n7350 0.00942857
R25815 VSS.n7356 VSS.n7351 0.00942857
R25816 VSS.n7494 VSS.n7477 0.00942857
R25817 VSS.n7515 VSS.n7463 0.00942857
R25818 VSS.n7542 VSS.n7541 0.00942857
R25819 VSS.n7428 VSS.n7422 0.00942857
R25820 VSS.n8088 VSS.n8087 0.00942857
R25821 VSS.n8160 VSS.n7840 0.00942857
R25822 VSS.n7843 VSS.n7841 0.00942857
R25823 VSS.n7998 VSS.n7963 0.00942857
R25824 VSS.n7967 VSS.n7966 0.00942857
R25825 VSS.n8060 VSS.n8059 0.00942857
R25826 VSS.n7986 VSS.n7964 0.00942857
R25827 VSS.n8023 VSS.n7946 0.00942857
R25828 VSS.n7931 VSS.n7921 0.00942857
R25829 VSS.n8058 VSS.n7912 0.00942857
R25830 VSS.n8253 VSS.n7796 0.00942857
R25831 VSS.n8258 VSS.n8257 0.00942857
R25832 VSS.n8269 VSS.n8267 0.00942857
R25833 VSS.n8313 VSS.n7771 0.00942857
R25834 VSS.n8327 VSS.n7764 0.00942857
R25835 VSS.n7770 VSS.n7765 0.00942857
R25836 VSS.n8086 VSS.n7891 0.00942857
R25837 VSS.n8107 VSS.n7877 0.00942857
R25838 VSS.n8134 VSS.n8133 0.00942857
R25839 VSS.n7842 VSS.n7836 0.00942857
R25840 VSS.n8559 VSS.n260 0.00942857
R25841 VSS.n264 VSS.n263 0.00942857
R25842 VSS.n8621 VSS.n8620 0.00942857
R25843 VSS.n8707 VSS.n8706 0.00942857
R25844 VSS.n9013 VSS.n9012 0.00942857
R25845 VSS.n8757 VSS.n8756 0.00942857
R25846 VSS.n8705 VSS.n8704 0.00942857
R25847 VSS.n8718 VSS.n8647 0.00942857
R25848 VSS.n8661 VSS.n8658 0.00942857
R25849 VSS.n8758 VSS.n8684 0.00942857
R25850 VSS.n8840 VSS.n8839 0.00942857
R25851 VSS.n8963 VSS.n8818 0.00942857
R25852 VSS.n8866 VSS.n8857 0.00942857
R25853 VSS.n8945 VSS.n8882 0.00942857
R25854 VSS.n8941 VSS.n8886 0.00942857
R25855 VSS.n8940 VSS.n8939 0.00942857
R25856 VSS.n8547 VSS.n261 0.00942857
R25857 VSS.n8584 VSS.n243 0.00942857
R25858 VSS.n228 VSS.n218 0.00942857
R25859 VSS.n8619 VSS.n209 0.00942857
R25860 VSS.n1241 VSS.n1206 0.00942857
R25861 VSS.n1210 VSS.n1209 0.00942857
R25862 VSS.n1303 VSS.n1302 0.00942857
R25863 VSS.n1389 VSS.n1388 0.00942857
R25864 VSS.n1676 VSS.n1675 0.00942857
R25865 VSS.n1439 VSS.n1438 0.00942857
R25866 VSS.n1387 VSS.n1386 0.00942857
R25867 VSS.n1400 VSS.n1329 0.00942857
R25868 VSS.n1343 VSS.n1340 0.00942857
R25869 VSS.n1440 VSS.n1366 0.00942857
R25870 VSS.n1522 VSS.n1513 0.00942857
R25871 VSS.n1527 VSS.n1526 0.00942857
R25872 VSS.n1574 VSS.n1573 0.00942857
R25873 VSS.n1551 VSS.n1543 0.00942857
R25874 VSS.n1595 VSS.n1564 0.00942857
R25875 VSS.n1563 VSS.n1550 0.00942857
R25876 VSS.n1229 VSS.n1207 0.00942857
R25877 VSS.n1266 VSS.n1189 0.00942857
R25878 VSS.n1174 VSS.n1164 0.00942857
R25879 VSS.n1301 VSS.n1155 0.00942857
R25880 VSS.n1814 VSS.n1779 0.00942857
R25881 VSS.n1783 VSS.n1782 0.00942857
R25882 VSS.n1876 VSS.n1875 0.00942857
R25883 VSS.n1962 VSS.n1961 0.00942857
R25884 VSS.n2268 VSS.n2267 0.00942857
R25885 VSS.n2012 VSS.n2011 0.00942857
R25886 VSS.n1960 VSS.n1959 0.00942857
R25887 VSS.n1973 VSS.n1902 0.00942857
R25888 VSS.n1916 VSS.n1913 0.00942857
R25889 VSS.n2013 VSS.n1939 0.00942857
R25890 VSS.n2095 VSS.n2086 0.00942857
R25891 VSS.n2100 VSS.n2099 0.00942857
R25892 VSS.n2134 VSS.n2133 0.00942857
R25893 VSS.n2124 VSS.n2116 0.00942857
R25894 VSS.n2187 VSS.n2125 0.00942857
R25895 VSS.n2162 VSS.n2123 0.00942857
R25896 VSS.n1802 VSS.n1780 0.00942857
R25897 VSS.n1839 VSS.n1762 0.00942857
R25898 VSS.n1747 VSS.n1737 0.00942857
R25899 VSS.n1874 VSS.n1728 0.00942857
R25900 VSS.n3608 VSS.n3573 0.00942857
R25901 VSS.n3577 VSS.n3576 0.00942857
R25902 VSS.n3670 VSS.n3669 0.00942857
R25903 VSS.n3698 VSS.n3697 0.00942857
R25904 VSS.n3770 VSS.n3450 0.00942857
R25905 VSS.n3453 VSS.n3451 0.00942857
R25906 VSS.n3696 VSS.n3501 0.00942857
R25907 VSS.n3717 VSS.n3487 0.00942857
R25908 VSS.n3744 VSS.n3743 0.00942857
R25909 VSS.n3452 VSS.n3446 0.00942857
R25910 VSS.n3863 VSS.n3406 0.00942857
R25911 VSS.n3868 VSS.n3867 0.00942857
R25912 VSS.n3879 VSS.n3877 0.00942857
R25913 VSS.n3923 VSS.n3381 0.00942857
R25914 VSS.n3938 VSS.n3375 0.00942857
R25915 VSS.n3937 VSS.n3377 0.00942857
R25916 VSS.n3596 VSS.n3574 0.00942857
R25917 VSS.n3633 VSS.n3556 0.00942857
R25918 VSS.n3541 VSS.n3531 0.00942857
R25919 VSS.n3668 VSS.n3522 0.00942857
R25920 VSS.n4200 VSS.n4165 0.00942857
R25921 VSS.n4169 VSS.n4168 0.00942857
R25922 VSS.n4262 VSS.n4261 0.00942857
R25923 VSS.n4290 VSS.n4289 0.00942857
R25924 VSS.n4362 VSS.n4042 0.00942857
R25925 VSS.n4045 VSS.n4043 0.00942857
R25926 VSS.n4288 VSS.n4093 0.00942857
R25927 VSS.n4309 VSS.n4079 0.00942857
R25928 VSS.n4336 VSS.n4335 0.00942857
R25929 VSS.n4044 VSS.n4038 0.00942857
R25930 VSS.n4455 VSS.n3998 0.00942857
R25931 VSS.n4460 VSS.n4459 0.00942857
R25932 VSS.n4471 VSS.n4469 0.00942857
R25933 VSS.n4515 VSS.n3973 0.00942857
R25934 VSS.n4530 VSS.n3967 0.00942857
R25935 VSS.n4529 VSS.n3969 0.00942857
R25936 VSS.n4188 VSS.n4166 0.00942857
R25937 VSS.n4225 VSS.n4148 0.00942857
R25938 VSS.n4133 VSS.n4123 0.00942857
R25939 VSS.n4260 VSS.n4114 0.00942857
R25940 VSS.n4792 VSS.n4757 0.00942857
R25941 VSS.n4761 VSS.n4760 0.00942857
R25942 VSS.n4854 VSS.n4853 0.00942857
R25943 VSS.n4882 VSS.n4881 0.00942857
R25944 VSS.n4954 VSS.n4634 0.00942857
R25945 VSS.n4637 VSS.n4635 0.00942857
R25946 VSS.n4880 VSS.n4685 0.00942857
R25947 VSS.n4901 VSS.n4671 0.00942857
R25948 VSS.n4928 VSS.n4927 0.00942857
R25949 VSS.n4636 VSS.n4630 0.00942857
R25950 VSS.n5047 VSS.n4590 0.00942857
R25951 VSS.n5052 VSS.n5051 0.00942857
R25952 VSS.n5063 VSS.n5061 0.00942857
R25953 VSS.n5107 VSS.n4565 0.00942857
R25954 VSS.n5122 VSS.n4559 0.00942857
R25955 VSS.n5121 VSS.n4561 0.00942857
R25956 VSS.n4780 VSS.n4758 0.00942857
R25957 VSS.n4817 VSS.n4740 0.00942857
R25958 VSS.n4725 VSS.n4715 0.00942857
R25959 VSS.n4852 VSS.n4706 0.00942857
R25960 VSS.n5384 VSS.n5349 0.00942857
R25961 VSS.n5353 VSS.n5352 0.00942857
R25962 VSS.n5446 VSS.n5445 0.00942857
R25963 VSS.n5474 VSS.n5473 0.00942857
R25964 VSS.n5546 VSS.n5226 0.00942857
R25965 VSS.n5229 VSS.n5227 0.00942857
R25966 VSS.n5472 VSS.n5277 0.00942857
R25967 VSS.n5493 VSS.n5263 0.00942857
R25968 VSS.n5520 VSS.n5519 0.00942857
R25969 VSS.n5228 VSS.n5222 0.00942857
R25970 VSS.n5639 VSS.n5182 0.00942857
R25971 VSS.n5644 VSS.n5643 0.00942857
R25972 VSS.n5655 VSS.n5653 0.00942857
R25973 VSS.n5699 VSS.n5157 0.00942857
R25974 VSS.n5714 VSS.n5151 0.00942857
R25975 VSS.n5713 VSS.n5153 0.00942857
R25976 VSS.n5372 VSS.n5350 0.00942857
R25977 VSS.n5409 VSS.n5332 0.00942857
R25978 VSS.n5317 VSS.n5307 0.00942857
R25979 VSS.n5444 VSS.n5298 0.00942857
R25980 VSS.n5976 VSS.n5941 0.00942857
R25981 VSS.n5945 VSS.n5944 0.00942857
R25982 VSS.n6038 VSS.n6037 0.00942857
R25983 VSS.n6066 VSS.n6065 0.00942857
R25984 VSS.n6138 VSS.n5818 0.00942857
R25985 VSS.n5821 VSS.n5819 0.00942857
R25986 VSS.n6064 VSS.n5869 0.00942857
R25987 VSS.n6085 VSS.n5855 0.00942857
R25988 VSS.n6112 VSS.n6111 0.00942857
R25989 VSS.n5820 VSS.n5814 0.00942857
R25990 VSS.n6231 VSS.n5774 0.00942857
R25991 VSS.n6236 VSS.n6235 0.00942857
R25992 VSS.n6247 VSS.n6245 0.00942857
R25993 VSS.n6291 VSS.n5749 0.00942857
R25994 VSS.n6306 VSS.n5743 0.00942857
R25995 VSS.n6305 VSS.n5745 0.00942857
R25996 VSS.n5964 VSS.n5942 0.00942857
R25997 VSS.n6001 VSS.n5924 0.00942857
R25998 VSS.n5909 VSS.n5899 0.00942857
R25999 VSS.n6036 VSS.n5890 0.00942857
R26000 VSS.n6568 VSS.n6533 0.00942857
R26001 VSS.n6537 VSS.n6536 0.00942857
R26002 VSS.n6630 VSS.n6629 0.00942857
R26003 VSS.n6658 VSS.n6657 0.00942857
R26004 VSS.n6730 VSS.n6410 0.00942857
R26005 VSS.n6413 VSS.n6411 0.00942857
R26006 VSS.n6656 VSS.n6461 0.00942857
R26007 VSS.n6677 VSS.n6447 0.00942857
R26008 VSS.n6704 VSS.n6703 0.00942857
R26009 VSS.n6412 VSS.n6406 0.00942857
R26010 VSS.n6823 VSS.n6366 0.00942857
R26011 VSS.n6828 VSS.n6827 0.00942857
R26012 VSS.n6839 VSS.n6837 0.00942857
R26013 VSS.n6883 VSS.n6341 0.00942857
R26014 VSS.n6898 VSS.n6335 0.00942857
R26015 VSS.n6897 VSS.n6337 0.00942857
R26016 VSS.n6556 VSS.n6534 0.00942857
R26017 VSS.n6593 VSS.n6516 0.00942857
R26018 VSS.n6501 VSS.n6491 0.00942857
R26019 VSS.n6628 VSS.n6482 0.00942857
R26020 VSS.n2412 VSS.n2377 0.00942857
R26021 VSS.n2381 VSS.n2380 0.00942857
R26022 VSS.n2474 VSS.n2473 0.00942857
R26023 VSS.n2560 VSS.n2559 0.00942857
R26024 VSS.n7012 VSS.n7011 0.00942857
R26025 VSS.n2610 VSS.n2609 0.00942857
R26026 VSS.n2558 VSS.n2557 0.00942857
R26027 VSS.n2571 VSS.n2500 0.00942857
R26028 VSS.n2514 VSS.n2511 0.00942857
R26029 VSS.n2611 VSS.n2537 0.00942857
R26030 VSS.n2693 VSS.n2684 0.00942857
R26031 VSS.n2698 VSS.n2697 0.00942857
R26032 VSS.n2732 VSS.n2731 0.00942857
R26033 VSS.n2722 VSS.n2714 0.00942857
R26034 VSS.n6931 VSS.n2723 0.00942857
R26035 VSS.n2760 VSS.n2721 0.00942857
R26036 VSS.n2400 VSS.n2378 0.00942857
R26037 VSS.n2437 VSS.n2360 0.00942857
R26038 VSS.n2345 VSS.n2335 0.00942857
R26039 VSS.n2472 VSS.n2326 0.00942857
R26040 VSS.n3009 VSS.n2976 0.00942857
R26041 VSS.n2979 VSS.n2978 0.00942857
R26042 VSS.n3079 VSS.n2927 0.00942857
R26043 VSS.n3106 VSS.n3105 0.00942857
R26044 VSS.n3178 VSS.n2857 0.00942857
R26045 VSS.n2860 VSS.n2858 0.00942857
R26046 VSS.n3104 VSS.n2908 0.00942857
R26047 VSS.n3125 VSS.n2894 0.00942857
R26048 VSS.n3152 VSS.n3151 0.00942857
R26049 VSS.n2859 VSS.n2853 0.00942857
R26050 VSS.n3271 VSS.n2813 0.00942857
R26051 VSS.n3276 VSS.n3275 0.00942857
R26052 VSS.n3287 VSS.n3285 0.00942857
R26053 VSS.n3331 VSS.n2788 0.00942857
R26054 VSS.n3346 VSS.n2782 0.00942857
R26055 VSS.n3345 VSS.n2784 0.00942857
R26056 VSS.n2997 VSS.n2977 0.00942857
R26057 VSS.n3023 VSS.n2952 0.00942857
R26058 VSS.n3059 VSS.n3058 0.00942857
R26059 VSS.n3081 VSS.n3080 0.00942857
R26060 VSS.n338 VSS.n330 0.00942857
R26061 VSS.n427 VSS.n426 0.00942857
R26062 VSS.n396 VSS.n395 0.00942857
R26063 VSS.n9066 VSS.n9065 0.00942857
R26064 VSS.n9138 VSS.n124 0.00942857
R26065 VSS.n127 VSS.n125 0.00942857
R26066 VSS.n9064 VSS.n175 0.00942857
R26067 VSS.n9085 VSS.n161 0.00942857
R26068 VSS.n9112 VSS.n9111 0.00942857
R26069 VSS.n126 VSS.n120 0.00942857
R26070 VSS.n9231 VSS.n80 0.00942857
R26071 VSS.n9236 VSS.n9235 0.00942857
R26072 VSS.n9247 VSS.n9245 0.00942857
R26073 VSS.n9291 VSS.n55 0.00942857
R26074 VSS.n9306 VSS.n49 0.00942857
R26075 VSS.n9305 VSS.n51 0.00942857
R26076 VSS.n337 VSS.n336 0.00942857
R26077 VSS.n417 VSS.n290 0.00942857
R26078 VSS.n374 VSS.n303 0.00942857
R26079 VSS.n397 VSS.n308 0.00942857
R26080 VSS.n552 VSS.n482 0.00942857
R26081 VSS.n831 VSS.n830 0.00942857
R26082 VSS.n602 VSS.n601 0.00942857
R26083 VSS.n551 VSS.n483 0.00942857
R26084 VSS.n563 VSS.n489 0.00942857
R26085 VSS.n503 VSS.n500 0.00942857
R26086 VSS.n603 VSS.n526 0.00942857
R26087 VSS.n685 VSS.n676 0.00942857
R26088 VSS.n690 VSS.n689 0.00942857
R26089 VSS.n733 VSS.n732 0.00942857
R26090 VSS.n714 VSS.n706 0.00942857
R26091 VSS.n750 VSS.n726 0.00942857
R26092 VSS.n725 VSS.n713 0.00942857
R26093 VSS.n902 VSS.n901 0.00942857
R26094 VSS.n982 VSS.n456 0.00942857
R26095 VSS.n932 VSS.n469 0.00942857
R26096 VSS.n948 VSS.n475 0.00942857
R26097 VSS.n7261 VSS.n7252 0.00942857
R26098 VSS.n7266 VSS.n7265 0.00942857
R26099 VSS.n7300 VSS.n7299 0.00942857
R26100 VSS.n7290 VSS.n7282 0.00942857
R26101 VSS.n8359 VSS.n7291 0.00942857
R26102 VSS.n7328 VSS.n7289 0.00942857
R26103 VSS.n7104 VSS.n7095 0.00853571
R26104 VSS.n7180 VSS.n7093 0.00853571
R26105 VSS.n7097 VSS.n7094 0.00853571
R26106 VSS.n897 VSS.n896 0.00853571
R26107 VSS.n908 VSS.n907 0.00853571
R26108 VSS.n7573 VSS.n7421 0.00853571
R26109 VSS.n1078 VSS.n1077 0.00853571
R26110 VSS.n1089 VSS.n1088 0.00853571
R26111 VSS.n8519 VSS.n8518 0.00853571
R26112 VSS.n1076 VSS.n1075 0.00853571
R26113 VSS.n1086 VSS.n1018 0.00853571
R26114 VSS.n7651 VSS.n7650 0.00853571
R26115 VSS.n7690 VSS.n7377 0.00853571
R26116 VSS.n7703 VSS.n7702 0.00853571
R26117 VSS.n7615 VSS.n7410 0.00853571
R26118 VSS.n7622 VSS.n7407 0.00853571
R26119 VSS.n7652 VSS.n7385 0.00853571
R26120 VSS.n7657 VSS.n7656 0.00853571
R26121 VSS.n7704 VSS.n7367 0.00853571
R26122 VSS.n7704 VSS.n7368 0.00853571
R26123 VSS.n7731 VSS.n7353 0.00853571
R26124 VSS.n7727 VSS.n7353 0.00853571
R26125 VSS.n7749 VSS.n7340 0.00853571
R26126 VSS.n7575 VSS.n7574 0.00853571
R26127 VSS.n7611 VSS.n7412 0.00853571
R26128 VSS.n8165 VSS.n7835 0.00853571
R26129 VSS.n7990 VSS.n7989 0.00853571
R26130 VSS.n8013 VSS.n7952 0.00853571
R26131 VSS.n7982 VSS.n7970 0.00853571
R26132 VSS.n7988 VSS.n7971 0.00853571
R26133 VSS.n7953 VSS.n7951 0.00853571
R26134 VSS.n8243 VSS.n8242 0.00853571
R26135 VSS.n8282 VSS.n7791 0.00853571
R26136 VSS.n8295 VSS.n8294 0.00853571
R26137 VSS.n8207 VSS.n7824 0.00853571
R26138 VSS.n8214 VSS.n7821 0.00853571
R26139 VSS.n8244 VSS.n7799 0.00853571
R26140 VSS.n8249 VSS.n8248 0.00853571
R26141 VSS.n8296 VSS.n7781 0.00853571
R26142 VSS.n8296 VSS.n7782 0.00853571
R26143 VSS.n8323 VSS.n7767 0.00853571
R26144 VSS.n8319 VSS.n7767 0.00853571
R26145 VSS.n8341 VSS.n7754 0.00853571
R26146 VSS.n8167 VSS.n8166 0.00853571
R26147 VSS.n8203 VSS.n7826 0.00853571
R26148 VSS.n8551 VSS.n8550 0.00853571
R26149 VSS.n8574 VSS.n249 0.00853571
R26150 VSS.n8683 VSS.n8674 0.00853571
R26151 VSS.n8759 VSS.n8672 0.00853571
R26152 VSS.n8676 VSS.n8673 0.00853571
R26153 VSS.n8971 VSS.n8805 0.00853571
R26154 VSS.n8865 VSS.n8864 0.00853571
R26155 VSS.n8951 VSS.n8852 0.00853571
R26156 VSS.n8793 VSS.n8789 0.00853571
R26157 VSS.n8798 VSS.n8782 0.00853571
R26158 VSS.n8812 VSS.n8811 0.00853571
R26159 VSS.n8968 VSS.n8809 0.00853571
R26160 VSS.n8950 VSS.n8853 0.00853571
R26161 VSS.n8950 VSS.n8854 0.00853571
R26162 VSS.n8934 VSS.n8890 0.00853571
R26163 VSS.n8894 VSS.n8890 0.00853571
R26164 VSS.n8930 VSS.n8929 0.00853571
R26165 VSS.n8543 VSS.n267 0.00853571
R26166 VSS.n8549 VSS.n268 0.00853571
R26167 VSS.n250 VSS.n248 0.00853571
R26168 VSS.n1233 VSS.n1232 0.00853571
R26169 VSS.n1256 VSS.n1195 0.00853571
R26170 VSS.n1365 VSS.n1356 0.00853571
R26171 VSS.n1441 VSS.n1354 0.00853571
R26172 VSS.n1358 VSS.n1355 0.00853571
R26173 VSS.n1632 VSS.n1631 0.00853571
R26174 VSS.n1620 VSS.n1508 0.00853571
R26175 VSS.n1608 VSS.n1536 0.00853571
R26176 VSS.n1474 VSS.n1470 0.00853571
R26177 VSS.n1479 VSS.n1464 0.00853571
R26178 VSS.n1633 VSS.n1491 0.00853571
R26179 VSS.n1518 VSS.n1517 0.00853571
R26180 VSS.n1546 VSS.n1540 0.00853571
R26181 VSS.n1607 VSS.n1540 0.00853571
R26182 VSS.n1555 VSS.n1553 0.00853571
R26183 VSS.n1556 VSS.n1555 0.00853571
R26184 VSS.n9349 VSS.n2 0.00853571
R26185 VSS.n1225 VSS.n1213 0.00853571
R26186 VSS.n1231 VSS.n1214 0.00853571
R26187 VSS.n1196 VSS.n1194 0.00853571
R26188 VSS.n1806 VSS.n1805 0.00853571
R26189 VSS.n1829 VSS.n1768 0.00853571
R26190 VSS.n1938 VSS.n1929 0.00853571
R26191 VSS.n2014 VSS.n1927 0.00853571
R26192 VSS.n1931 VSS.n1928 0.00853571
R26193 VSS.n2224 VSS.n2223 0.00853571
R26194 VSS.n2212 VSS.n2081 0.00853571
R26195 VSS.n2200 VSS.n2109 0.00853571
R26196 VSS.n2047 VSS.n2043 0.00853571
R26197 VSS.n2052 VSS.n2037 0.00853571
R26198 VSS.n2225 VSS.n2064 0.00853571
R26199 VSS.n2091 VSS.n2090 0.00853571
R26200 VSS.n2119 VSS.n2113 0.00853571
R26201 VSS.n2199 VSS.n2113 0.00853571
R26202 VSS.n2170 VSS.n2168 0.00853571
R26203 VSS.n2170 VSS.n2169 0.00853571
R26204 VSS.n2175 VSS.n2155 0.00853571
R26205 VSS.n1798 VSS.n1786 0.00853571
R26206 VSS.n1804 VSS.n1787 0.00853571
R26207 VSS.n1769 VSS.n1767 0.00853571
R26208 VSS.n3600 VSS.n3599 0.00853571
R26209 VSS.n3623 VSS.n3562 0.00853571
R26210 VSS.n3775 VSS.n3445 0.00853571
R26211 VSS.n3777 VSS.n3776 0.00853571
R26212 VSS.n3813 VSS.n3436 0.00853571
R26213 VSS.n3853 VSS.n3852 0.00853571
R26214 VSS.n3892 VSS.n3401 0.00853571
R26215 VSS.n3905 VSS.n3904 0.00853571
R26216 VSS.n3817 VSS.n3434 0.00853571
R26217 VSS.n3824 VSS.n3431 0.00853571
R26218 VSS.n3854 VSS.n3409 0.00853571
R26219 VSS.n3859 VSS.n3858 0.00853571
R26220 VSS.n3906 VSS.n3391 0.00853571
R26221 VSS.n3906 VSS.n3392 0.00853571
R26222 VSS.n3929 VSS.n3378 0.00853571
R26223 VSS.n3930 VSS.n3929 0.00853571
R26224 VSS.n3952 VSS.n3365 0.00853571
R26225 VSS.n3592 VSS.n3580 0.00853571
R26226 VSS.n3598 VSS.n3581 0.00853571
R26227 VSS.n3563 VSS.n3561 0.00853571
R26228 VSS.n4192 VSS.n4191 0.00853571
R26229 VSS.n4215 VSS.n4154 0.00853571
R26230 VSS.n4367 VSS.n4037 0.00853571
R26231 VSS.n4369 VSS.n4368 0.00853571
R26232 VSS.n4405 VSS.n4028 0.00853571
R26233 VSS.n4445 VSS.n4444 0.00853571
R26234 VSS.n4484 VSS.n3993 0.00853571
R26235 VSS.n4497 VSS.n4496 0.00853571
R26236 VSS.n4409 VSS.n4026 0.00853571
R26237 VSS.n4416 VSS.n4023 0.00853571
R26238 VSS.n4446 VSS.n4001 0.00853571
R26239 VSS.n4451 VSS.n4450 0.00853571
R26240 VSS.n4498 VSS.n3983 0.00853571
R26241 VSS.n4498 VSS.n3984 0.00853571
R26242 VSS.n4521 VSS.n3970 0.00853571
R26243 VSS.n4522 VSS.n4521 0.00853571
R26244 VSS.n4544 VSS.n3957 0.00853571
R26245 VSS.n4184 VSS.n4172 0.00853571
R26246 VSS.n4190 VSS.n4173 0.00853571
R26247 VSS.n4155 VSS.n4153 0.00853571
R26248 VSS.n4784 VSS.n4783 0.00853571
R26249 VSS.n4807 VSS.n4746 0.00853571
R26250 VSS.n4959 VSS.n4629 0.00853571
R26251 VSS.n4961 VSS.n4960 0.00853571
R26252 VSS.n4997 VSS.n4620 0.00853571
R26253 VSS.n5037 VSS.n5036 0.00853571
R26254 VSS.n5076 VSS.n4585 0.00853571
R26255 VSS.n5089 VSS.n5088 0.00853571
R26256 VSS.n5001 VSS.n4618 0.00853571
R26257 VSS.n5008 VSS.n4615 0.00853571
R26258 VSS.n5038 VSS.n4593 0.00853571
R26259 VSS.n5043 VSS.n5042 0.00853571
R26260 VSS.n5090 VSS.n4575 0.00853571
R26261 VSS.n5090 VSS.n4576 0.00853571
R26262 VSS.n5113 VSS.n4562 0.00853571
R26263 VSS.n5114 VSS.n5113 0.00853571
R26264 VSS.n5136 VSS.n4549 0.00853571
R26265 VSS.n4776 VSS.n4764 0.00853571
R26266 VSS.n4782 VSS.n4765 0.00853571
R26267 VSS.n4747 VSS.n4745 0.00853571
R26268 VSS.n5376 VSS.n5375 0.00853571
R26269 VSS.n5399 VSS.n5338 0.00853571
R26270 VSS.n5551 VSS.n5221 0.00853571
R26271 VSS.n5553 VSS.n5552 0.00853571
R26272 VSS.n5589 VSS.n5212 0.00853571
R26273 VSS.n5629 VSS.n5628 0.00853571
R26274 VSS.n5668 VSS.n5177 0.00853571
R26275 VSS.n5681 VSS.n5680 0.00853571
R26276 VSS.n5593 VSS.n5210 0.00853571
R26277 VSS.n5600 VSS.n5207 0.00853571
R26278 VSS.n5630 VSS.n5185 0.00853571
R26279 VSS.n5635 VSS.n5634 0.00853571
R26280 VSS.n5682 VSS.n5167 0.00853571
R26281 VSS.n5682 VSS.n5168 0.00853571
R26282 VSS.n5705 VSS.n5154 0.00853571
R26283 VSS.n5706 VSS.n5705 0.00853571
R26284 VSS.n5728 VSS.n5141 0.00853571
R26285 VSS.n5368 VSS.n5356 0.00853571
R26286 VSS.n5374 VSS.n5357 0.00853571
R26287 VSS.n5339 VSS.n5337 0.00853571
R26288 VSS.n5968 VSS.n5967 0.00853571
R26289 VSS.n5991 VSS.n5930 0.00853571
R26290 VSS.n6143 VSS.n5813 0.00853571
R26291 VSS.n6145 VSS.n6144 0.00853571
R26292 VSS.n6181 VSS.n5804 0.00853571
R26293 VSS.n6221 VSS.n6220 0.00853571
R26294 VSS.n6260 VSS.n5769 0.00853571
R26295 VSS.n6273 VSS.n6272 0.00853571
R26296 VSS.n6185 VSS.n5802 0.00853571
R26297 VSS.n6192 VSS.n5799 0.00853571
R26298 VSS.n6222 VSS.n5777 0.00853571
R26299 VSS.n6227 VSS.n6226 0.00853571
R26300 VSS.n6274 VSS.n5759 0.00853571
R26301 VSS.n6274 VSS.n5760 0.00853571
R26302 VSS.n6297 VSS.n5746 0.00853571
R26303 VSS.n6298 VSS.n6297 0.00853571
R26304 VSS.n6320 VSS.n5733 0.00853571
R26305 VSS.n5960 VSS.n5948 0.00853571
R26306 VSS.n5966 VSS.n5949 0.00853571
R26307 VSS.n5931 VSS.n5929 0.00853571
R26308 VSS.n6560 VSS.n6559 0.00853571
R26309 VSS.n6583 VSS.n6522 0.00853571
R26310 VSS.n6735 VSS.n6405 0.00853571
R26311 VSS.n6737 VSS.n6736 0.00853571
R26312 VSS.n6773 VSS.n6396 0.00853571
R26313 VSS.n6813 VSS.n6812 0.00853571
R26314 VSS.n6852 VSS.n6361 0.00853571
R26315 VSS.n6865 VSS.n6864 0.00853571
R26316 VSS.n6777 VSS.n6394 0.00853571
R26317 VSS.n6784 VSS.n6391 0.00853571
R26318 VSS.n6814 VSS.n6369 0.00853571
R26319 VSS.n6819 VSS.n6818 0.00853571
R26320 VSS.n6866 VSS.n6351 0.00853571
R26321 VSS.n6866 VSS.n6352 0.00853571
R26322 VSS.n6889 VSS.n6338 0.00853571
R26323 VSS.n6890 VSS.n6889 0.00853571
R26324 VSS.n6912 VSS.n6325 0.00853571
R26325 VSS.n6552 VSS.n6540 0.00853571
R26326 VSS.n6558 VSS.n6541 0.00853571
R26327 VSS.n6523 VSS.n6521 0.00853571
R26328 VSS.n2404 VSS.n2403 0.00853571
R26329 VSS.n2427 VSS.n2366 0.00853571
R26330 VSS.n2536 VSS.n2527 0.00853571
R26331 VSS.n2612 VSS.n2525 0.00853571
R26332 VSS.n2529 VSS.n2526 0.00853571
R26333 VSS.n6968 VSS.n6967 0.00853571
R26334 VSS.n6956 VSS.n2679 0.00853571
R26335 VSS.n6944 VSS.n2707 0.00853571
R26336 VSS.n2645 VSS.n2641 0.00853571
R26337 VSS.n2650 VSS.n2635 0.00853571
R26338 VSS.n6969 VSS.n2662 0.00853571
R26339 VSS.n2689 VSS.n2688 0.00853571
R26340 VSS.n2717 VSS.n2711 0.00853571
R26341 VSS.n6943 VSS.n2711 0.00853571
R26342 VSS.n2768 VSS.n2766 0.00853571
R26343 VSS.n2768 VSS.n2767 0.00853571
R26344 VSS.n6919 VSS.n2753 0.00853571
R26345 VSS.n2396 VSS.n2384 0.00853571
R26346 VSS.n2402 VSS.n2385 0.00853571
R26347 VSS.n2367 VSS.n2365 0.00853571
R26348 VSS.n3001 VSS.n3000 0.00853571
R26349 VSS.n3019 VSS.n3018 0.00853571
R26350 VSS.n3183 VSS.n2852 0.00853571
R26351 VSS.n3185 VSS.n3184 0.00853571
R26352 VSS.n3221 VSS.n2843 0.00853571
R26353 VSS.n3261 VSS.n3260 0.00853571
R26354 VSS.n3300 VSS.n2808 0.00853571
R26355 VSS.n3313 VSS.n3312 0.00853571
R26356 VSS.n3225 VSS.n2841 0.00853571
R26357 VSS.n3232 VSS.n2838 0.00853571
R26358 VSS.n3262 VSS.n2816 0.00853571
R26359 VSS.n3267 VSS.n3266 0.00853571
R26360 VSS.n3314 VSS.n2798 0.00853571
R26361 VSS.n3314 VSS.n2799 0.00853571
R26362 VSS.n3337 VSS.n2785 0.00853571
R26363 VSS.n3338 VSS.n3337 0.00853571
R26364 VSS.n3360 VSS.n2772 0.00853571
R26365 VSS.n2993 VSS.n2982 0.00853571
R26366 VSS.n2999 VSS.n2983 0.00853571
R26367 VSS.n3028 VSS.n2966 0.00853571
R26368 VSS.n333 VSS.n332 0.00853571
R26369 VSS.n351 VSS.n350 0.00853571
R26370 VSS.n9143 VSS.n119 0.00853571
R26371 VSS.n9145 VSS.n9144 0.00853571
R26372 VSS.n9181 VSS.n110 0.00853571
R26373 VSS.n9221 VSS.n9220 0.00853571
R26374 VSS.n9260 VSS.n75 0.00853571
R26375 VSS.n9273 VSS.n9272 0.00853571
R26376 VSS.n9185 VSS.n108 0.00853571
R26377 VSS.n9192 VSS.n105 0.00853571
R26378 VSS.n9222 VSS.n83 0.00853571
R26379 VSS.n9227 VSS.n9226 0.00853571
R26380 VSS.n9274 VSS.n65 0.00853571
R26381 VSS.n9274 VSS.n66 0.00853571
R26382 VSS.n9297 VSS.n52 0.00853571
R26383 VSS.n9298 VSS.n9297 0.00853571
R26384 VSS.n9320 VSS.n39 0.00853571
R26385 VSS.n433 VSS.n432 0.00853571
R26386 VSS.n334 VSS.n331 0.00853571
R26387 VSS.n352 VSS.n285 0.00853571
R26388 VSS.n525 VSS.n516 0.00853571
R26389 VSS.n604 VSS.n514 0.00853571
R26390 VSS.n518 VSS.n515 0.00853571
R26391 VSS.n787 VSS.n786 0.00853571
R26392 VSS.n775 VSS.n671 0.00853571
R26393 VSS.n763 VSS.n699 0.00853571
R26394 VSS.n637 VSS.n633 0.00853571
R26395 VSS.n642 VSS.n627 0.00853571
R26396 VSS.n788 VSS.n654 0.00853571
R26397 VSS.n681 VSS.n680 0.00853571
R26398 VSS.n709 VSS.n703 0.00853571
R26399 VSS.n762 VSS.n703 0.00853571
R26400 VSS.n719 VSS.n718 0.00853571
R26401 VSS.n718 VSS.n716 0.00853571
R26402 VSS.n9326 VSS.n35 0.00853571
R26403 VSS.n998 VSS.n997 0.00853571
R26404 VSS.n895 VSS.n894 0.00853571
R26405 VSS.n905 VSS.n451 0.00853571
R26406 VSS.n8396 VSS.n8395 0.00853571
R26407 VSS.n8384 VSS.n7247 0.00853571
R26408 VSS.n8372 VSS.n7275 0.00853571
R26409 VSS.n7213 VSS.n7209 0.00853571
R26410 VSS.n7218 VSS.n7203 0.00853571
R26411 VSS.n8397 VSS.n7230 0.00853571
R26412 VSS.n7257 VSS.n7256 0.00853571
R26413 VSS.n7285 VSS.n7279 0.00853571
R26414 VSS.n8371 VSS.n7279 0.00853571
R26415 VSS.n7336 VSS.n7334 0.00853571
R26416 VSS.n7336 VSS.n7335 0.00853571
R26417 VSS.n8347 VSS.n7321 0.00853571
R26418 VSS.n8517 VSS.n1009 0.00822143
R26419 VSS.n8509 VSS.n1011 0.00822143
R26420 VSS.n8492 VSS.n1035 0.00822143
R26421 VSS.n7486 VSS.n1041 0.00822143
R26422 VSS.n7487 VSS.n7475 0.00822143
R26423 VSS.n7517 VSS.n7461 0.00822143
R26424 VSS.n7548 VSS.n7423 0.00822143
R26425 VSS.n7612 VSS.n7411 0.00822143
R26426 VSS.n7981 VSS.n7969 0.00822143
R26427 VSS.n8016 VSS.n7949 0.00822143
R26428 VSS.n8049 VSS.n7918 0.00822143
R26429 VSS.n8078 VSS.n7900 0.00822143
R26430 VSS.n8079 VSS.n7889 0.00822143
R26431 VSS.n8109 VSS.n7875 0.00822143
R26432 VSS.n8140 VSS.n7837 0.00822143
R26433 VSS.n8204 VSS.n7825 0.00822143
R26434 VSS.n8542 VSS.n266 0.00822143
R26435 VSS.n8577 VSS.n246 0.00822143
R26436 VSS.n8610 VSS.n215 0.00822143
R26437 VSS.n8639 VSS.n197 0.00822143
R26438 VSS.n9041 VSS.n8640 0.00822143
R26439 VSS.n9033 VSS.n8642 0.00822143
R26440 VSS.n9016 VSS.n8665 0.00822143
R26441 VSS.n8790 VSS.n8671 0.00822143
R26442 VSS.n1224 VSS.n1212 0.00822143
R26443 VSS.n1259 VSS.n1192 0.00822143
R26444 VSS.n1292 VSS.n1161 0.00822143
R26445 VSS.n1321 VSS.n1143 0.00822143
R26446 VSS.n1704 VSS.n1322 0.00822143
R26447 VSS.n1696 VSS.n1324 0.00822143
R26448 VSS.n1679 VSS.n1347 0.00822143
R26449 VSS.n1471 VSS.n1353 0.00822143
R26450 VSS.n1797 VSS.n1785 0.00822143
R26451 VSS.n1832 VSS.n1765 0.00822143
R26452 VSS.n1865 VSS.n1734 0.00822143
R26453 VSS.n1894 VSS.n1716 0.00822143
R26454 VSS.n2296 VSS.n1895 0.00822143
R26455 VSS.n2288 VSS.n1897 0.00822143
R26456 VSS.n2271 VSS.n1920 0.00822143
R26457 VSS.n2044 VSS.n1926 0.00822143
R26458 VSS.n3591 VSS.n3579 0.00822143
R26459 VSS.n3626 VSS.n3559 0.00822143
R26460 VSS.n3659 VSS.n3528 0.00822143
R26461 VSS.n3688 VSS.n3510 0.00822143
R26462 VSS.n3689 VSS.n3499 0.00822143
R26463 VSS.n3719 VSS.n3485 0.00822143
R26464 VSS.n3750 VSS.n3447 0.00822143
R26465 VSS.n3814 VSS.n3435 0.00822143
R26466 VSS.n4183 VSS.n4171 0.00822143
R26467 VSS.n4218 VSS.n4151 0.00822143
R26468 VSS.n4251 VSS.n4120 0.00822143
R26469 VSS.n4280 VSS.n4102 0.00822143
R26470 VSS.n4281 VSS.n4091 0.00822143
R26471 VSS.n4311 VSS.n4077 0.00822143
R26472 VSS.n4342 VSS.n4039 0.00822143
R26473 VSS.n4406 VSS.n4027 0.00822143
R26474 VSS.n4775 VSS.n4763 0.00822143
R26475 VSS.n4810 VSS.n4743 0.00822143
R26476 VSS.n4843 VSS.n4712 0.00822143
R26477 VSS.n4872 VSS.n4694 0.00822143
R26478 VSS.n4873 VSS.n4683 0.00822143
R26479 VSS.n4903 VSS.n4669 0.00822143
R26480 VSS.n4934 VSS.n4631 0.00822143
R26481 VSS.n4998 VSS.n4619 0.00822143
R26482 VSS.n5367 VSS.n5355 0.00822143
R26483 VSS.n5402 VSS.n5335 0.00822143
R26484 VSS.n5435 VSS.n5304 0.00822143
R26485 VSS.n5464 VSS.n5286 0.00822143
R26486 VSS.n5465 VSS.n5275 0.00822143
R26487 VSS.n5495 VSS.n5261 0.00822143
R26488 VSS.n5526 VSS.n5223 0.00822143
R26489 VSS.n5590 VSS.n5211 0.00822143
R26490 VSS.n5959 VSS.n5947 0.00822143
R26491 VSS.n5994 VSS.n5927 0.00822143
R26492 VSS.n6027 VSS.n5896 0.00822143
R26493 VSS.n6056 VSS.n5878 0.00822143
R26494 VSS.n6057 VSS.n5867 0.00822143
R26495 VSS.n6087 VSS.n5853 0.00822143
R26496 VSS.n6118 VSS.n5815 0.00822143
R26497 VSS.n6182 VSS.n5803 0.00822143
R26498 VSS.n6551 VSS.n6539 0.00822143
R26499 VSS.n6586 VSS.n6519 0.00822143
R26500 VSS.n6619 VSS.n6488 0.00822143
R26501 VSS.n6648 VSS.n6470 0.00822143
R26502 VSS.n6649 VSS.n6459 0.00822143
R26503 VSS.n6679 VSS.n6445 0.00822143
R26504 VSS.n6710 VSS.n6407 0.00822143
R26505 VSS.n6774 VSS.n6395 0.00822143
R26506 VSS.n2395 VSS.n2383 0.00822143
R26507 VSS.n2430 VSS.n2363 0.00822143
R26508 VSS.n2463 VSS.n2332 0.00822143
R26509 VSS.n2492 VSS.n2314 0.00822143
R26510 VSS.n7040 VSS.n2493 0.00822143
R26511 VSS.n7032 VSS.n2495 0.00822143
R26512 VSS.n7015 VSS.n2518 0.00822143
R26513 VSS.n2642 VSS.n2524 0.00822143
R26514 VSS.n2992 VSS.n2981 0.00822143
R26515 VSS.n3022 VSS.n2969 0.00822143
R26516 VSS.n3053 VSS.n2929 0.00822143
R26517 VSS.n3096 VSS.n2917 0.00822143
R26518 VSS.n3097 VSS.n2906 0.00822143
R26519 VSS.n3127 VSS.n2892 0.00822143
R26520 VSS.n3158 VSS.n2854 0.00822143
R26521 VSS.n3222 VSS.n2842 0.00822143
R26522 VSS.n431 VSS.n276 0.00822143
R26523 VSS.n423 VSS.n278 0.00822143
R26524 VSS.n406 VSS.n302 0.00822143
R26525 VSS.n9056 VSS.n177 0.00822143
R26526 VSS.n9057 VSS.n173 0.00822143
R26527 VSS.n9087 VSS.n159 0.00822143
R26528 VSS.n9118 VSS.n121 0.00822143
R26529 VSS.n9182 VSS.n109 0.00822143
R26530 VSS.n996 VSS.n442 0.00822143
R26531 VSS.n988 VSS.n444 0.00822143
R26532 VSS.n971 VSS.n468 0.00822143
R26533 VSS.n864 VSS.n474 0.00822143
R26534 VSS.n863 VSS.n479 0.00822143
R26535 VSS.n851 VSS.n484 0.00822143
R26536 VSS.n834 VSS.n507 0.00822143
R26537 VSS.n634 VSS.n513 0.00822143
R26538 VSS.n8468 VSS.n7061 0.00822143
R26539 VSS.n8460 VSS.n7063 0.00822143
R26540 VSS.n8443 VSS.n7086 0.00822143
R26541 VSS.n7210 VSS.n7092 0.00822143
R26542 VSS.n7141 VSS.n7140 0.00764286
R26543 VSS.n7164 VSS.n7163 0.00764286
R26544 VSS.n8470 VSS.n8469 0.00764286
R26545 VSS.n8461 VSS.n7068 0.00764286
R26546 VSS.n7138 VSS.n7070 0.00764286
R26547 VSS.n7075 VSS.n7074 0.00764286
R26548 VSS.n7083 VSS.n7082 0.00764286
R26549 VSS.n7166 VSS.n7084 0.00764286
R26550 VSS.n934 VSS.n931 0.00764286
R26551 VSS.n7513 VSS.n7465 0.00764286
R26552 VSS.n7551 VSS.n7437 0.00764286
R26553 VSS.n1115 VSS.n1112 0.00764286
R26554 VSS.n1023 VSS.n1022 0.00764286
R26555 VSS.n1032 VSS.n1031 0.00764286
R26556 VSS.n1114 VSS.n1113 0.00764286
R26557 VSS.n8491 VSS.n1036 0.00764286
R26558 VSS.n1046 VSS.n1043 0.00764286
R26559 VSS.n7621 VSS.n7620 0.00764286
R26560 VSS.n7619 VSS.n7402 0.00764286
R26561 VSS.n7651 VSS.n7388 0.00764286
R26562 VSS.n7703 VSS.n7369 0.00764286
R26563 VSS.n7735 VSS.n7734 0.00764286
R26564 VSS.n7734 VSS.n7352 0.00764286
R26565 VSS.n7616 VSS.n7615 0.00764286
R26566 VSS.n7616 VSS.n7407 0.00764286
R26567 VSS.n7622 VSS.n7408 0.00764286
R26568 VSS.n7618 VSS.n7404 0.00764286
R26569 VSS.n7637 VSS.n7636 0.00764286
R26570 VSS.n7652 VSS.n7387 0.00764286
R26571 VSS.n7674 VSS.n7673 0.00764286
R26572 VSS.n7710 VSS.n7365 0.00764286
R26573 VSS.n7733 VSS.n7351 0.00764286
R26574 VSS.n7733 VSS.n7732 0.00764286
R26575 VSS.n7488 VSS.n7476 0.00764286
R26576 VSS.n7516 VSS.n7515 0.00764286
R26577 VSS.n7523 VSS.n7458 0.00764286
R26578 VSS.n7519 VSS.n7518 0.00764286
R26579 VSS.n7541 VSS.n7444 0.00764286
R26580 VSS.n7555 VSS.n7438 0.00764286
R26581 VSS.n8105 VSS.n7879 0.00764286
R26582 VSS.n8143 VSS.n7851 0.00764286
R26583 VSS.n7932 VSS.n7926 0.00764286
R26584 VSS.n8019 VSS.n7946 0.00764286
R26585 VSS.n8027 VSS.n8026 0.00764286
R26586 VSS.n7931 VSS.n7930 0.00764286
R26587 VSS.n8050 VSS.n7921 0.00764286
R26588 VSS.n8077 VSS.n7901 0.00764286
R26589 VSS.n8213 VSS.n8212 0.00764286
R26590 VSS.n8211 VSS.n7816 0.00764286
R26591 VSS.n8243 VSS.n7802 0.00764286
R26592 VSS.n8295 VSS.n7783 0.00764286
R26593 VSS.n8327 VSS.n8326 0.00764286
R26594 VSS.n8326 VSS.n7766 0.00764286
R26595 VSS.n8208 VSS.n8207 0.00764286
R26596 VSS.n8208 VSS.n7821 0.00764286
R26597 VSS.n8214 VSS.n7822 0.00764286
R26598 VSS.n8210 VSS.n7818 0.00764286
R26599 VSS.n8229 VSS.n8228 0.00764286
R26600 VSS.n8244 VSS.n7801 0.00764286
R26601 VSS.n8266 VSS.n8265 0.00764286
R26602 VSS.n8302 VSS.n7779 0.00764286
R26603 VSS.n8325 VSS.n7765 0.00764286
R26604 VSS.n8325 VSS.n8324 0.00764286
R26605 VSS.n8080 VSS.n7890 0.00764286
R26606 VSS.n8108 VSS.n8107 0.00764286
R26607 VSS.n8115 VSS.n7872 0.00764286
R26608 VSS.n8111 VSS.n8110 0.00764286
R26609 VSS.n8133 VSS.n7858 0.00764286
R26610 VSS.n8147 VSS.n7852 0.00764286
R26611 VSS.n229 VSS.n223 0.00764286
R26612 VSS.n8720 VSS.n8719 0.00764286
R26613 VSS.n8743 VSS.n8742 0.00764286
R26614 VSS.n9043 VSS.n9042 0.00764286
R26615 VSS.n9034 VSS.n8647 0.00764286
R26616 VSS.n8717 VSS.n8649 0.00764286
R26617 VSS.n8654 VSS.n8653 0.00764286
R26618 VSS.n8662 VSS.n8661 0.00764286
R26619 VSS.n8745 VSS.n8663 0.00764286
R26620 VSS.n8797 VSS.n8796 0.00764286
R26621 VSS.n8989 VSS.n8777 0.00764286
R26622 VSS.n8975 VSS.n8805 0.00764286
R26623 VSS.n8952 VSS.n8951 0.00764286
R26624 VSS.n8937 VSS.n8886 0.00764286
R26625 VSS.n8937 VSS.n8936 0.00764286
R26626 VSS.n8794 VSS.n8793 0.00764286
R26627 VSS.n8794 VSS.n8782 0.00764286
R26628 VSS.n8798 VSS.n8784 0.00764286
R26629 VSS.n8783 VSS.n8778 0.00764286
R26630 VSS.n8978 VSS.n8977 0.00764286
R26631 VSS.n8811 VSS.n8804 0.00764286
R26632 VSS.n8875 VSS.n8874 0.00764286
R26633 VSS.n8908 VSS.n8907 0.00764286
R26634 VSS.n8939 VSS.n8938 0.00764286
R26635 VSS.n8938 VSS.n8888 0.00764286
R26636 VSS.n8580 VSS.n243 0.00764286
R26637 VSS.n8588 VSS.n8587 0.00764286
R26638 VSS.n228 VSS.n227 0.00764286
R26639 VSS.n8611 VSS.n218 0.00764286
R26640 VSS.n8638 VSS.n198 0.00764286
R26641 VSS.n1175 VSS.n1169 0.00764286
R26642 VSS.n1402 VSS.n1401 0.00764286
R26643 VSS.n1425 VSS.n1424 0.00764286
R26644 VSS.n1706 VSS.n1705 0.00764286
R26645 VSS.n1697 VSS.n1329 0.00764286
R26646 VSS.n1399 VSS.n1331 0.00764286
R26647 VSS.n1336 VSS.n1335 0.00764286
R26648 VSS.n1344 VSS.n1343 0.00764286
R26649 VSS.n1427 VSS.n1345 0.00764286
R26650 VSS.n1478 VSS.n1477 0.00764286
R26651 VSS.n1652 VSS.n1459 0.00764286
R26652 VSS.n1632 VSS.n1489 0.00764286
R26653 VSS.n1612 VSS.n1536 0.00764286
R26654 VSS.n1564 VSS.n1552 0.00764286
R26655 VSS.n1560 VSS.n1552 0.00764286
R26656 VSS.n1475 VSS.n1474 0.00764286
R26657 VSS.n1475 VSS.n1464 0.00764286
R26658 VSS.n1479 VSS.n1465 0.00764286
R26659 VSS.n1651 VSS.n1461 0.00764286
R26660 VSS.n1635 VSS.n1490 0.00764286
R26661 VSS.n1634 VSS.n1633 0.00764286
R26662 VSS.n1545 VSS.n1534 0.00764286
R26663 VSS.n1606 VSS.n1605 0.00764286
R26664 VSS.n1563 VSS.n1562 0.00764286
R26665 VSS.n1562 VSS.n1561 0.00764286
R26666 VSS.n1262 VSS.n1189 0.00764286
R26667 VSS.n1270 VSS.n1269 0.00764286
R26668 VSS.n1174 VSS.n1173 0.00764286
R26669 VSS.n1293 VSS.n1164 0.00764286
R26670 VSS.n1320 VSS.n1144 0.00764286
R26671 VSS.n1748 VSS.n1742 0.00764286
R26672 VSS.n1975 VSS.n1974 0.00764286
R26673 VSS.n1998 VSS.n1997 0.00764286
R26674 VSS.n2298 VSS.n2297 0.00764286
R26675 VSS.n2289 VSS.n1902 0.00764286
R26676 VSS.n1972 VSS.n1904 0.00764286
R26677 VSS.n1909 VSS.n1908 0.00764286
R26678 VSS.n1917 VSS.n1916 0.00764286
R26679 VSS.n2000 VSS.n1918 0.00764286
R26680 VSS.n2051 VSS.n2050 0.00764286
R26681 VSS.n2244 VSS.n2032 0.00764286
R26682 VSS.n2224 VSS.n2062 0.00764286
R26683 VSS.n2204 VSS.n2109 0.00764286
R26684 VSS.n2164 VSS.n2125 0.00764286
R26685 VSS.n2165 VSS.n2164 0.00764286
R26686 VSS.n2048 VSS.n2047 0.00764286
R26687 VSS.n2048 VSS.n2037 0.00764286
R26688 VSS.n2052 VSS.n2038 0.00764286
R26689 VSS.n2243 VSS.n2034 0.00764286
R26690 VSS.n2227 VSS.n2063 0.00764286
R26691 VSS.n2226 VSS.n2225 0.00764286
R26692 VSS.n2118 VSS.n2107 0.00764286
R26693 VSS.n2198 VSS.n2197 0.00764286
R26694 VSS.n2163 VSS.n2162 0.00764286
R26695 VSS.n2163 VSS.n2161 0.00764286
R26696 VSS.n1835 VSS.n1762 0.00764286
R26697 VSS.n1843 VSS.n1842 0.00764286
R26698 VSS.n1747 VSS.n1746 0.00764286
R26699 VSS.n1866 VSS.n1737 0.00764286
R26700 VSS.n1893 VSS.n1717 0.00764286
R26701 VSS.n3542 VSS.n3536 0.00764286
R26702 VSS.n3715 VSS.n3489 0.00764286
R26703 VSS.n3753 VSS.n3461 0.00764286
R26704 VSS.n3690 VSS.n3500 0.00764286
R26705 VSS.n3718 VSS.n3717 0.00764286
R26706 VSS.n3725 VSS.n3482 0.00764286
R26707 VSS.n3721 VSS.n3720 0.00764286
R26708 VSS.n3743 VSS.n3468 0.00764286
R26709 VSS.n3757 VSS.n3462 0.00764286
R26710 VSS.n3823 VSS.n3822 0.00764286
R26711 VSS.n3821 VSS.n3426 0.00764286
R26712 VSS.n3853 VSS.n3412 0.00764286
R26713 VSS.n3905 VSS.n3393 0.00764286
R26714 VSS.n3938 VSS.n3376 0.00764286
R26715 VSS.n3934 VSS.n3376 0.00764286
R26716 VSS.n3818 VSS.n3817 0.00764286
R26717 VSS.n3818 VSS.n3431 0.00764286
R26718 VSS.n3824 VSS.n3432 0.00764286
R26719 VSS.n3820 VSS.n3428 0.00764286
R26720 VSS.n3839 VSS.n3838 0.00764286
R26721 VSS.n3854 VSS.n3411 0.00764286
R26722 VSS.n3876 VSS.n3875 0.00764286
R26723 VSS.n3912 VSS.n3389 0.00764286
R26724 VSS.n3937 VSS.n3936 0.00764286
R26725 VSS.n3936 VSS.n3935 0.00764286
R26726 VSS.n3629 VSS.n3556 0.00764286
R26727 VSS.n3637 VSS.n3636 0.00764286
R26728 VSS.n3541 VSS.n3540 0.00764286
R26729 VSS.n3660 VSS.n3531 0.00764286
R26730 VSS.n3687 VSS.n3511 0.00764286
R26731 VSS.n4134 VSS.n4128 0.00764286
R26732 VSS.n4307 VSS.n4081 0.00764286
R26733 VSS.n4345 VSS.n4053 0.00764286
R26734 VSS.n4282 VSS.n4092 0.00764286
R26735 VSS.n4310 VSS.n4309 0.00764286
R26736 VSS.n4317 VSS.n4074 0.00764286
R26737 VSS.n4313 VSS.n4312 0.00764286
R26738 VSS.n4335 VSS.n4060 0.00764286
R26739 VSS.n4349 VSS.n4054 0.00764286
R26740 VSS.n4415 VSS.n4414 0.00764286
R26741 VSS.n4413 VSS.n4018 0.00764286
R26742 VSS.n4445 VSS.n4004 0.00764286
R26743 VSS.n4497 VSS.n3985 0.00764286
R26744 VSS.n4530 VSS.n3968 0.00764286
R26745 VSS.n4526 VSS.n3968 0.00764286
R26746 VSS.n4410 VSS.n4409 0.00764286
R26747 VSS.n4410 VSS.n4023 0.00764286
R26748 VSS.n4416 VSS.n4024 0.00764286
R26749 VSS.n4412 VSS.n4020 0.00764286
R26750 VSS.n4431 VSS.n4430 0.00764286
R26751 VSS.n4446 VSS.n4003 0.00764286
R26752 VSS.n4468 VSS.n4467 0.00764286
R26753 VSS.n4504 VSS.n3981 0.00764286
R26754 VSS.n4529 VSS.n4528 0.00764286
R26755 VSS.n4528 VSS.n4527 0.00764286
R26756 VSS.n4221 VSS.n4148 0.00764286
R26757 VSS.n4229 VSS.n4228 0.00764286
R26758 VSS.n4133 VSS.n4132 0.00764286
R26759 VSS.n4252 VSS.n4123 0.00764286
R26760 VSS.n4279 VSS.n4103 0.00764286
R26761 VSS.n4726 VSS.n4720 0.00764286
R26762 VSS.n4899 VSS.n4673 0.00764286
R26763 VSS.n4937 VSS.n4645 0.00764286
R26764 VSS.n4874 VSS.n4684 0.00764286
R26765 VSS.n4902 VSS.n4901 0.00764286
R26766 VSS.n4909 VSS.n4666 0.00764286
R26767 VSS.n4905 VSS.n4904 0.00764286
R26768 VSS.n4927 VSS.n4652 0.00764286
R26769 VSS.n4941 VSS.n4646 0.00764286
R26770 VSS.n5007 VSS.n5006 0.00764286
R26771 VSS.n5005 VSS.n4610 0.00764286
R26772 VSS.n5037 VSS.n4596 0.00764286
R26773 VSS.n5089 VSS.n4577 0.00764286
R26774 VSS.n5122 VSS.n4560 0.00764286
R26775 VSS.n5118 VSS.n4560 0.00764286
R26776 VSS.n5002 VSS.n5001 0.00764286
R26777 VSS.n5002 VSS.n4615 0.00764286
R26778 VSS.n5008 VSS.n4616 0.00764286
R26779 VSS.n5004 VSS.n4612 0.00764286
R26780 VSS.n5023 VSS.n5022 0.00764286
R26781 VSS.n5038 VSS.n4595 0.00764286
R26782 VSS.n5060 VSS.n5059 0.00764286
R26783 VSS.n5096 VSS.n4573 0.00764286
R26784 VSS.n5121 VSS.n5120 0.00764286
R26785 VSS.n5120 VSS.n5119 0.00764286
R26786 VSS.n4813 VSS.n4740 0.00764286
R26787 VSS.n4821 VSS.n4820 0.00764286
R26788 VSS.n4725 VSS.n4724 0.00764286
R26789 VSS.n4844 VSS.n4715 0.00764286
R26790 VSS.n4871 VSS.n4695 0.00764286
R26791 VSS.n5318 VSS.n5312 0.00764286
R26792 VSS.n5491 VSS.n5265 0.00764286
R26793 VSS.n5529 VSS.n5237 0.00764286
R26794 VSS.n5466 VSS.n5276 0.00764286
R26795 VSS.n5494 VSS.n5493 0.00764286
R26796 VSS.n5501 VSS.n5258 0.00764286
R26797 VSS.n5497 VSS.n5496 0.00764286
R26798 VSS.n5519 VSS.n5244 0.00764286
R26799 VSS.n5533 VSS.n5238 0.00764286
R26800 VSS.n5599 VSS.n5598 0.00764286
R26801 VSS.n5597 VSS.n5202 0.00764286
R26802 VSS.n5629 VSS.n5188 0.00764286
R26803 VSS.n5681 VSS.n5169 0.00764286
R26804 VSS.n5714 VSS.n5152 0.00764286
R26805 VSS.n5710 VSS.n5152 0.00764286
R26806 VSS.n5594 VSS.n5593 0.00764286
R26807 VSS.n5594 VSS.n5207 0.00764286
R26808 VSS.n5600 VSS.n5208 0.00764286
R26809 VSS.n5596 VSS.n5204 0.00764286
R26810 VSS.n5615 VSS.n5614 0.00764286
R26811 VSS.n5630 VSS.n5187 0.00764286
R26812 VSS.n5652 VSS.n5651 0.00764286
R26813 VSS.n5688 VSS.n5165 0.00764286
R26814 VSS.n5713 VSS.n5712 0.00764286
R26815 VSS.n5712 VSS.n5711 0.00764286
R26816 VSS.n5405 VSS.n5332 0.00764286
R26817 VSS.n5413 VSS.n5412 0.00764286
R26818 VSS.n5317 VSS.n5316 0.00764286
R26819 VSS.n5436 VSS.n5307 0.00764286
R26820 VSS.n5463 VSS.n5287 0.00764286
R26821 VSS.n5910 VSS.n5904 0.00764286
R26822 VSS.n6083 VSS.n5857 0.00764286
R26823 VSS.n6121 VSS.n5829 0.00764286
R26824 VSS.n6058 VSS.n5868 0.00764286
R26825 VSS.n6086 VSS.n6085 0.00764286
R26826 VSS.n6093 VSS.n5850 0.00764286
R26827 VSS.n6089 VSS.n6088 0.00764286
R26828 VSS.n6111 VSS.n5836 0.00764286
R26829 VSS.n6125 VSS.n5830 0.00764286
R26830 VSS.n6191 VSS.n6190 0.00764286
R26831 VSS.n6189 VSS.n5794 0.00764286
R26832 VSS.n6221 VSS.n5780 0.00764286
R26833 VSS.n6273 VSS.n5761 0.00764286
R26834 VSS.n6306 VSS.n5744 0.00764286
R26835 VSS.n6302 VSS.n5744 0.00764286
R26836 VSS.n6186 VSS.n6185 0.00764286
R26837 VSS.n6186 VSS.n5799 0.00764286
R26838 VSS.n6192 VSS.n5800 0.00764286
R26839 VSS.n6188 VSS.n5796 0.00764286
R26840 VSS.n6207 VSS.n6206 0.00764286
R26841 VSS.n6222 VSS.n5779 0.00764286
R26842 VSS.n6244 VSS.n6243 0.00764286
R26843 VSS.n6280 VSS.n5757 0.00764286
R26844 VSS.n6305 VSS.n6304 0.00764286
R26845 VSS.n6304 VSS.n6303 0.00764286
R26846 VSS.n5997 VSS.n5924 0.00764286
R26847 VSS.n6005 VSS.n6004 0.00764286
R26848 VSS.n5909 VSS.n5908 0.00764286
R26849 VSS.n6028 VSS.n5899 0.00764286
R26850 VSS.n6055 VSS.n5879 0.00764286
R26851 VSS.n6502 VSS.n6496 0.00764286
R26852 VSS.n6675 VSS.n6449 0.00764286
R26853 VSS.n6713 VSS.n6421 0.00764286
R26854 VSS.n6650 VSS.n6460 0.00764286
R26855 VSS.n6678 VSS.n6677 0.00764286
R26856 VSS.n6685 VSS.n6442 0.00764286
R26857 VSS.n6681 VSS.n6680 0.00764286
R26858 VSS.n6703 VSS.n6428 0.00764286
R26859 VSS.n6717 VSS.n6422 0.00764286
R26860 VSS.n6783 VSS.n6782 0.00764286
R26861 VSS.n6781 VSS.n6386 0.00764286
R26862 VSS.n6813 VSS.n6372 0.00764286
R26863 VSS.n6865 VSS.n6353 0.00764286
R26864 VSS.n6898 VSS.n6336 0.00764286
R26865 VSS.n6894 VSS.n6336 0.00764286
R26866 VSS.n6778 VSS.n6777 0.00764286
R26867 VSS.n6778 VSS.n6391 0.00764286
R26868 VSS.n6784 VSS.n6392 0.00764286
R26869 VSS.n6780 VSS.n6388 0.00764286
R26870 VSS.n6799 VSS.n6798 0.00764286
R26871 VSS.n6814 VSS.n6371 0.00764286
R26872 VSS.n6836 VSS.n6835 0.00764286
R26873 VSS.n6872 VSS.n6349 0.00764286
R26874 VSS.n6897 VSS.n6896 0.00764286
R26875 VSS.n6896 VSS.n6895 0.00764286
R26876 VSS.n6589 VSS.n6516 0.00764286
R26877 VSS.n6597 VSS.n6596 0.00764286
R26878 VSS.n6501 VSS.n6500 0.00764286
R26879 VSS.n6620 VSS.n6491 0.00764286
R26880 VSS.n6647 VSS.n6471 0.00764286
R26881 VSS.n2346 VSS.n2340 0.00764286
R26882 VSS.n2573 VSS.n2572 0.00764286
R26883 VSS.n2596 VSS.n2595 0.00764286
R26884 VSS.n7042 VSS.n7041 0.00764286
R26885 VSS.n7033 VSS.n2500 0.00764286
R26886 VSS.n2570 VSS.n2502 0.00764286
R26887 VSS.n2507 VSS.n2506 0.00764286
R26888 VSS.n2515 VSS.n2514 0.00764286
R26889 VSS.n2598 VSS.n2516 0.00764286
R26890 VSS.n2649 VSS.n2648 0.00764286
R26891 VSS.n6988 VSS.n2630 0.00764286
R26892 VSS.n6968 VSS.n2660 0.00764286
R26893 VSS.n6948 VSS.n2707 0.00764286
R26894 VSS.n2762 VSS.n2723 0.00764286
R26895 VSS.n2763 VSS.n2762 0.00764286
R26896 VSS.n2646 VSS.n2645 0.00764286
R26897 VSS.n2646 VSS.n2635 0.00764286
R26898 VSS.n2650 VSS.n2636 0.00764286
R26899 VSS.n6987 VSS.n2632 0.00764286
R26900 VSS.n6971 VSS.n2661 0.00764286
R26901 VSS.n6970 VSS.n6969 0.00764286
R26902 VSS.n2716 VSS.n2705 0.00764286
R26903 VSS.n6942 VSS.n6941 0.00764286
R26904 VSS.n2761 VSS.n2760 0.00764286
R26905 VSS.n2761 VSS.n2759 0.00764286
R26906 VSS.n2433 VSS.n2360 0.00764286
R26907 VSS.n2441 VSS.n2440 0.00764286
R26908 VSS.n2345 VSS.n2344 0.00764286
R26909 VSS.n2464 VSS.n2335 0.00764286
R26910 VSS.n2491 VSS.n2315 0.00764286
R26911 VSS.n3061 VSS.n2943 0.00764286
R26912 VSS.n3123 VSS.n2896 0.00764286
R26913 VSS.n3161 VSS.n2868 0.00764286
R26914 VSS.n3098 VSS.n2907 0.00764286
R26915 VSS.n3126 VSS.n3125 0.00764286
R26916 VSS.n3133 VSS.n2889 0.00764286
R26917 VSS.n3129 VSS.n3128 0.00764286
R26918 VSS.n3151 VSS.n2875 0.00764286
R26919 VSS.n3165 VSS.n2869 0.00764286
R26920 VSS.n3231 VSS.n3230 0.00764286
R26921 VSS.n3229 VSS.n2833 0.00764286
R26922 VSS.n3261 VSS.n2819 0.00764286
R26923 VSS.n3313 VSS.n2800 0.00764286
R26924 VSS.n3346 VSS.n2783 0.00764286
R26925 VSS.n3342 VSS.n2783 0.00764286
R26926 VSS.n3226 VSS.n3225 0.00764286
R26927 VSS.n3226 VSS.n2838 0.00764286
R26928 VSS.n3232 VSS.n2839 0.00764286
R26929 VSS.n3228 VSS.n2835 0.00764286
R26930 VSS.n3247 VSS.n3246 0.00764286
R26931 VSS.n3262 VSS.n2818 0.00764286
R26932 VSS.n3284 VSS.n3283 0.00764286
R26933 VSS.n3320 VSS.n2796 0.00764286
R26934 VSS.n3345 VSS.n3344 0.00764286
R26935 VSS.n3344 VSS.n3343 0.00764286
R26936 VSS.n3024 VSS.n3023 0.00764286
R26937 VSS.n3046 VSS.n2950 0.00764286
R26938 VSS.n3060 VSS.n3059 0.00764286
R26939 VSS.n3058 VSS.n3054 0.00764286
R26940 VSS.n3095 VSS.n2918 0.00764286
R26941 VSS.n375 VSS.n372 0.00764286
R26942 VSS.n9083 VSS.n163 0.00764286
R26943 VSS.n9121 VSS.n135 0.00764286
R26944 VSS.n9058 VSS.n174 0.00764286
R26945 VSS.n9086 VSS.n9085 0.00764286
R26946 VSS.n9093 VSS.n156 0.00764286
R26947 VSS.n9089 VSS.n9088 0.00764286
R26948 VSS.n9111 VSS.n142 0.00764286
R26949 VSS.n9125 VSS.n136 0.00764286
R26950 VSS.n9191 VSS.n9190 0.00764286
R26951 VSS.n9189 VSS.n100 0.00764286
R26952 VSS.n9221 VSS.n86 0.00764286
R26953 VSS.n9273 VSS.n67 0.00764286
R26954 VSS.n9306 VSS.n50 0.00764286
R26955 VSS.n9302 VSS.n50 0.00764286
R26956 VSS.n9186 VSS.n9185 0.00764286
R26957 VSS.n9186 VSS.n105 0.00764286
R26958 VSS.n9192 VSS.n106 0.00764286
R26959 VSS.n9188 VSS.n102 0.00764286
R26960 VSS.n9207 VSS.n9206 0.00764286
R26961 VSS.n9222 VSS.n85 0.00764286
R26962 VSS.n9244 VSS.n9243 0.00764286
R26963 VSS.n9280 VSS.n63 0.00764286
R26964 VSS.n9305 VSS.n9304 0.00764286
R26965 VSS.n9304 VSS.n9303 0.00764286
R26966 VSS.n290 VSS.n289 0.00764286
R26967 VSS.n299 VSS.n298 0.00764286
R26968 VSS.n374 VSS.n373 0.00764286
R26969 VSS.n405 VSS.n303 0.00764286
R26970 VSS.n9055 VSS.n178 0.00764286
R26971 VSS.n565 VSS.n564 0.00764286
R26972 VSS.n588 VSS.n587 0.00764286
R26973 VSS.n862 VSS.n480 0.00764286
R26974 VSS.n852 VSS.n489 0.00764286
R26975 VSS.n562 VSS.n491 0.00764286
R26976 VSS.n496 VSS.n495 0.00764286
R26977 VSS.n504 VSS.n503 0.00764286
R26978 VSS.n590 VSS.n505 0.00764286
R26979 VSS.n641 VSS.n640 0.00764286
R26980 VSS.n807 VSS.n622 0.00764286
R26981 VSS.n787 VSS.n652 0.00764286
R26982 VSS.n767 VSS.n699 0.00764286
R26983 VSS.n726 VSS.n715 0.00764286
R26984 VSS.n722 VSS.n715 0.00764286
R26985 VSS.n638 VSS.n637 0.00764286
R26986 VSS.n638 VSS.n627 0.00764286
R26987 VSS.n642 VSS.n628 0.00764286
R26988 VSS.n806 VSS.n624 0.00764286
R26989 VSS.n790 VSS.n653 0.00764286
R26990 VSS.n789 VSS.n788 0.00764286
R26991 VSS.n708 VSS.n697 0.00764286
R26992 VSS.n761 VSS.n760 0.00764286
R26993 VSS.n725 VSS.n724 0.00764286
R26994 VSS.n724 VSS.n723 0.00764286
R26995 VSS.n456 VSS.n455 0.00764286
R26996 VSS.n465 VSS.n464 0.00764286
R26997 VSS.n933 VSS.n932 0.00764286
R26998 VSS.n970 VSS.n469 0.00764286
R26999 VSS.n865 VSS.n476 0.00764286
R27000 VSS.n7217 VSS.n7216 0.00764286
R27001 VSS.n8416 VSS.n7198 0.00764286
R27002 VSS.n8396 VSS.n7228 0.00764286
R27003 VSS.n8376 VSS.n7275 0.00764286
R27004 VSS.n7330 VSS.n7291 0.00764286
R27005 VSS.n7331 VSS.n7330 0.00764286
R27006 VSS.n7214 VSS.n7213 0.00764286
R27007 VSS.n7214 VSS.n7203 0.00764286
R27008 VSS.n7218 VSS.n7204 0.00764286
R27009 VSS.n8415 VSS.n7200 0.00764286
R27010 VSS.n8399 VSS.n7229 0.00764286
R27011 VSS.n8398 VSS.n8397 0.00764286
R27012 VSS.n7284 VSS.n7273 0.00764286
R27013 VSS.n8370 VSS.n8369 0.00764286
R27014 VSS.n7329 VSS.n7328 0.00764286
R27015 VSS.n7329 VSS.n7327 0.00764286
R27016 VSS.n7140 VSS.n7137 0.00675
R27017 VSS.n8457 VSS.n8456 0.00675
R27018 VSS.n7167 VSS.n7164 0.00675
R27019 VSS.n7139 VSS.n7138 0.00675
R27020 VSS.n8458 VSS.n7071 0.00675
R27021 VSS.n8446 VSS.n7083 0.00675
R27022 VSS.n7166 VSS.n7165 0.00675
R27023 VSS.n8442 VSS.n7087 0.00675
R27024 VSS.n898 VSS.n893 0.00675
R27025 VSS.n885 VSS.n453 0.00675
R27026 VSS.n975 VSS.n463 0.00675
R27027 VSS.n931 VSS.n930 0.00675
R27028 VSS.n7465 VSS.n7456 0.00675
R27029 VSS.n7459 VSS.n7457 0.00675
R27030 VSS.n7556 VSS.n7437 0.00675
R27031 VSS.n1079 VSS.n1074 0.00675
R27032 VSS.n1066 VSS.n1020 0.00675
R27033 VSS.n8496 VSS.n1030 0.00675
R27034 VSS.n1112 VSS.n1111 0.00675
R27035 VSS.n1022 VSS.n1019 0.00675
R27036 VSS.n8495 VSS.n8494 0.00675
R27037 VSS.n1114 VSS.n1033 0.00675
R27038 VSS.n7620 VSS.n7619 0.00675
R27039 VSS.n7638 VSS.n7388 0.00675
R27040 VSS.n7659 VSS.n7384 0.00675
R27041 VSS.n7661 VSS.n7660 0.00675
R27042 VSS.n7684 VSS.n7682 0.00675
R27043 VSS.n7730 VSS.n7352 0.00675
R27044 VSS.n7618 VSS.n7408 0.00675
R27045 VSS.n7637 VSS.n7387 0.00675
R27046 VSS.n7658 VSS.n7657 0.00675
R27047 VSS.n7685 VSS.n7672 0.00675
R27048 VSS.n7732 VSS.n7731 0.00675
R27049 VSS.n7727 VSS.n7340 0.00675
R27050 VSS.n7463 VSS.n7458 0.00675
R27051 VSS.n7522 VSS.n7460 0.00675
R27052 VSS.n7444 VSS.n7441 0.00675
R27053 VSS.n7555 VSS.n7554 0.00675
R27054 VSS.n7553 VSS.n7549 0.00675
R27055 VSS.n7879 VSS.n7870 0.00675
R27056 VSS.n7873 VSS.n7871 0.00675
R27057 VSS.n8148 VSS.n7851 0.00675
R27058 VSS.n7984 VSS.n7963 0.00675
R27059 VSS.n7955 VSS.n7954 0.00675
R27060 VSS.n8046 VSS.n7925 0.00675
R27061 VSS.n7933 VSS.n7932 0.00675
R27062 VSS.n8020 VSS.n8019 0.00675
R27063 VSS.n8047 VSS.n7923 0.00675
R27064 VSS.n7930 VSS.n7924 0.00675
R27065 VSS.n8212 VSS.n8211 0.00675
R27066 VSS.n8230 VSS.n7802 0.00675
R27067 VSS.n8251 VSS.n7798 0.00675
R27068 VSS.n8253 VSS.n8252 0.00675
R27069 VSS.n8276 VSS.n8274 0.00675
R27070 VSS.n8322 VSS.n7766 0.00675
R27071 VSS.n8210 VSS.n7822 0.00675
R27072 VSS.n8229 VSS.n7801 0.00675
R27073 VSS.n8250 VSS.n8249 0.00675
R27074 VSS.n8277 VSS.n8264 0.00675
R27075 VSS.n8324 VSS.n8323 0.00675
R27076 VSS.n8319 VSS.n7754 0.00675
R27077 VSS.n7877 VSS.n7872 0.00675
R27078 VSS.n8114 VSS.n7874 0.00675
R27079 VSS.n7858 VSS.n7855 0.00675
R27080 VSS.n8147 VSS.n8146 0.00675
R27081 VSS.n8145 VSS.n8141 0.00675
R27082 VSS.n8545 VSS.n260 0.00675
R27083 VSS.n252 VSS.n251 0.00675
R27084 VSS.n8607 VSS.n222 0.00675
R27085 VSS.n230 VSS.n229 0.00675
R27086 VSS.n8719 VSS.n8716 0.00675
R27087 VSS.n9030 VSS.n9029 0.00675
R27088 VSS.n8746 VSS.n8743 0.00675
R27089 VSS.n8718 VSS.n8717 0.00675
R27090 VSS.n9031 VSS.n8650 0.00675
R27091 VSS.n9019 VSS.n8662 0.00675
R27092 VSS.n8745 VSS.n8744 0.00675
R27093 VSS.n9015 VSS.n8666 0.00675
R27094 VSS.n8796 VSS.n8777 0.00675
R27095 VSS.n8976 VSS.n8975 0.00675
R27096 VSS.n8969 VSS.n8808 0.00675
R27097 VSS.n8841 VSS.n8840 0.00675
R27098 VSS.n8872 VSS.n8871 0.00675
R27099 VSS.n8936 VSS.n8935 0.00675
R27100 VSS.n8784 VSS.n8783 0.00675
R27101 VSS.n8977 VSS.n8804 0.00675
R27102 VSS.n8968 VSS.n8810 0.00675
R27103 VSS.n8873 VSS.n8856 0.00675
R27104 VSS.n8934 VSS.n8888 0.00675
R27105 VSS.n8930 VSS.n8894 0.00675
R27106 VSS.n8581 VSS.n8580 0.00675
R27107 VSS.n8608 VSS.n220 0.00675
R27108 VSS.n227 VSS.n221 0.00675
R27109 VSS.n1227 VSS.n1206 0.00675
R27110 VSS.n1198 VSS.n1197 0.00675
R27111 VSS.n1289 VSS.n1168 0.00675
R27112 VSS.n1176 VSS.n1175 0.00675
R27113 VSS.n1401 VSS.n1398 0.00675
R27114 VSS.n1693 VSS.n1692 0.00675
R27115 VSS.n1428 VSS.n1425 0.00675
R27116 VSS.n1400 VSS.n1399 0.00675
R27117 VSS.n1694 VSS.n1332 0.00675
R27118 VSS.n1682 VSS.n1344 0.00675
R27119 VSS.n1427 VSS.n1426 0.00675
R27120 VSS.n1678 VSS.n1348 0.00675
R27121 VSS.n1477 VSS.n1459 0.00675
R27122 VSS.n1636 VSS.n1489 0.00675
R27123 VSS.n1520 VSS.n1514 0.00675
R27124 VSS.n1522 VSS.n1521 0.00675
R27125 VSS.n1614 VSS.n1535 0.00675
R27126 VSS.n1560 VSS.n1559 0.00675
R27127 VSS.n1465 VSS.n1461 0.00675
R27128 VSS.n1635 VSS.n1634 0.00675
R27129 VSS.n1519 VSS.n1518 0.00675
R27130 VSS.n1615 VSS.n1533 0.00675
R27131 VSS.n1561 VSS.n1553 0.00675
R27132 VSS.n1556 VSS.n2 0.00675
R27133 VSS.n1263 VSS.n1262 0.00675
R27134 VSS.n1290 VSS.n1166 0.00675
R27135 VSS.n1173 VSS.n1167 0.00675
R27136 VSS.n1800 VSS.n1779 0.00675
R27137 VSS.n1771 VSS.n1770 0.00675
R27138 VSS.n1862 VSS.n1741 0.00675
R27139 VSS.n1749 VSS.n1748 0.00675
R27140 VSS.n1974 VSS.n1971 0.00675
R27141 VSS.n2285 VSS.n2284 0.00675
R27142 VSS.n2001 VSS.n1998 0.00675
R27143 VSS.n1973 VSS.n1972 0.00675
R27144 VSS.n2286 VSS.n1905 0.00675
R27145 VSS.n2274 VSS.n1917 0.00675
R27146 VSS.n2000 VSS.n1999 0.00675
R27147 VSS.n2270 VSS.n1921 0.00675
R27148 VSS.n2050 VSS.n2032 0.00675
R27149 VSS.n2228 VSS.n2062 0.00675
R27150 VSS.n2093 VSS.n2087 0.00675
R27151 VSS.n2095 VSS.n2094 0.00675
R27152 VSS.n2206 VSS.n2108 0.00675
R27153 VSS.n2167 VSS.n2165 0.00675
R27154 VSS.n2038 VSS.n2034 0.00675
R27155 VSS.n2227 VSS.n2226 0.00675
R27156 VSS.n2092 VSS.n2091 0.00675
R27157 VSS.n2207 VSS.n2106 0.00675
R27158 VSS.n2168 VSS.n2161 0.00675
R27159 VSS.n2169 VSS.n2155 0.00675
R27160 VSS.n1836 VSS.n1835 0.00675
R27161 VSS.n1863 VSS.n1739 0.00675
R27162 VSS.n1746 VSS.n1740 0.00675
R27163 VSS.n3594 VSS.n3573 0.00675
R27164 VSS.n3565 VSS.n3564 0.00675
R27165 VSS.n3656 VSS.n3535 0.00675
R27166 VSS.n3543 VSS.n3542 0.00675
R27167 VSS.n3489 VSS.n3480 0.00675
R27168 VSS.n3483 VSS.n3481 0.00675
R27169 VSS.n3758 VSS.n3461 0.00675
R27170 VSS.n3487 VSS.n3482 0.00675
R27171 VSS.n3724 VSS.n3484 0.00675
R27172 VSS.n3468 VSS.n3465 0.00675
R27173 VSS.n3757 VSS.n3756 0.00675
R27174 VSS.n3755 VSS.n3751 0.00675
R27175 VSS.n3822 VSS.n3821 0.00675
R27176 VSS.n3840 VSS.n3412 0.00675
R27177 VSS.n3861 VSS.n3408 0.00675
R27178 VSS.n3863 VSS.n3862 0.00675
R27179 VSS.n3886 VSS.n3884 0.00675
R27180 VSS.n3934 VSS.n3933 0.00675
R27181 VSS.n3820 VSS.n3432 0.00675
R27182 VSS.n3839 VSS.n3411 0.00675
R27183 VSS.n3860 VSS.n3859 0.00675
R27184 VSS.n3887 VSS.n3874 0.00675
R27185 VSS.n3935 VSS.n3378 0.00675
R27186 VSS.n3930 VSS.n3365 0.00675
R27187 VSS.n3630 VSS.n3629 0.00675
R27188 VSS.n3657 VSS.n3533 0.00675
R27189 VSS.n3540 VSS.n3534 0.00675
R27190 VSS.n4186 VSS.n4165 0.00675
R27191 VSS.n4157 VSS.n4156 0.00675
R27192 VSS.n4248 VSS.n4127 0.00675
R27193 VSS.n4135 VSS.n4134 0.00675
R27194 VSS.n4081 VSS.n4072 0.00675
R27195 VSS.n4075 VSS.n4073 0.00675
R27196 VSS.n4350 VSS.n4053 0.00675
R27197 VSS.n4079 VSS.n4074 0.00675
R27198 VSS.n4316 VSS.n4076 0.00675
R27199 VSS.n4060 VSS.n4057 0.00675
R27200 VSS.n4349 VSS.n4348 0.00675
R27201 VSS.n4347 VSS.n4343 0.00675
R27202 VSS.n4414 VSS.n4413 0.00675
R27203 VSS.n4432 VSS.n4004 0.00675
R27204 VSS.n4453 VSS.n4000 0.00675
R27205 VSS.n4455 VSS.n4454 0.00675
R27206 VSS.n4478 VSS.n4476 0.00675
R27207 VSS.n4526 VSS.n4525 0.00675
R27208 VSS.n4412 VSS.n4024 0.00675
R27209 VSS.n4431 VSS.n4003 0.00675
R27210 VSS.n4452 VSS.n4451 0.00675
R27211 VSS.n4479 VSS.n4466 0.00675
R27212 VSS.n4527 VSS.n3970 0.00675
R27213 VSS.n4522 VSS.n3957 0.00675
R27214 VSS.n4222 VSS.n4221 0.00675
R27215 VSS.n4249 VSS.n4125 0.00675
R27216 VSS.n4132 VSS.n4126 0.00675
R27217 VSS.n4778 VSS.n4757 0.00675
R27218 VSS.n4749 VSS.n4748 0.00675
R27219 VSS.n4840 VSS.n4719 0.00675
R27220 VSS.n4727 VSS.n4726 0.00675
R27221 VSS.n4673 VSS.n4664 0.00675
R27222 VSS.n4667 VSS.n4665 0.00675
R27223 VSS.n4942 VSS.n4645 0.00675
R27224 VSS.n4671 VSS.n4666 0.00675
R27225 VSS.n4908 VSS.n4668 0.00675
R27226 VSS.n4652 VSS.n4649 0.00675
R27227 VSS.n4941 VSS.n4940 0.00675
R27228 VSS.n4939 VSS.n4935 0.00675
R27229 VSS.n5006 VSS.n5005 0.00675
R27230 VSS.n5024 VSS.n4596 0.00675
R27231 VSS.n5045 VSS.n4592 0.00675
R27232 VSS.n5047 VSS.n5046 0.00675
R27233 VSS.n5070 VSS.n5068 0.00675
R27234 VSS.n5118 VSS.n5117 0.00675
R27235 VSS.n5004 VSS.n4616 0.00675
R27236 VSS.n5023 VSS.n4595 0.00675
R27237 VSS.n5044 VSS.n5043 0.00675
R27238 VSS.n5071 VSS.n5058 0.00675
R27239 VSS.n5119 VSS.n4562 0.00675
R27240 VSS.n5114 VSS.n4549 0.00675
R27241 VSS.n4814 VSS.n4813 0.00675
R27242 VSS.n4841 VSS.n4717 0.00675
R27243 VSS.n4724 VSS.n4718 0.00675
R27244 VSS.n5370 VSS.n5349 0.00675
R27245 VSS.n5341 VSS.n5340 0.00675
R27246 VSS.n5432 VSS.n5311 0.00675
R27247 VSS.n5319 VSS.n5318 0.00675
R27248 VSS.n5265 VSS.n5256 0.00675
R27249 VSS.n5259 VSS.n5257 0.00675
R27250 VSS.n5534 VSS.n5237 0.00675
R27251 VSS.n5263 VSS.n5258 0.00675
R27252 VSS.n5500 VSS.n5260 0.00675
R27253 VSS.n5244 VSS.n5241 0.00675
R27254 VSS.n5533 VSS.n5532 0.00675
R27255 VSS.n5531 VSS.n5527 0.00675
R27256 VSS.n5598 VSS.n5597 0.00675
R27257 VSS.n5616 VSS.n5188 0.00675
R27258 VSS.n5637 VSS.n5184 0.00675
R27259 VSS.n5639 VSS.n5638 0.00675
R27260 VSS.n5662 VSS.n5660 0.00675
R27261 VSS.n5710 VSS.n5709 0.00675
R27262 VSS.n5596 VSS.n5208 0.00675
R27263 VSS.n5615 VSS.n5187 0.00675
R27264 VSS.n5636 VSS.n5635 0.00675
R27265 VSS.n5663 VSS.n5650 0.00675
R27266 VSS.n5711 VSS.n5154 0.00675
R27267 VSS.n5706 VSS.n5141 0.00675
R27268 VSS.n5406 VSS.n5405 0.00675
R27269 VSS.n5433 VSS.n5309 0.00675
R27270 VSS.n5316 VSS.n5310 0.00675
R27271 VSS.n5962 VSS.n5941 0.00675
R27272 VSS.n5933 VSS.n5932 0.00675
R27273 VSS.n6024 VSS.n5903 0.00675
R27274 VSS.n5911 VSS.n5910 0.00675
R27275 VSS.n5857 VSS.n5848 0.00675
R27276 VSS.n5851 VSS.n5849 0.00675
R27277 VSS.n6126 VSS.n5829 0.00675
R27278 VSS.n5855 VSS.n5850 0.00675
R27279 VSS.n6092 VSS.n5852 0.00675
R27280 VSS.n5836 VSS.n5833 0.00675
R27281 VSS.n6125 VSS.n6124 0.00675
R27282 VSS.n6123 VSS.n6119 0.00675
R27283 VSS.n6190 VSS.n6189 0.00675
R27284 VSS.n6208 VSS.n5780 0.00675
R27285 VSS.n6229 VSS.n5776 0.00675
R27286 VSS.n6231 VSS.n6230 0.00675
R27287 VSS.n6254 VSS.n6252 0.00675
R27288 VSS.n6302 VSS.n6301 0.00675
R27289 VSS.n6188 VSS.n5800 0.00675
R27290 VSS.n6207 VSS.n5779 0.00675
R27291 VSS.n6228 VSS.n6227 0.00675
R27292 VSS.n6255 VSS.n6242 0.00675
R27293 VSS.n6303 VSS.n5746 0.00675
R27294 VSS.n6298 VSS.n5733 0.00675
R27295 VSS.n5998 VSS.n5997 0.00675
R27296 VSS.n6025 VSS.n5901 0.00675
R27297 VSS.n5908 VSS.n5902 0.00675
R27298 VSS.n6554 VSS.n6533 0.00675
R27299 VSS.n6525 VSS.n6524 0.00675
R27300 VSS.n6616 VSS.n6495 0.00675
R27301 VSS.n6503 VSS.n6502 0.00675
R27302 VSS.n6449 VSS.n6440 0.00675
R27303 VSS.n6443 VSS.n6441 0.00675
R27304 VSS.n6718 VSS.n6421 0.00675
R27305 VSS.n6447 VSS.n6442 0.00675
R27306 VSS.n6684 VSS.n6444 0.00675
R27307 VSS.n6428 VSS.n6425 0.00675
R27308 VSS.n6717 VSS.n6716 0.00675
R27309 VSS.n6715 VSS.n6711 0.00675
R27310 VSS.n6782 VSS.n6781 0.00675
R27311 VSS.n6800 VSS.n6372 0.00675
R27312 VSS.n6821 VSS.n6368 0.00675
R27313 VSS.n6823 VSS.n6822 0.00675
R27314 VSS.n6846 VSS.n6844 0.00675
R27315 VSS.n6894 VSS.n6893 0.00675
R27316 VSS.n6780 VSS.n6392 0.00675
R27317 VSS.n6799 VSS.n6371 0.00675
R27318 VSS.n6820 VSS.n6819 0.00675
R27319 VSS.n6847 VSS.n6834 0.00675
R27320 VSS.n6895 VSS.n6338 0.00675
R27321 VSS.n6890 VSS.n6325 0.00675
R27322 VSS.n6590 VSS.n6589 0.00675
R27323 VSS.n6617 VSS.n6493 0.00675
R27324 VSS.n6500 VSS.n6494 0.00675
R27325 VSS.n2398 VSS.n2377 0.00675
R27326 VSS.n2369 VSS.n2368 0.00675
R27327 VSS.n2460 VSS.n2339 0.00675
R27328 VSS.n2347 VSS.n2346 0.00675
R27329 VSS.n2572 VSS.n2569 0.00675
R27330 VSS.n7029 VSS.n7028 0.00675
R27331 VSS.n2599 VSS.n2596 0.00675
R27332 VSS.n2571 VSS.n2570 0.00675
R27333 VSS.n7030 VSS.n2503 0.00675
R27334 VSS.n7018 VSS.n2515 0.00675
R27335 VSS.n2598 VSS.n2597 0.00675
R27336 VSS.n7014 VSS.n2519 0.00675
R27337 VSS.n2648 VSS.n2630 0.00675
R27338 VSS.n6972 VSS.n2660 0.00675
R27339 VSS.n2691 VSS.n2685 0.00675
R27340 VSS.n2693 VSS.n2692 0.00675
R27341 VSS.n6950 VSS.n2706 0.00675
R27342 VSS.n2765 VSS.n2763 0.00675
R27343 VSS.n2636 VSS.n2632 0.00675
R27344 VSS.n6971 VSS.n6970 0.00675
R27345 VSS.n2690 VSS.n2689 0.00675
R27346 VSS.n6951 VSS.n2704 0.00675
R27347 VSS.n2766 VSS.n2759 0.00675
R27348 VSS.n2767 VSS.n2753 0.00675
R27349 VSS.n2434 VSS.n2433 0.00675
R27350 VSS.n2461 VSS.n2337 0.00675
R27351 VSS.n2344 VSS.n2338 0.00675
R27352 VSS.n2995 VSS.n2976 0.00675
R27353 VSS.n3030 VSS.n3029 0.00675
R27354 VSS.n3050 VSS.n3049 0.00675
R27355 VSS.n3056 VSS.n2943 0.00675
R27356 VSS.n2896 VSS.n2887 0.00675
R27357 VSS.n2890 VSS.n2888 0.00675
R27358 VSS.n3166 VSS.n2868 0.00675
R27359 VSS.n2894 VSS.n2889 0.00675
R27360 VSS.n3132 VSS.n2891 0.00675
R27361 VSS.n2875 VSS.n2872 0.00675
R27362 VSS.n3165 VSS.n3164 0.00675
R27363 VSS.n3163 VSS.n3159 0.00675
R27364 VSS.n3230 VSS.n3229 0.00675
R27365 VSS.n3248 VSS.n2819 0.00675
R27366 VSS.n3269 VSS.n2815 0.00675
R27367 VSS.n3271 VSS.n3270 0.00675
R27368 VSS.n3294 VSS.n3292 0.00675
R27369 VSS.n3342 VSS.n3341 0.00675
R27370 VSS.n3228 VSS.n2839 0.00675
R27371 VSS.n3247 VSS.n2818 0.00675
R27372 VSS.n3268 VSS.n3267 0.00675
R27373 VSS.n3295 VSS.n3282 0.00675
R27374 VSS.n3343 VSS.n2785 0.00675
R27375 VSS.n3338 VSS.n2772 0.00675
R27376 VSS.n3024 VSS.n2968 0.00675
R27377 VSS.n3051 VSS.n2947 0.00675
R27378 VSS.n3060 VSS.n2944 0.00675
R27379 VSS.n339 VSS.n338 0.00675
R27380 VSS.n354 VSS.n287 0.00675
R27381 VSS.n410 VSS.n297 0.00675
R27382 VSS.n376 VSS.n375 0.00675
R27383 VSS.n163 VSS.n154 0.00675
R27384 VSS.n157 VSS.n155 0.00675
R27385 VSS.n9126 VSS.n135 0.00675
R27386 VSS.n161 VSS.n156 0.00675
R27387 VSS.n9092 VSS.n158 0.00675
R27388 VSS.n142 VSS.n139 0.00675
R27389 VSS.n9125 VSS.n9124 0.00675
R27390 VSS.n9123 VSS.n9119 0.00675
R27391 VSS.n9190 VSS.n9189 0.00675
R27392 VSS.n9208 VSS.n86 0.00675
R27393 VSS.n9229 VSS.n82 0.00675
R27394 VSS.n9231 VSS.n9230 0.00675
R27395 VSS.n9254 VSS.n9252 0.00675
R27396 VSS.n9302 VSS.n9301 0.00675
R27397 VSS.n9188 VSS.n106 0.00675
R27398 VSS.n9207 VSS.n85 0.00675
R27399 VSS.n9228 VSS.n9227 0.00675
R27400 VSS.n9255 VSS.n9242 0.00675
R27401 VSS.n9303 VSS.n52 0.00675
R27402 VSS.n9298 VSS.n39 0.00675
R27403 VSS.n289 VSS.n286 0.00675
R27404 VSS.n409 VSS.n408 0.00675
R27405 VSS.n373 VSS.n300 0.00675
R27406 VSS.n564 VSS.n561 0.00675
R27407 VSS.n848 VSS.n847 0.00675
R27408 VSS.n591 VSS.n588 0.00675
R27409 VSS.n563 VSS.n562 0.00675
R27410 VSS.n849 VSS.n492 0.00675
R27411 VSS.n837 VSS.n504 0.00675
R27412 VSS.n590 VSS.n589 0.00675
R27413 VSS.n833 VSS.n508 0.00675
R27414 VSS.n640 VSS.n622 0.00675
R27415 VSS.n791 VSS.n652 0.00675
R27416 VSS.n683 VSS.n677 0.00675
R27417 VSS.n685 VSS.n684 0.00675
R27418 VSS.n769 VSS.n698 0.00675
R27419 VSS.n722 VSS.n721 0.00675
R27420 VSS.n628 VSS.n624 0.00675
R27421 VSS.n790 VSS.n789 0.00675
R27422 VSS.n682 VSS.n681 0.00675
R27423 VSS.n770 VSS.n696 0.00675
R27424 VSS.n723 VSS.n719 0.00675
R27425 VSS.n716 VSS.n35 0.00675
R27426 VSS.n455 VSS.n452 0.00675
R27427 VSS.n974 VSS.n973 0.00675
R27428 VSS.n933 VSS.n466 0.00675
R27429 VSS.n7216 VSS.n7198 0.00675
R27430 VSS.n8400 VSS.n7228 0.00675
R27431 VSS.n7259 VSS.n7253 0.00675
R27432 VSS.n7261 VSS.n7260 0.00675
R27433 VSS.n8378 VSS.n7274 0.00675
R27434 VSS.n7333 VSS.n7331 0.00675
R27435 VSS.n7204 VSS.n7200 0.00675
R27436 VSS.n8399 VSS.n8398 0.00675
R27437 VSS.n7258 VSS.n7257 0.00675
R27438 VSS.n8379 VSS.n7272 0.00675
R27439 VSS.n7334 VSS.n7327 0.00675
R27440 VSS.n7335 VSS.n7321 0.00675
R27441 VSS.n7589 VSS.n7588 0.00636816
R27442 VSS.n8181 VSS.n8180 0.00636816
R27443 VSS.n8787 VSS.n8771 0.00636816
R27444 VSS.n1468 VSS.n1453 0.00636816
R27445 VSS.n2041 VSS.n2026 0.00636816
R27446 VSS.n3791 VSS.n3790 0.00636816
R27447 VSS.n4383 VSS.n4382 0.00636816
R27448 VSS.n4975 VSS.n4974 0.00636816
R27449 VSS.n5567 VSS.n5566 0.00636816
R27450 VSS.n6159 VSS.n6158 0.00636816
R27451 VSS.n6751 VSS.n6750 0.00636816
R27452 VSS.n2639 VSS.n2624 0.00636816
R27453 VSS.n3199 VSS.n3198 0.00636816
R27454 VSS.n9159 VSS.n9158 0.00636816
R27455 VSS.n631 VSS.n616 0.00636816
R27456 VSS.n7207 VSS.n7192 0.00636816
R27457 VSS.n7747 VSS.n7341 0.00636785
R27458 VSS.n8339 VSS.n7755 0.00636785
R27459 VSS.n8927 VSS.n8895 0.00636785
R27460 VSS.n9347 VSS.n3 0.00636785
R27461 VSS.n2160 VSS.n2154 0.00636785
R27462 VSS.n3950 VSS.n3366 0.00636785
R27463 VSS.n4542 VSS.n3958 0.00636785
R27464 VSS.n5134 VSS.n4550 0.00636785
R27465 VSS.n5726 VSS.n5142 0.00636785
R27466 VSS.n6318 VSS.n5734 0.00636785
R27467 VSS.n6910 VSS.n6326 0.00636785
R27468 VSS.n2758 VSS.n2752 0.00636785
R27469 VSS.n3358 VSS.n2773 0.00636785
R27470 VSS.n9318 VSS.n40 0.00636785
R27471 VSS.n34 VSS.n28 0.00636785
R27472 VSS.n7326 VSS.n7320 0.00636785
R27473 VSS.n7625 VSS.n7624 0.00620714
R27474 VSS.n7624 VSS.n7386 0.00620714
R27475 VSS.n7706 VSS.n7354 0.00620714
R27476 VSS.n7724 VSS.n7354 0.00620714
R27477 VSS.n8217 VSS.n8216 0.00620714
R27478 VSS.n8216 VSS.n7800 0.00620714
R27479 VSS.n8298 VSS.n7768 0.00620714
R27480 VSS.n8316 VSS.n7768 0.00620714
R27481 VSS.n8985 VSS.n8984 0.00620714
R27482 VSS.n8984 VSS.n8983 0.00620714
R27483 VSS.n8948 VSS.n8878 0.00620714
R27484 VSS.n8891 VSS.n8878 0.00620714
R27485 VSS.n1492 VSS.n1481 0.00620714
R27486 VSS.n1497 VSS.n1492 0.00620714
R27487 VSS.n1600 VSS.n1599 0.00620714
R27488 VSS.n1599 VSS.n1598 0.00620714
R27489 VSS.n2065 VSS.n2054 0.00620714
R27490 VSS.n2070 VSS.n2065 0.00620714
R27491 VSS.n2192 VSS.n2191 0.00620714
R27492 VSS.n2191 VSS.n2190 0.00620714
R27493 VSS.n3827 VSS.n3826 0.00620714
R27494 VSS.n3826 VSS.n3410 0.00620714
R27495 VSS.n3908 VSS.n3379 0.00620714
R27496 VSS.n3926 VSS.n3379 0.00620714
R27497 VSS.n4419 VSS.n4418 0.00620714
R27498 VSS.n4418 VSS.n4002 0.00620714
R27499 VSS.n4500 VSS.n3971 0.00620714
R27500 VSS.n4518 VSS.n3971 0.00620714
R27501 VSS.n5011 VSS.n5010 0.00620714
R27502 VSS.n5010 VSS.n4594 0.00620714
R27503 VSS.n5092 VSS.n4563 0.00620714
R27504 VSS.n5110 VSS.n4563 0.00620714
R27505 VSS.n5603 VSS.n5602 0.00620714
R27506 VSS.n5602 VSS.n5186 0.00620714
R27507 VSS.n5684 VSS.n5155 0.00620714
R27508 VSS.n5702 VSS.n5155 0.00620714
R27509 VSS.n6195 VSS.n6194 0.00620714
R27510 VSS.n6194 VSS.n5778 0.00620714
R27511 VSS.n6276 VSS.n5747 0.00620714
R27512 VSS.n6294 VSS.n5747 0.00620714
R27513 VSS.n6787 VSS.n6786 0.00620714
R27514 VSS.n6786 VSS.n6370 0.00620714
R27515 VSS.n6868 VSS.n6339 0.00620714
R27516 VSS.n6886 VSS.n6339 0.00620714
R27517 VSS.n2663 VSS.n2652 0.00620714
R27518 VSS.n2668 VSS.n2663 0.00620714
R27519 VSS.n6936 VSS.n6935 0.00620714
R27520 VSS.n6935 VSS.n6934 0.00620714
R27521 VSS.n3235 VSS.n3234 0.00620714
R27522 VSS.n3234 VSS.n2817 0.00620714
R27523 VSS.n3316 VSS.n2786 0.00620714
R27524 VSS.n3334 VSS.n2786 0.00620714
R27525 VSS.n9195 VSS.n9194 0.00620714
R27526 VSS.n9194 VSS.n84 0.00620714
R27527 VSS.n9276 VSS.n53 0.00620714
R27528 VSS.n9294 VSS.n53 0.00620714
R27529 VSS.n655 VSS.n644 0.00620714
R27530 VSS.n660 VSS.n655 0.00620714
R27531 VSS.n755 VSS.n754 0.00620714
R27532 VSS.n754 VSS.n753 0.00620714
R27533 VSS.n7231 VSS.n7220 0.00620714
R27534 VSS.n7236 VSS.n7231 0.00620714
R27535 VSS.n8364 VSS.n8363 0.00620714
R27536 VSS.n8363 VSS.n8362 0.00620714
R27537 VSS.n7614 VSS.n7406 0.00587143
R27538 VSS.n7655 VSS.n7654 0.00587143
R27539 VSS.n7671 VSS.n7366 0.00587143
R27540 VSS.n7725 VSS.n7339 0.00587143
R27541 VSS.n8206 VSS.n7820 0.00587143
R27542 VSS.n8247 VSS.n8246 0.00587143
R27543 VSS.n8263 VSS.n7780 0.00587143
R27544 VSS.n8317 VSS.n7753 0.00587143
R27545 VSS.n8792 VSS.n8781 0.00587143
R27546 VSS.n8814 VSS.n8813 0.00587143
R27547 VSS.n8877 VSS.n8876 0.00587143
R27548 VSS.n8932 VSS.n8931 0.00587143
R27549 VSS.n1473 VSS.n1463 0.00587143
R27550 VSS.n1516 VSS.n1515 0.00587143
R27551 VSS.n1547 VSS.n1532 0.00587143
R27552 VSS.n1554 VSS.n1 0.00587143
R27553 VSS.n2046 VSS.n2036 0.00587143
R27554 VSS.n2089 VSS.n2088 0.00587143
R27555 VSS.n2120 VSS.n2105 0.00587143
R27556 VSS.n2172 VSS.n2171 0.00587143
R27557 VSS.n3816 VSS.n3430 0.00587143
R27558 VSS.n3857 VSS.n3856 0.00587143
R27559 VSS.n3873 VSS.n3390 0.00587143
R27560 VSS.n3928 VSS.n3364 0.00587143
R27561 VSS.n4408 VSS.n4022 0.00587143
R27562 VSS.n4449 VSS.n4448 0.00587143
R27563 VSS.n4465 VSS.n3982 0.00587143
R27564 VSS.n4520 VSS.n3956 0.00587143
R27565 VSS.n5000 VSS.n4614 0.00587143
R27566 VSS.n5041 VSS.n5040 0.00587143
R27567 VSS.n5057 VSS.n4574 0.00587143
R27568 VSS.n5112 VSS.n4548 0.00587143
R27569 VSS.n5592 VSS.n5206 0.00587143
R27570 VSS.n5633 VSS.n5632 0.00587143
R27571 VSS.n5649 VSS.n5166 0.00587143
R27572 VSS.n5704 VSS.n5140 0.00587143
R27573 VSS.n6184 VSS.n5798 0.00587143
R27574 VSS.n6225 VSS.n6224 0.00587143
R27575 VSS.n6241 VSS.n5758 0.00587143
R27576 VSS.n6296 VSS.n5732 0.00587143
R27577 VSS.n6776 VSS.n6390 0.00587143
R27578 VSS.n6817 VSS.n6816 0.00587143
R27579 VSS.n6833 VSS.n6350 0.00587143
R27580 VSS.n6888 VSS.n6324 0.00587143
R27581 VSS.n2644 VSS.n2634 0.00587143
R27582 VSS.n2687 VSS.n2686 0.00587143
R27583 VSS.n2718 VSS.n2703 0.00587143
R27584 VSS.n2770 VSS.n2769 0.00587143
R27585 VSS.n3224 VSS.n2837 0.00587143
R27586 VSS.n3265 VSS.n3264 0.00587143
R27587 VSS.n3281 VSS.n2797 0.00587143
R27588 VSS.n3336 VSS.n2771 0.00587143
R27589 VSS.n9184 VSS.n104 0.00587143
R27590 VSS.n9225 VSS.n9224 0.00587143
R27591 VSS.n9241 VSS.n64 0.00587143
R27592 VSS.n9296 VSS.n38 0.00587143
R27593 VSS.n636 VSS.n626 0.00587143
R27594 VSS.n679 VSS.n678 0.00587143
R27595 VSS.n710 VSS.n695 0.00587143
R27596 VSS.n717 VSS.n36 0.00587143
R27597 VSS.n7212 VSS.n7202 0.00587143
R27598 VSS.n7255 VSS.n7254 0.00587143
R27599 VSS.n7286 VSS.n7271 0.00587143
R27600 VSS.n7338 VSS.n7337 0.00587143
R27601 VSS.n7129 VSS.n7124 0.00585714
R27602 VSS.n7116 VSS.n7072 0.00585714
R27603 VSS.n8447 VSS.n7081 0.00585714
R27604 VSS.n7168 VSS.n7161 0.00585714
R27605 VSS.n7178 VSS.n7103 0.00585714
R27606 VSS.n8462 VSS.n7065 0.00585714
R27607 VSS.n7074 VSS.n7071 0.00585714
R27608 VSS.n8446 VSS.n8445 0.00585714
R27609 VSS.n907 VSS.n906 0.00585714
R27610 VSS.n985 VSS.n984 0.00585714
R27611 VSS.n7490 VSS.n7470 0.00585714
R27612 VSS.n7525 VSS.n7524 0.00585714
R27613 VSS.n7545 VSS.n7544 0.00585714
R27614 VSS.n7557 VSS.n7436 0.00585714
R27615 VSS.n7427 VSS.n7420 0.00585714
R27616 VSS.n1088 VSS.n1087 0.00585714
R27617 VSS.n8506 VSS.n8505 0.00585714
R27618 VSS.n1086 VSS.n1016 0.00585714
R27619 VSS.n8507 VSS.n1019 0.00585714
R27620 VSS.n8495 VSS.n1032 0.00585714
R27621 VSS.n8490 VSS.n1037 0.00585714
R27622 VSS.n7639 VSS.n7398 0.00585714
R27623 VSS.n7681 VSS.n7680 0.00585714
R27624 VSS.n7702 VSS.n7363 0.00585714
R27625 VSS.n7712 VSS.n7711 0.00585714
R27626 VSS.n7368 VSS.n7365 0.00585714
R27627 VSS.n7474 VSS.n7462 0.00585714
R27628 VSS.n7519 VSS.n7460 0.00585714
R27629 VSS.n7546 VSS.n7441 0.00585714
R27630 VSS.n8082 VSS.n7884 0.00585714
R27631 VSS.n8117 VSS.n8116 0.00585714
R27632 VSS.n8137 VSS.n8136 0.00585714
R27633 VSS.n8149 VSS.n7850 0.00585714
R27634 VSS.n7841 VSS.n7834 0.00585714
R27635 VSS.n8013 VSS.n8012 0.00585714
R27636 VSS.n8021 VSS.n7947 0.00585714
R27637 VSS.n8014 VSS.n7951 0.00585714
R27638 VSS.n8020 VSS.n7948 0.00585714
R27639 VSS.n8026 VSS.n7923 0.00585714
R27640 VSS.n8051 VSS.n7919 0.00585714
R27641 VSS.n8231 VSS.n7812 0.00585714
R27642 VSS.n8273 VSS.n8272 0.00585714
R27643 VSS.n8294 VSS.n7777 0.00585714
R27644 VSS.n8304 VSS.n8303 0.00585714
R27645 VSS.n7782 VSS.n7779 0.00585714
R27646 VSS.n7888 VSS.n7876 0.00585714
R27647 VSS.n8111 VSS.n7874 0.00585714
R27648 VSS.n8138 VSS.n7855 0.00585714
R27649 VSS.n8574 VSS.n8573 0.00585714
R27650 VSS.n8582 VSS.n244 0.00585714
R27651 VSS.n8708 VSS.n8703 0.00585714
R27652 VSS.n8695 VSS.n8651 0.00585714
R27653 VSS.n9020 VSS.n8660 0.00585714
R27654 VSS.n8747 VSS.n8740 0.00585714
R27655 VSS.n8757 VSS.n8682 0.00585714
R27656 VSS.n9035 VSS.n8644 0.00585714
R27657 VSS.n8653 VSS.n8650 0.00585714
R27658 VSS.n9019 VSS.n9018 0.00585714
R27659 VSS.n8979 VSS.n8803 0.00585714
R27660 VSS.n8870 VSS.n8869 0.00585714
R27661 VSS.n8906 VSS.n8852 0.00585714
R27662 VSS.n8910 VSS.n8909 0.00585714
R27663 VSS.n8907 VSS.n8854 0.00585714
R27664 VSS.n8575 VSS.n248 0.00585714
R27665 VSS.n8581 VSS.n245 0.00585714
R27666 VSS.n8587 VSS.n220 0.00585714
R27667 VSS.n8612 VSS.n216 0.00585714
R27668 VSS.n1256 VSS.n1255 0.00585714
R27669 VSS.n1264 VSS.n1190 0.00585714
R27670 VSS.n1390 VSS.n1385 0.00585714
R27671 VSS.n1377 VSS.n1333 0.00585714
R27672 VSS.n1683 VSS.n1342 0.00585714
R27673 VSS.n1429 VSS.n1422 0.00585714
R27674 VSS.n1439 VSS.n1364 0.00585714
R27675 VSS.n1698 VSS.n1326 0.00585714
R27676 VSS.n1335 VSS.n1332 0.00585714
R27677 VSS.n1682 VSS.n1681 0.00585714
R27678 VSS.n1637 VSS.n1488 0.00585714
R27679 VSS.n1577 VSS.n1576 0.00585714
R27680 VSS.n1608 VSS.n1539 0.00585714
R27681 VSS.n1604 VSS.n1542 0.00585714
R27682 VSS.n1607 VSS.n1606 0.00585714
R27683 VSS.n1257 VSS.n1194 0.00585714
R27684 VSS.n1263 VSS.n1191 0.00585714
R27685 VSS.n1269 VSS.n1166 0.00585714
R27686 VSS.n1294 VSS.n1162 0.00585714
R27687 VSS.n1829 VSS.n1828 0.00585714
R27688 VSS.n1837 VSS.n1763 0.00585714
R27689 VSS.n1963 VSS.n1958 0.00585714
R27690 VSS.n1950 VSS.n1906 0.00585714
R27691 VSS.n2275 VSS.n1915 0.00585714
R27692 VSS.n2002 VSS.n1995 0.00585714
R27693 VSS.n2012 VSS.n1937 0.00585714
R27694 VSS.n2290 VSS.n1899 0.00585714
R27695 VSS.n1908 VSS.n1905 0.00585714
R27696 VSS.n2274 VSS.n2273 0.00585714
R27697 VSS.n2229 VSS.n2061 0.00585714
R27698 VSS.n2137 VSS.n2136 0.00585714
R27699 VSS.n2200 VSS.n2112 0.00585714
R27700 VSS.n2196 VSS.n2115 0.00585714
R27701 VSS.n2199 VSS.n2198 0.00585714
R27702 VSS.n1830 VSS.n1767 0.00585714
R27703 VSS.n1836 VSS.n1764 0.00585714
R27704 VSS.n1842 VSS.n1739 0.00585714
R27705 VSS.n1867 VSS.n1735 0.00585714
R27706 VSS.n3623 VSS.n3622 0.00585714
R27707 VSS.n3631 VSS.n3557 0.00585714
R27708 VSS.n3692 VSS.n3494 0.00585714
R27709 VSS.n3727 VSS.n3726 0.00585714
R27710 VSS.n3747 VSS.n3746 0.00585714
R27711 VSS.n3759 VSS.n3460 0.00585714
R27712 VSS.n3451 VSS.n3444 0.00585714
R27713 VSS.n3498 VSS.n3486 0.00585714
R27714 VSS.n3721 VSS.n3484 0.00585714
R27715 VSS.n3748 VSS.n3465 0.00585714
R27716 VSS.n3841 VSS.n3422 0.00585714
R27717 VSS.n3883 VSS.n3882 0.00585714
R27718 VSS.n3904 VSS.n3387 0.00585714
R27719 VSS.n3914 VSS.n3913 0.00585714
R27720 VSS.n3392 VSS.n3389 0.00585714
R27721 VSS.n3624 VSS.n3561 0.00585714
R27722 VSS.n3630 VSS.n3558 0.00585714
R27723 VSS.n3636 VSS.n3533 0.00585714
R27724 VSS.n3661 VSS.n3529 0.00585714
R27725 VSS.n4215 VSS.n4214 0.00585714
R27726 VSS.n4223 VSS.n4149 0.00585714
R27727 VSS.n4284 VSS.n4086 0.00585714
R27728 VSS.n4319 VSS.n4318 0.00585714
R27729 VSS.n4339 VSS.n4338 0.00585714
R27730 VSS.n4351 VSS.n4052 0.00585714
R27731 VSS.n4043 VSS.n4036 0.00585714
R27732 VSS.n4090 VSS.n4078 0.00585714
R27733 VSS.n4313 VSS.n4076 0.00585714
R27734 VSS.n4340 VSS.n4057 0.00585714
R27735 VSS.n4433 VSS.n4014 0.00585714
R27736 VSS.n4475 VSS.n4474 0.00585714
R27737 VSS.n4496 VSS.n3979 0.00585714
R27738 VSS.n4506 VSS.n4505 0.00585714
R27739 VSS.n3984 VSS.n3981 0.00585714
R27740 VSS.n4216 VSS.n4153 0.00585714
R27741 VSS.n4222 VSS.n4150 0.00585714
R27742 VSS.n4228 VSS.n4125 0.00585714
R27743 VSS.n4253 VSS.n4121 0.00585714
R27744 VSS.n4807 VSS.n4806 0.00585714
R27745 VSS.n4815 VSS.n4741 0.00585714
R27746 VSS.n4876 VSS.n4678 0.00585714
R27747 VSS.n4911 VSS.n4910 0.00585714
R27748 VSS.n4931 VSS.n4930 0.00585714
R27749 VSS.n4943 VSS.n4644 0.00585714
R27750 VSS.n4635 VSS.n4628 0.00585714
R27751 VSS.n4682 VSS.n4670 0.00585714
R27752 VSS.n4905 VSS.n4668 0.00585714
R27753 VSS.n4932 VSS.n4649 0.00585714
R27754 VSS.n5025 VSS.n4606 0.00585714
R27755 VSS.n5067 VSS.n5066 0.00585714
R27756 VSS.n5088 VSS.n4571 0.00585714
R27757 VSS.n5098 VSS.n5097 0.00585714
R27758 VSS.n4576 VSS.n4573 0.00585714
R27759 VSS.n4808 VSS.n4745 0.00585714
R27760 VSS.n4814 VSS.n4742 0.00585714
R27761 VSS.n4820 VSS.n4717 0.00585714
R27762 VSS.n4845 VSS.n4713 0.00585714
R27763 VSS.n5399 VSS.n5398 0.00585714
R27764 VSS.n5407 VSS.n5333 0.00585714
R27765 VSS.n5468 VSS.n5270 0.00585714
R27766 VSS.n5503 VSS.n5502 0.00585714
R27767 VSS.n5523 VSS.n5522 0.00585714
R27768 VSS.n5535 VSS.n5236 0.00585714
R27769 VSS.n5227 VSS.n5220 0.00585714
R27770 VSS.n5274 VSS.n5262 0.00585714
R27771 VSS.n5497 VSS.n5260 0.00585714
R27772 VSS.n5524 VSS.n5241 0.00585714
R27773 VSS.n5617 VSS.n5198 0.00585714
R27774 VSS.n5659 VSS.n5658 0.00585714
R27775 VSS.n5680 VSS.n5163 0.00585714
R27776 VSS.n5690 VSS.n5689 0.00585714
R27777 VSS.n5168 VSS.n5165 0.00585714
R27778 VSS.n5400 VSS.n5337 0.00585714
R27779 VSS.n5406 VSS.n5334 0.00585714
R27780 VSS.n5412 VSS.n5309 0.00585714
R27781 VSS.n5437 VSS.n5305 0.00585714
R27782 VSS.n5991 VSS.n5990 0.00585714
R27783 VSS.n5999 VSS.n5925 0.00585714
R27784 VSS.n6060 VSS.n5862 0.00585714
R27785 VSS.n6095 VSS.n6094 0.00585714
R27786 VSS.n6115 VSS.n6114 0.00585714
R27787 VSS.n6127 VSS.n5828 0.00585714
R27788 VSS.n5819 VSS.n5812 0.00585714
R27789 VSS.n5866 VSS.n5854 0.00585714
R27790 VSS.n6089 VSS.n5852 0.00585714
R27791 VSS.n6116 VSS.n5833 0.00585714
R27792 VSS.n6209 VSS.n5790 0.00585714
R27793 VSS.n6251 VSS.n6250 0.00585714
R27794 VSS.n6272 VSS.n5755 0.00585714
R27795 VSS.n6282 VSS.n6281 0.00585714
R27796 VSS.n5760 VSS.n5757 0.00585714
R27797 VSS.n5992 VSS.n5929 0.00585714
R27798 VSS.n5998 VSS.n5926 0.00585714
R27799 VSS.n6004 VSS.n5901 0.00585714
R27800 VSS.n6029 VSS.n5897 0.00585714
R27801 VSS.n6583 VSS.n6582 0.00585714
R27802 VSS.n6591 VSS.n6517 0.00585714
R27803 VSS.n6652 VSS.n6454 0.00585714
R27804 VSS.n6687 VSS.n6686 0.00585714
R27805 VSS.n6707 VSS.n6706 0.00585714
R27806 VSS.n6719 VSS.n6420 0.00585714
R27807 VSS.n6411 VSS.n6404 0.00585714
R27808 VSS.n6458 VSS.n6446 0.00585714
R27809 VSS.n6681 VSS.n6444 0.00585714
R27810 VSS.n6708 VSS.n6425 0.00585714
R27811 VSS.n6801 VSS.n6382 0.00585714
R27812 VSS.n6843 VSS.n6842 0.00585714
R27813 VSS.n6864 VSS.n6347 0.00585714
R27814 VSS.n6874 VSS.n6873 0.00585714
R27815 VSS.n6352 VSS.n6349 0.00585714
R27816 VSS.n6584 VSS.n6521 0.00585714
R27817 VSS.n6590 VSS.n6518 0.00585714
R27818 VSS.n6596 VSS.n6493 0.00585714
R27819 VSS.n6621 VSS.n6489 0.00585714
R27820 VSS.n2427 VSS.n2426 0.00585714
R27821 VSS.n2435 VSS.n2361 0.00585714
R27822 VSS.n2561 VSS.n2556 0.00585714
R27823 VSS.n2548 VSS.n2504 0.00585714
R27824 VSS.n7019 VSS.n2513 0.00585714
R27825 VSS.n2600 VSS.n2593 0.00585714
R27826 VSS.n2610 VSS.n2535 0.00585714
R27827 VSS.n7034 VSS.n2497 0.00585714
R27828 VSS.n2506 VSS.n2503 0.00585714
R27829 VSS.n7018 VSS.n7017 0.00585714
R27830 VSS.n6973 VSS.n2659 0.00585714
R27831 VSS.n2735 VSS.n2734 0.00585714
R27832 VSS.n6944 VSS.n2710 0.00585714
R27833 VSS.n6940 VSS.n2713 0.00585714
R27834 VSS.n6943 VSS.n6942 0.00585714
R27835 VSS.n2428 VSS.n2365 0.00585714
R27836 VSS.n2434 VSS.n2362 0.00585714
R27837 VSS.n2440 VSS.n2337 0.00585714
R27838 VSS.n2465 VSS.n2333 0.00585714
R27839 VSS.n3019 VSS.n2964 0.00585714
R27840 VSS.n2967 VSS.n2965 0.00585714
R27841 VSS.n3100 VSS.n2901 0.00585714
R27842 VSS.n3135 VSS.n3134 0.00585714
R27843 VSS.n3155 VSS.n3154 0.00585714
R27844 VSS.n3167 VSS.n2867 0.00585714
R27845 VSS.n2858 VSS.n2851 0.00585714
R27846 VSS.n2905 VSS.n2893 0.00585714
R27847 VSS.n3129 VSS.n2891 0.00585714
R27848 VSS.n3156 VSS.n2872 0.00585714
R27849 VSS.n3249 VSS.n2829 0.00585714
R27850 VSS.n3291 VSS.n3290 0.00585714
R27851 VSS.n3312 VSS.n2794 0.00585714
R27852 VSS.n3322 VSS.n3321 0.00585714
R27853 VSS.n2799 VSS.n2796 0.00585714
R27854 VSS.n3020 VSS.n2966 0.00585714
R27855 VSS.n3027 VSS.n2968 0.00585714
R27856 VSS.n2950 VSS.n2947 0.00585714
R27857 VSS.n2945 VSS.n2930 0.00585714
R27858 VSS.n353 VSS.n351 0.00585714
R27859 VSS.n420 VSS.n419 0.00585714
R27860 VSS.n9060 VSS.n168 0.00585714
R27861 VSS.n9095 VSS.n9094 0.00585714
R27862 VSS.n9115 VSS.n9114 0.00585714
R27863 VSS.n9127 VSS.n134 0.00585714
R27864 VSS.n125 VSS.n118 0.00585714
R27865 VSS.n172 VSS.n160 0.00585714
R27866 VSS.n9089 VSS.n158 0.00585714
R27867 VSS.n9116 VSS.n139 0.00585714
R27868 VSS.n9209 VSS.n96 0.00585714
R27869 VSS.n9251 VSS.n9250 0.00585714
R27870 VSS.n9272 VSS.n61 0.00585714
R27871 VSS.n9282 VSS.n9281 0.00585714
R27872 VSS.n66 VSS.n63 0.00585714
R27873 VSS.n352 VSS.n283 0.00585714
R27874 VSS.n421 VSS.n286 0.00585714
R27875 VSS.n409 VSS.n299 0.00585714
R27876 VSS.n404 VSS.n304 0.00585714
R27877 VSS.n553 VSS.n550 0.00585714
R27878 VSS.n537 VSS.n493 0.00585714
R27879 VSS.n838 VSS.n502 0.00585714
R27880 VSS.n592 VSS.n585 0.00585714
R27881 VSS.n602 VSS.n524 0.00585714
R27882 VSS.n853 VSS.n486 0.00585714
R27883 VSS.n495 VSS.n492 0.00585714
R27884 VSS.n837 VSS.n836 0.00585714
R27885 VSS.n792 VSS.n651 0.00585714
R27886 VSS.n736 VSS.n735 0.00585714
R27887 VSS.n763 VSS.n702 0.00585714
R27888 VSS.n759 VSS.n705 0.00585714
R27889 VSS.n762 VSS.n761 0.00585714
R27890 VSS.n905 VSS.n449 0.00585714
R27891 VSS.n986 VSS.n452 0.00585714
R27892 VSS.n974 VSS.n465 0.00585714
R27893 VSS.n969 VSS.n470 0.00585714
R27894 VSS.n8401 VSS.n7227 0.00585714
R27895 VSS.n7303 VSS.n7302 0.00585714
R27896 VSS.n8372 VSS.n7278 0.00585714
R27897 VSS.n8368 VSS.n7281 0.00585714
R27898 VSS.n8371 VSS.n8370 0.00585714
R27899 VSS.n961 VSS.n478 0.00565497
R27900 VSS.n8482 VSS.n1045 0.00565497
R27901 VSS.n8076 VSS.n7903 0.00565497
R27902 VSS.n8637 VSS.n200 0.00565497
R27903 VSS.n1319 VSS.n1146 0.00565497
R27904 VSS.n1892 VSS.n1719 0.00565497
R27905 VSS.n3686 VSS.n3513 0.00565497
R27906 VSS.n4278 VSS.n4105 0.00565497
R27907 VSS.n4870 VSS.n4697 0.00565497
R27908 VSS.n5462 VSS.n5289 0.00565497
R27909 VSS.n6054 VSS.n5881 0.00565497
R27910 VSS.n6646 VSS.n6473 0.00565497
R27911 VSS.n2490 VSS.n2317 0.00565497
R27912 VSS.n3094 VSS.n2920 0.00565497
R27913 VSS.n9054 VSS.n180 0.00565497
R27914 VSS.n8433 VSS.n7096 0.00511752
R27915 VSS.n7610 VSS.n7414 0.00511752
R27916 VSS.n8202 VSS.n7828 0.00511752
R27917 VSS.n9006 VSS.n8675 0.00511752
R27918 VSS.n1669 VSS.n1357 0.00511752
R27919 VSS.n2261 VSS.n1930 0.00511752
R27920 VSS.n3812 VSS.n3438 0.00511752
R27921 VSS.n4404 VSS.n4030 0.00511752
R27922 VSS.n4996 VSS.n4622 0.00511752
R27923 VSS.n5588 VSS.n5214 0.00511752
R27924 VSS.n6180 VSS.n5806 0.00511752
R27925 VSS.n6772 VSS.n6398 0.00511752
R27926 VSS.n7005 VSS.n2528 0.00511752
R27927 VSS.n3220 VSS.n2845 0.00511752
R27928 VSS.n9180 VSS.n112 0.00511752
R27929 VSS.n824 VSS.n517 0.00511752
R27930 VSS.n8469 VSS.n7062 0.00496429
R27931 VSS.n8465 VSS.n7065 0.00496429
R27932 VSS.n8441 VSS.n7088 0.00496429
R27933 VSS.n8438 VSS.n7088 0.00496429
R27934 VSS.n8435 VSS.n7094 0.00496429
R27935 VSS.n935 VSS.n928 0.00496429
R27936 VSS.n946 VSS.n871 0.00496429
R27937 VSS.n1116 VSS.n1109 0.00496429
R27938 VSS.n1127 VSS.n1052 0.00496429
R27939 VSS.n8518 VSS.n1010 0.00496429
R27940 VSS.n8514 VSS.n1013 0.00496429
R27941 VSS.n8511 VSS.n1013 0.00496429
R27942 VSS.n8487 VSS.n1037 0.00496429
R27943 VSS.n8484 VSS.n1043 0.00496429
R27944 VSS.n7722 VSS.n7350 0.00496429
R27945 VSS.n7668 VSS.n7667 0.00496429
R27946 VSS.n7723 VSS.n7356 0.00496429
R27947 VSS.n7498 VSS.n7476 0.00496429
R27948 VSS.n7501 VSS.n7474 0.00496429
R27949 VSS.n7439 VSS.n7424 0.00496429
R27950 VSS.n7569 VSS.n7424 0.00496429
R27951 VSS.n7572 VSS.n7412 0.00496429
R27952 VSS.n8045 VSS.n8044 0.00496429
R27953 VSS.n7913 VSS.n7910 0.00496429
R27954 VSS.n7992 VSS.n7970 0.00496429
R27955 VSS.n7995 VSS.n7968 0.00496429
R27956 VSS.n7968 VSS.n7950 0.00496429
R27957 VSS.n8054 VSS.n7919 0.00496429
R27958 VSS.n8057 VSS.n7901 0.00496429
R27959 VSS.n8314 VSS.n7764 0.00496429
R27960 VSS.n8260 VSS.n8259 0.00496429
R27961 VSS.n8315 VSS.n7770 0.00496429
R27962 VSS.n8090 VSS.n7890 0.00496429
R27963 VSS.n8093 VSS.n7888 0.00496429
R27964 VSS.n7853 VSS.n7838 0.00496429
R27965 VSS.n8161 VSS.n7838 0.00496429
R27966 VSS.n8164 VSS.n7826 0.00496429
R27967 VSS.n8606 VSS.n8605 0.00496429
R27968 VSS.n210 VSS.n207 0.00496429
R27969 VSS.n9042 VSS.n8641 0.00496429
R27970 VSS.n9038 VSS.n8644 0.00496429
R27971 VSS.n9014 VSS.n8667 0.00496429
R27972 VSS.n9011 VSS.n8667 0.00496429
R27973 VSS.n9008 VSS.n8673 0.00496429
R27974 VSS.n8941 VSS.n8885 0.00496429
R27975 VSS.n8965 VSS.n8964 0.00496429
R27976 VSS.n8940 VSS.n8887 0.00496429
R27977 VSS.n8553 VSS.n267 0.00496429
R27978 VSS.n8556 VSS.n265 0.00496429
R27979 VSS.n265 VSS.n247 0.00496429
R27980 VSS.n8615 VSS.n216 0.00496429
R27981 VSS.n8618 VSS.n198 0.00496429
R27982 VSS.n1288 VSS.n1287 0.00496429
R27983 VSS.n1156 VSS.n1153 0.00496429
R27984 VSS.n1705 VSS.n1323 0.00496429
R27985 VSS.n1701 VSS.n1326 0.00496429
R27986 VSS.n1677 VSS.n1349 0.00496429
R27987 VSS.n1674 VSS.n1349 0.00496429
R27988 VSS.n1671 VSS.n1355 0.00496429
R27989 VSS.n1596 VSS.n1595 0.00496429
R27990 VSS.n1529 VSS.n1528 0.00496429
R27991 VSS.n1597 VSS.n1550 0.00496429
R27992 VSS.n1235 VSS.n1213 0.00496429
R27993 VSS.n1238 VSS.n1211 0.00496429
R27994 VSS.n1211 VSS.n1193 0.00496429
R27995 VSS.n1297 VSS.n1162 0.00496429
R27996 VSS.n1300 VSS.n1144 0.00496429
R27997 VSS.n1861 VSS.n1860 0.00496429
R27998 VSS.n1729 VSS.n1726 0.00496429
R27999 VSS.n2297 VSS.n1896 0.00496429
R28000 VSS.n2293 VSS.n1899 0.00496429
R28001 VSS.n2269 VSS.n1922 0.00496429
R28002 VSS.n2266 VSS.n1922 0.00496429
R28003 VSS.n2263 VSS.n1928 0.00496429
R28004 VSS.n2188 VSS.n2187 0.00496429
R28005 VSS.n2102 VSS.n2101 0.00496429
R28006 VSS.n2189 VSS.n2123 0.00496429
R28007 VSS.n1808 VSS.n1786 0.00496429
R28008 VSS.n1811 VSS.n1784 0.00496429
R28009 VSS.n1784 VSS.n1766 0.00496429
R28010 VSS.n1870 VSS.n1735 0.00496429
R28011 VSS.n1873 VSS.n1717 0.00496429
R28012 VSS.n3655 VSS.n3654 0.00496429
R28013 VSS.n3523 VSS.n3520 0.00496429
R28014 VSS.n3700 VSS.n3500 0.00496429
R28015 VSS.n3703 VSS.n3498 0.00496429
R28016 VSS.n3463 VSS.n3448 0.00496429
R28017 VSS.n3771 VSS.n3448 0.00496429
R28018 VSS.n3774 VSS.n3436 0.00496429
R28019 VSS.n3924 VSS.n3375 0.00496429
R28020 VSS.n3870 VSS.n3869 0.00496429
R28021 VSS.n3925 VSS.n3377 0.00496429
R28022 VSS.n3602 VSS.n3580 0.00496429
R28023 VSS.n3605 VSS.n3578 0.00496429
R28024 VSS.n3578 VSS.n3560 0.00496429
R28025 VSS.n3664 VSS.n3529 0.00496429
R28026 VSS.n3667 VSS.n3511 0.00496429
R28027 VSS.n4247 VSS.n4246 0.00496429
R28028 VSS.n4115 VSS.n4112 0.00496429
R28029 VSS.n4292 VSS.n4092 0.00496429
R28030 VSS.n4295 VSS.n4090 0.00496429
R28031 VSS.n4055 VSS.n4040 0.00496429
R28032 VSS.n4363 VSS.n4040 0.00496429
R28033 VSS.n4366 VSS.n4028 0.00496429
R28034 VSS.n4516 VSS.n3967 0.00496429
R28035 VSS.n4462 VSS.n4461 0.00496429
R28036 VSS.n4517 VSS.n3969 0.00496429
R28037 VSS.n4194 VSS.n4172 0.00496429
R28038 VSS.n4197 VSS.n4170 0.00496429
R28039 VSS.n4170 VSS.n4152 0.00496429
R28040 VSS.n4256 VSS.n4121 0.00496429
R28041 VSS.n4259 VSS.n4103 0.00496429
R28042 VSS.n4839 VSS.n4838 0.00496429
R28043 VSS.n4707 VSS.n4704 0.00496429
R28044 VSS.n4884 VSS.n4684 0.00496429
R28045 VSS.n4887 VSS.n4682 0.00496429
R28046 VSS.n4647 VSS.n4632 0.00496429
R28047 VSS.n4955 VSS.n4632 0.00496429
R28048 VSS.n4958 VSS.n4620 0.00496429
R28049 VSS.n5108 VSS.n4559 0.00496429
R28050 VSS.n5054 VSS.n5053 0.00496429
R28051 VSS.n5109 VSS.n4561 0.00496429
R28052 VSS.n4786 VSS.n4764 0.00496429
R28053 VSS.n4789 VSS.n4762 0.00496429
R28054 VSS.n4762 VSS.n4744 0.00496429
R28055 VSS.n4848 VSS.n4713 0.00496429
R28056 VSS.n4851 VSS.n4695 0.00496429
R28057 VSS.n5431 VSS.n5430 0.00496429
R28058 VSS.n5299 VSS.n5296 0.00496429
R28059 VSS.n5476 VSS.n5276 0.00496429
R28060 VSS.n5479 VSS.n5274 0.00496429
R28061 VSS.n5239 VSS.n5224 0.00496429
R28062 VSS.n5547 VSS.n5224 0.00496429
R28063 VSS.n5550 VSS.n5212 0.00496429
R28064 VSS.n5700 VSS.n5151 0.00496429
R28065 VSS.n5646 VSS.n5645 0.00496429
R28066 VSS.n5701 VSS.n5153 0.00496429
R28067 VSS.n5378 VSS.n5356 0.00496429
R28068 VSS.n5381 VSS.n5354 0.00496429
R28069 VSS.n5354 VSS.n5336 0.00496429
R28070 VSS.n5440 VSS.n5305 0.00496429
R28071 VSS.n5443 VSS.n5287 0.00496429
R28072 VSS.n6023 VSS.n6022 0.00496429
R28073 VSS.n5891 VSS.n5888 0.00496429
R28074 VSS.n6068 VSS.n5868 0.00496429
R28075 VSS.n6071 VSS.n5866 0.00496429
R28076 VSS.n5831 VSS.n5816 0.00496429
R28077 VSS.n6139 VSS.n5816 0.00496429
R28078 VSS.n6142 VSS.n5804 0.00496429
R28079 VSS.n6292 VSS.n5743 0.00496429
R28080 VSS.n6238 VSS.n6237 0.00496429
R28081 VSS.n6293 VSS.n5745 0.00496429
R28082 VSS.n5970 VSS.n5948 0.00496429
R28083 VSS.n5973 VSS.n5946 0.00496429
R28084 VSS.n5946 VSS.n5928 0.00496429
R28085 VSS.n6032 VSS.n5897 0.00496429
R28086 VSS.n6035 VSS.n5879 0.00496429
R28087 VSS.n6615 VSS.n6614 0.00496429
R28088 VSS.n6483 VSS.n6480 0.00496429
R28089 VSS.n6660 VSS.n6460 0.00496429
R28090 VSS.n6663 VSS.n6458 0.00496429
R28091 VSS.n6423 VSS.n6408 0.00496429
R28092 VSS.n6731 VSS.n6408 0.00496429
R28093 VSS.n6734 VSS.n6396 0.00496429
R28094 VSS.n6884 VSS.n6335 0.00496429
R28095 VSS.n6830 VSS.n6829 0.00496429
R28096 VSS.n6885 VSS.n6337 0.00496429
R28097 VSS.n6562 VSS.n6540 0.00496429
R28098 VSS.n6565 VSS.n6538 0.00496429
R28099 VSS.n6538 VSS.n6520 0.00496429
R28100 VSS.n6624 VSS.n6489 0.00496429
R28101 VSS.n6627 VSS.n6471 0.00496429
R28102 VSS.n2459 VSS.n2458 0.00496429
R28103 VSS.n2327 VSS.n2324 0.00496429
R28104 VSS.n7041 VSS.n2494 0.00496429
R28105 VSS.n7037 VSS.n2497 0.00496429
R28106 VSS.n7013 VSS.n2520 0.00496429
R28107 VSS.n7010 VSS.n2520 0.00496429
R28108 VSS.n7007 VSS.n2526 0.00496429
R28109 VSS.n6932 VSS.n6931 0.00496429
R28110 VSS.n2700 VSS.n2699 0.00496429
R28111 VSS.n6933 VSS.n2721 0.00496429
R28112 VSS.n2406 VSS.n2384 0.00496429
R28113 VSS.n2409 VSS.n2382 0.00496429
R28114 VSS.n2382 VSS.n2364 0.00496429
R28115 VSS.n2468 VSS.n2333 0.00496429
R28116 VSS.n2471 VSS.n2315 0.00496429
R28117 VSS.n3062 VSS.n2942 0.00496429
R28118 VSS.n2933 VSS.n2926 0.00496429
R28119 VSS.n3108 VSS.n2907 0.00496429
R28120 VSS.n3111 VSS.n2905 0.00496429
R28121 VSS.n2870 VSS.n2855 0.00496429
R28122 VSS.n3179 VSS.n2855 0.00496429
R28123 VSS.n3182 VSS.n2843 0.00496429
R28124 VSS.n3332 VSS.n2782 0.00496429
R28125 VSS.n3278 VSS.n3277 0.00496429
R28126 VSS.n3333 VSS.n2784 0.00496429
R28127 VSS.n3003 VSS.n2982 0.00496429
R28128 VSS.n3006 VSS.n2980 0.00496429
R28129 VSS.n2980 VSS.n2970 0.00496429
R28130 VSS.n3075 VSS.n2930 0.00496429
R28131 VSS.n3078 VSS.n2918 0.00496429
R28132 VSS.n371 VSS.n317 0.00496429
R28133 VSS.n391 VSS.n390 0.00496429
R28134 VSS.n9068 VSS.n174 0.00496429
R28135 VSS.n9071 VSS.n172 0.00496429
R28136 VSS.n137 VSS.n122 0.00496429
R28137 VSS.n9139 VSS.n122 0.00496429
R28138 VSS.n9142 VSS.n110 0.00496429
R28139 VSS.n9292 VSS.n49 0.00496429
R28140 VSS.n9238 VSS.n9237 0.00496429
R28141 VSS.n9293 VSS.n51 0.00496429
R28142 VSS.n432 VSS.n277 0.00496429
R28143 VSS.n428 VSS.n280 0.00496429
R28144 VSS.n425 VSS.n280 0.00496429
R28145 VSS.n401 VSS.n304 0.00496429
R28146 VSS.n398 VSS.n178 0.00496429
R28147 VSS.n859 VSS.n480 0.00496429
R28148 VSS.n856 VSS.n486 0.00496429
R28149 VSS.n832 VSS.n509 0.00496429
R28150 VSS.n829 VSS.n509 0.00496429
R28151 VSS.n826 VSS.n515 0.00496429
R28152 VSS.n751 VSS.n750 0.00496429
R28153 VSS.n692 VSS.n691 0.00496429
R28154 VSS.n752 VSS.n713 0.00496429
R28155 VSS.n997 VSS.n443 0.00496429
R28156 VSS.n993 VSS.n446 0.00496429
R28157 VSS.n990 VSS.n446 0.00496429
R28158 VSS.n966 VSS.n470 0.00496429
R28159 VSS.n963 VSS.n476 0.00496429
R28160 VSS.n8360 VSS.n8359 0.00496429
R28161 VSS.n7268 VSS.n7267 0.00496429
R28162 VSS.n8361 VSS.n7289 0.00496429
R28163 VSS.n8508 VSS.n1017 0.00486429
R28164 VSS.n8501 VSS.n1025 0.00486429
R28165 VSS.n8500 VSS.n1026 0.00486429
R28166 VSS.n8493 VSS.n1034 0.00486429
R28167 VSS.n7521 VSS.n7520 0.00486429
R28168 VSS.n7538 VSS.n7445 0.00486429
R28169 VSS.n7540 VSS.n7539 0.00486429
R28170 VSS.n7547 VSS.n7440 0.00486429
R28171 VSS.n8018 VSS.n8017 0.00486429
R28172 VSS.n8025 VSS.n7945 0.00486429
R28173 VSS.n8029 VSS.n8028 0.00486429
R28174 VSS.n8048 VSS.n7922 0.00486429
R28175 VSS.n8113 VSS.n8112 0.00486429
R28176 VSS.n8130 VSS.n7859 0.00486429
R28177 VSS.n8132 VSS.n8131 0.00486429
R28178 VSS.n8139 VSS.n7854 0.00486429
R28179 VSS.n8579 VSS.n8578 0.00486429
R28180 VSS.n8586 VSS.n242 0.00486429
R28181 VSS.n8590 VSS.n8589 0.00486429
R28182 VSS.n8609 VSS.n219 0.00486429
R28183 VSS.n9032 VSS.n8648 0.00486429
R28184 VSS.n9025 VSS.n8656 0.00486429
R28185 VSS.n9024 VSS.n8657 0.00486429
R28186 VSS.n9017 VSS.n8664 0.00486429
R28187 VSS.n1261 VSS.n1260 0.00486429
R28188 VSS.n1268 VSS.n1188 0.00486429
R28189 VSS.n1272 VSS.n1271 0.00486429
R28190 VSS.n1291 VSS.n1165 0.00486429
R28191 VSS.n1695 VSS.n1330 0.00486429
R28192 VSS.n1688 VSS.n1338 0.00486429
R28193 VSS.n1687 VSS.n1339 0.00486429
R28194 VSS.n1680 VSS.n1346 0.00486429
R28195 VSS.n1834 VSS.n1833 0.00486429
R28196 VSS.n1841 VSS.n1761 0.00486429
R28197 VSS.n1845 VSS.n1844 0.00486429
R28198 VSS.n1864 VSS.n1738 0.00486429
R28199 VSS.n2287 VSS.n1903 0.00486429
R28200 VSS.n2280 VSS.n1911 0.00486429
R28201 VSS.n2279 VSS.n1912 0.00486429
R28202 VSS.n2272 VSS.n1919 0.00486429
R28203 VSS.n3628 VSS.n3627 0.00486429
R28204 VSS.n3635 VSS.n3555 0.00486429
R28205 VSS.n3639 VSS.n3638 0.00486429
R28206 VSS.n3658 VSS.n3532 0.00486429
R28207 VSS.n3723 VSS.n3722 0.00486429
R28208 VSS.n3740 VSS.n3469 0.00486429
R28209 VSS.n3742 VSS.n3741 0.00486429
R28210 VSS.n3749 VSS.n3464 0.00486429
R28211 VSS.n4220 VSS.n4219 0.00486429
R28212 VSS.n4227 VSS.n4147 0.00486429
R28213 VSS.n4231 VSS.n4230 0.00486429
R28214 VSS.n4250 VSS.n4124 0.00486429
R28215 VSS.n4315 VSS.n4314 0.00486429
R28216 VSS.n4332 VSS.n4061 0.00486429
R28217 VSS.n4334 VSS.n4333 0.00486429
R28218 VSS.n4341 VSS.n4056 0.00486429
R28219 VSS.n4812 VSS.n4811 0.00486429
R28220 VSS.n4819 VSS.n4739 0.00486429
R28221 VSS.n4823 VSS.n4822 0.00486429
R28222 VSS.n4842 VSS.n4716 0.00486429
R28223 VSS.n4907 VSS.n4906 0.00486429
R28224 VSS.n4924 VSS.n4653 0.00486429
R28225 VSS.n4926 VSS.n4925 0.00486429
R28226 VSS.n4933 VSS.n4648 0.00486429
R28227 VSS.n5404 VSS.n5403 0.00486429
R28228 VSS.n5411 VSS.n5331 0.00486429
R28229 VSS.n5415 VSS.n5414 0.00486429
R28230 VSS.n5434 VSS.n5308 0.00486429
R28231 VSS.n5499 VSS.n5498 0.00486429
R28232 VSS.n5516 VSS.n5245 0.00486429
R28233 VSS.n5518 VSS.n5517 0.00486429
R28234 VSS.n5525 VSS.n5240 0.00486429
R28235 VSS.n5996 VSS.n5995 0.00486429
R28236 VSS.n6003 VSS.n5923 0.00486429
R28237 VSS.n6007 VSS.n6006 0.00486429
R28238 VSS.n6026 VSS.n5900 0.00486429
R28239 VSS.n6091 VSS.n6090 0.00486429
R28240 VSS.n6108 VSS.n5837 0.00486429
R28241 VSS.n6110 VSS.n6109 0.00486429
R28242 VSS.n6117 VSS.n5832 0.00486429
R28243 VSS.n6588 VSS.n6587 0.00486429
R28244 VSS.n6595 VSS.n6515 0.00486429
R28245 VSS.n6599 VSS.n6598 0.00486429
R28246 VSS.n6618 VSS.n6492 0.00486429
R28247 VSS.n6683 VSS.n6682 0.00486429
R28248 VSS.n6700 VSS.n6429 0.00486429
R28249 VSS.n6702 VSS.n6701 0.00486429
R28250 VSS.n6709 VSS.n6424 0.00486429
R28251 VSS.n2432 VSS.n2431 0.00486429
R28252 VSS.n2439 VSS.n2359 0.00486429
R28253 VSS.n2443 VSS.n2442 0.00486429
R28254 VSS.n2462 VSS.n2336 0.00486429
R28255 VSS.n7031 VSS.n2501 0.00486429
R28256 VSS.n7024 VSS.n2509 0.00486429
R28257 VSS.n7023 VSS.n2510 0.00486429
R28258 VSS.n7016 VSS.n2517 0.00486429
R28259 VSS.n3026 VSS.n3025 0.00486429
R28260 VSS.n3043 VSS.n2951 0.00486429
R28261 VSS.n3045 VSS.n3044 0.00486429
R28262 VSS.n3052 VSS.n2946 0.00486429
R28263 VSS.n3131 VSS.n3130 0.00486429
R28264 VSS.n3148 VSS.n2876 0.00486429
R28265 VSS.n3150 VSS.n3149 0.00486429
R28266 VSS.n3157 VSS.n2871 0.00486429
R28267 VSS.n422 VSS.n284 0.00486429
R28268 VSS.n415 VSS.n292 0.00486429
R28269 VSS.n414 VSS.n293 0.00486429
R28270 VSS.n407 VSS.n301 0.00486429
R28271 VSS.n9091 VSS.n9090 0.00486429
R28272 VSS.n9108 VSS.n143 0.00486429
R28273 VSS.n9110 VSS.n9109 0.00486429
R28274 VSS.n9117 VSS.n138 0.00486429
R28275 VSS.n987 VSS.n450 0.00486429
R28276 VSS.n980 VSS.n458 0.00486429
R28277 VSS.n979 VSS.n459 0.00486429
R28278 VSS.n972 VSS.n467 0.00486429
R28279 VSS.n850 VSS.n490 0.00486429
R28280 VSS.n843 VSS.n498 0.00486429
R28281 VSS.n842 VSS.n499 0.00486429
R28282 VSS.n835 VSS.n506 0.00486429
R28283 VSS.n8459 VSS.n7069 0.00486429
R28284 VSS.n8452 VSS.n7077 0.00486429
R28285 VSS.n8451 VSS.n7078 0.00486429
R28286 VSS.n8444 VSS.n7085 0.00486429
R28287 VSS.n7751 VSS 0.00452857
R28288 VSS.n8343 VSS 0.00452857
R28289 VSS.n8892 VSS 0.00452857
R28290 VSS.n9351 VSS 0.00452857
R28291 VSS.n2173 VSS 0.00452857
R28292 VSS.n3954 VSS 0.00452857
R28293 VSS.n4546 VSS 0.00452857
R28294 VSS.n5138 VSS 0.00452857
R28295 VSS.n5730 VSS 0.00452857
R28296 VSS.n6322 VSS 0.00452857
R28297 VSS.n6914 VSS 0.00452857
R28298 VSS.n6917 VSS 0.00452857
R28299 VSS.n3362 VSS 0.00452857
R28300 VSS.n9322 VSS 0.00452857
R28301 VSS.n9324 VSS 0.00452857
R28302 VSS.n8345 VSS 0.00452857
R28303 VSS.n908 VSS.n448 0.00407143
R28304 VSS.n1089 VSS.n1015 0.00407143
R28305 VSS.n7587 VSS.n7409 0.00407143
R28306 VSS.n7628 VSS.n7403 0.00407143
R28307 VSS.n7634 VSS.n7633 0.00407143
R28308 VSS.n7748 VSS.n7342 0.00407143
R28309 VSS.n7627 VSS.n7626 0.00407143
R28310 VSS.n7635 VSS.n7399 0.00407143
R28311 VSS.n7689 VSS.n7688 0.00407143
R28312 VSS.n7965 VSS.n7952 0.00407143
R28313 VSS.n8179 VSS.n7823 0.00407143
R28314 VSS.n8220 VSS.n7817 0.00407143
R28315 VSS.n8226 VSS.n8225 0.00407143
R28316 VSS.n8340 VSS.n7756 0.00407143
R28317 VSS.n8219 VSS.n8218 0.00407143
R28318 VSS.n8227 VSS.n7813 0.00407143
R28319 VSS.n8281 VSS.n8280 0.00407143
R28320 VSS.n262 VSS.n249 0.00407143
R28321 VSS.n8788 VSS.n8786 0.00407143
R28322 VSS.n8988 VSS.n8779 0.00407143
R28323 VSS.n8981 VSS.n8980 0.00407143
R28324 VSS.n8928 VSS.n8897 0.00407143
R28325 VSS.n8987 VSS.n8986 0.00407143
R28326 VSS.n8982 VSS.n8801 0.00407143
R28327 VSS.n8863 VSS.n8862 0.00407143
R28328 VSS.n1208 VSS.n1195 0.00407143
R28329 VSS.n1469 VSS.n1467 0.00407143
R28330 VSS.n1648 VSS.n1460 0.00407143
R28331 VSS.n1495 VSS.n1494 0.00407143
R28332 VSS.n9348 VSS.n4 0.00407143
R28333 VSS.n1650 VSS.n1649 0.00407143
R28334 VSS.n1496 VSS.n1493 0.00407143
R28335 VSS.n1619 VSS.n1618 0.00407143
R28336 VSS.n1781 VSS.n1768 0.00407143
R28337 VSS.n2042 VSS.n2040 0.00407143
R28338 VSS.n2240 VSS.n2033 0.00407143
R28339 VSS.n2068 VSS.n2067 0.00407143
R28340 VSS.n2177 VSS.n2176 0.00407143
R28341 VSS.n2242 VSS.n2241 0.00407143
R28342 VSS.n2069 VSS.n2066 0.00407143
R28343 VSS.n2211 VSS.n2210 0.00407143
R28344 VSS.n3575 VSS.n3562 0.00407143
R28345 VSS.n3789 VSS.n3433 0.00407143
R28346 VSS.n3830 VSS.n3427 0.00407143
R28347 VSS.n3836 VSS.n3835 0.00407143
R28348 VSS.n3951 VSS.n3367 0.00407143
R28349 VSS.n3829 VSS.n3828 0.00407143
R28350 VSS.n3837 VSS.n3423 0.00407143
R28351 VSS.n3891 VSS.n3890 0.00407143
R28352 VSS.n4167 VSS.n4154 0.00407143
R28353 VSS.n4381 VSS.n4025 0.00407143
R28354 VSS.n4422 VSS.n4019 0.00407143
R28355 VSS.n4428 VSS.n4427 0.00407143
R28356 VSS.n4543 VSS.n3959 0.00407143
R28357 VSS.n4421 VSS.n4420 0.00407143
R28358 VSS.n4429 VSS.n4015 0.00407143
R28359 VSS.n4483 VSS.n4482 0.00407143
R28360 VSS.n4759 VSS.n4746 0.00407143
R28361 VSS.n4973 VSS.n4617 0.00407143
R28362 VSS.n5014 VSS.n4611 0.00407143
R28363 VSS.n5020 VSS.n5019 0.00407143
R28364 VSS.n5135 VSS.n4551 0.00407143
R28365 VSS.n5013 VSS.n5012 0.00407143
R28366 VSS.n5021 VSS.n4607 0.00407143
R28367 VSS.n5075 VSS.n5074 0.00407143
R28368 VSS.n5351 VSS.n5338 0.00407143
R28369 VSS.n5565 VSS.n5209 0.00407143
R28370 VSS.n5606 VSS.n5203 0.00407143
R28371 VSS.n5612 VSS.n5611 0.00407143
R28372 VSS.n5727 VSS.n5143 0.00407143
R28373 VSS.n5605 VSS.n5604 0.00407143
R28374 VSS.n5613 VSS.n5199 0.00407143
R28375 VSS.n5667 VSS.n5666 0.00407143
R28376 VSS.n5943 VSS.n5930 0.00407143
R28377 VSS.n6157 VSS.n5801 0.00407143
R28378 VSS.n6198 VSS.n5795 0.00407143
R28379 VSS.n6204 VSS.n6203 0.00407143
R28380 VSS.n6319 VSS.n5735 0.00407143
R28381 VSS.n6197 VSS.n6196 0.00407143
R28382 VSS.n6205 VSS.n5791 0.00407143
R28383 VSS.n6259 VSS.n6258 0.00407143
R28384 VSS.n6535 VSS.n6522 0.00407143
R28385 VSS.n6749 VSS.n6393 0.00407143
R28386 VSS.n6790 VSS.n6387 0.00407143
R28387 VSS.n6796 VSS.n6795 0.00407143
R28388 VSS.n6911 VSS.n6327 0.00407143
R28389 VSS.n6789 VSS.n6788 0.00407143
R28390 VSS.n6797 VSS.n6383 0.00407143
R28391 VSS.n6851 VSS.n6850 0.00407143
R28392 VSS.n2379 VSS.n2366 0.00407143
R28393 VSS.n2640 VSS.n2638 0.00407143
R28394 VSS.n6984 VSS.n2631 0.00407143
R28395 VSS.n2666 VSS.n2665 0.00407143
R28396 VSS.n6921 VSS.n6920 0.00407143
R28397 VSS.n6986 VSS.n6985 0.00407143
R28398 VSS.n2667 VSS.n2664 0.00407143
R28399 VSS.n6955 VSS.n6954 0.00407143
R28400 VSS.n3018 VSS.n2971 0.00407143
R28401 VSS.n3197 VSS.n2840 0.00407143
R28402 VSS.n3238 VSS.n2834 0.00407143
R28403 VSS.n3244 VSS.n3243 0.00407143
R28404 VSS.n3359 VSS.n2774 0.00407143
R28405 VSS.n3237 VSS.n3236 0.00407143
R28406 VSS.n3245 VSS.n2830 0.00407143
R28407 VSS.n3299 VSS.n3298 0.00407143
R28408 VSS.n350 VSS.n282 0.00407143
R28409 VSS.n9157 VSS.n107 0.00407143
R28410 VSS.n9198 VSS.n101 0.00407143
R28411 VSS.n9204 VSS.n9203 0.00407143
R28412 VSS.n9319 VSS.n41 0.00407143
R28413 VSS.n9197 VSS.n9196 0.00407143
R28414 VSS.n9205 VSS.n97 0.00407143
R28415 VSS.n9259 VSS.n9258 0.00407143
R28416 VSS.n632 VSS.n630 0.00407143
R28417 VSS.n803 VSS.n623 0.00407143
R28418 VSS.n658 VSS.n657 0.00407143
R28419 VSS.n9328 VSS.n9327 0.00407143
R28420 VSS.n805 VSS.n804 0.00407143
R28421 VSS.n659 VSS.n656 0.00407143
R28422 VSS.n774 VSS.n773 0.00407143
R28423 VSS.n7208 VSS.n7206 0.00407143
R28424 VSS.n8412 VSS.n7199 0.00407143
R28425 VSS.n7234 VSS.n7233 0.00407143
R28426 VSS.n8349 VSS.n8348 0.00407143
R28427 VSS.n8414 VSS.n8413 0.00407143
R28428 VSS.n7235 VSS.n7232 0.00407143
R28429 VSS.n8383 VSS.n8382 0.00407143
R28430 VSS.n7614 VSS.n7613 0.00352143
R28431 VSS.n7623 VSS.n7406 0.00352143
R28432 VSS.n7654 VSS.n7653 0.00352143
R28433 VSS.n7655 VSS.n7380 0.00352143
R28434 VSS.n7686 VSS.n7671 0.00352143
R28435 VSS.n7705 VSS.n7366 0.00352143
R28436 VSS.n7726 VSS.n7725 0.00352143
R28437 VSS.n7750 VSS.n7339 0.00352143
R28438 VSS.n8206 VSS.n8205 0.00352143
R28439 VSS.n8215 VSS.n7820 0.00352143
R28440 VSS.n8246 VSS.n8245 0.00352143
R28441 VSS.n8247 VSS.n7794 0.00352143
R28442 VSS.n8278 VSS.n8263 0.00352143
R28443 VSS.n8297 VSS.n7780 0.00352143
R28444 VSS.n8318 VSS.n8317 0.00352143
R28445 VSS.n8342 VSS.n7753 0.00352143
R28446 VSS.n8792 VSS.n8791 0.00352143
R28447 VSS.n8799 VSS.n8781 0.00352143
R28448 VSS.n8813 VSS.n8800 0.00352143
R28449 VSS.n8967 VSS.n8814 0.00352143
R28450 VSS.n8876 VSS.n8855 0.00352143
R28451 VSS.n8949 VSS.n8877 0.00352143
R28452 VSS.n8933 VSS.n8932 0.00352143
R28453 VSS.n8931 VSS.n8893 0.00352143
R28454 VSS.n1473 VSS.n1472 0.00352143
R28455 VSS.n1480 VSS.n1463 0.00352143
R28456 VSS.n1515 VSS.n1498 0.00352143
R28457 VSS.n1516 VSS.n1511 0.00352143
R28458 VSS.n1616 VSS.n1532 0.00352143
R28459 VSS.n1548 VSS.n1547 0.00352143
R28460 VSS.n1554 VSS.n1549 0.00352143
R28461 VSS.n9350 VSS.n1 0.00352143
R28462 VSS.n2046 VSS.n2045 0.00352143
R28463 VSS.n2053 VSS.n2036 0.00352143
R28464 VSS.n2088 VSS.n2071 0.00352143
R28465 VSS.n2089 VSS.n2084 0.00352143
R28466 VSS.n2208 VSS.n2105 0.00352143
R28467 VSS.n2121 VSS.n2120 0.00352143
R28468 VSS.n2171 VSS.n2122 0.00352143
R28469 VSS.n2174 VSS.n2172 0.00352143
R28470 VSS.n3816 VSS.n3815 0.00352143
R28471 VSS.n3825 VSS.n3430 0.00352143
R28472 VSS.n3856 VSS.n3855 0.00352143
R28473 VSS.n3857 VSS.n3404 0.00352143
R28474 VSS.n3888 VSS.n3873 0.00352143
R28475 VSS.n3907 VSS.n3390 0.00352143
R28476 VSS.n3928 VSS.n3927 0.00352143
R28477 VSS.n3953 VSS.n3364 0.00352143
R28478 VSS.n4408 VSS.n4407 0.00352143
R28479 VSS.n4417 VSS.n4022 0.00352143
R28480 VSS.n4448 VSS.n4447 0.00352143
R28481 VSS.n4449 VSS.n3996 0.00352143
R28482 VSS.n4480 VSS.n4465 0.00352143
R28483 VSS.n4499 VSS.n3982 0.00352143
R28484 VSS.n4520 VSS.n4519 0.00352143
R28485 VSS.n4545 VSS.n3956 0.00352143
R28486 VSS.n5000 VSS.n4999 0.00352143
R28487 VSS.n5009 VSS.n4614 0.00352143
R28488 VSS.n5040 VSS.n5039 0.00352143
R28489 VSS.n5041 VSS.n4588 0.00352143
R28490 VSS.n5072 VSS.n5057 0.00352143
R28491 VSS.n5091 VSS.n4574 0.00352143
R28492 VSS.n5112 VSS.n5111 0.00352143
R28493 VSS.n5137 VSS.n4548 0.00352143
R28494 VSS.n5592 VSS.n5591 0.00352143
R28495 VSS.n5601 VSS.n5206 0.00352143
R28496 VSS.n5632 VSS.n5631 0.00352143
R28497 VSS.n5633 VSS.n5180 0.00352143
R28498 VSS.n5664 VSS.n5649 0.00352143
R28499 VSS.n5683 VSS.n5166 0.00352143
R28500 VSS.n5704 VSS.n5703 0.00352143
R28501 VSS.n5729 VSS.n5140 0.00352143
R28502 VSS.n6184 VSS.n6183 0.00352143
R28503 VSS.n6193 VSS.n5798 0.00352143
R28504 VSS.n6224 VSS.n6223 0.00352143
R28505 VSS.n6225 VSS.n5772 0.00352143
R28506 VSS.n6256 VSS.n6241 0.00352143
R28507 VSS.n6275 VSS.n5758 0.00352143
R28508 VSS.n6296 VSS.n6295 0.00352143
R28509 VSS.n6321 VSS.n5732 0.00352143
R28510 VSS.n6776 VSS.n6775 0.00352143
R28511 VSS.n6785 VSS.n6390 0.00352143
R28512 VSS.n6816 VSS.n6815 0.00352143
R28513 VSS.n6817 VSS.n6364 0.00352143
R28514 VSS.n6848 VSS.n6833 0.00352143
R28515 VSS.n6867 VSS.n6350 0.00352143
R28516 VSS.n6888 VSS.n6887 0.00352143
R28517 VSS.n6913 VSS.n6324 0.00352143
R28518 VSS.n2644 VSS.n2643 0.00352143
R28519 VSS.n2651 VSS.n2634 0.00352143
R28520 VSS.n2686 VSS.n2669 0.00352143
R28521 VSS.n2687 VSS.n2682 0.00352143
R28522 VSS.n6952 VSS.n2703 0.00352143
R28523 VSS.n2719 VSS.n2718 0.00352143
R28524 VSS.n2769 VSS.n2720 0.00352143
R28525 VSS.n6918 VSS.n2770 0.00352143
R28526 VSS.n3224 VSS.n3223 0.00352143
R28527 VSS.n3233 VSS.n2837 0.00352143
R28528 VSS.n3264 VSS.n3263 0.00352143
R28529 VSS.n3265 VSS.n2811 0.00352143
R28530 VSS.n3296 VSS.n3281 0.00352143
R28531 VSS.n3315 VSS.n2797 0.00352143
R28532 VSS.n3336 VSS.n3335 0.00352143
R28533 VSS.n3361 VSS.n2771 0.00352143
R28534 VSS.n9184 VSS.n9183 0.00352143
R28535 VSS.n9193 VSS.n104 0.00352143
R28536 VSS.n9224 VSS.n9223 0.00352143
R28537 VSS.n9225 VSS.n78 0.00352143
R28538 VSS.n9256 VSS.n9241 0.00352143
R28539 VSS.n9275 VSS.n64 0.00352143
R28540 VSS.n9296 VSS.n9295 0.00352143
R28541 VSS.n9321 VSS.n38 0.00352143
R28542 VSS.n636 VSS.n635 0.00352143
R28543 VSS.n643 VSS.n626 0.00352143
R28544 VSS.n678 VSS.n661 0.00352143
R28545 VSS.n679 VSS.n674 0.00352143
R28546 VSS.n771 VSS.n695 0.00352143
R28547 VSS.n711 VSS.n710 0.00352143
R28548 VSS.n717 VSS.n712 0.00352143
R28549 VSS.n9325 VSS.n36 0.00352143
R28550 VSS.n7212 VSS.n7211 0.00352143
R28551 VSS.n7219 VSS.n7202 0.00352143
R28552 VSS.n7254 VSS.n7237 0.00352143
R28553 VSS.n7255 VSS.n7250 0.00352143
R28554 VSS.n8380 VSS.n7271 0.00352143
R28555 VSS.n7287 VSS.n7286 0.00352143
R28556 VSS.n7337 VSS.n7288 0.00352143
R28557 VSS.n8346 VSS.n7338 0.00352143
R28558 VSS.n1025 VSS.n1017 0.00318571
R28559 VSS.n1034 VSS.n1026 0.00318571
R28560 VSS.n7520 VSS.n7445 0.00318571
R28561 VSS.n7540 VSS.n7440 0.00318571
R28562 VSS.n8018 VSS.n7945 0.00318571
R28563 VSS.n8028 VSS.n7922 0.00318571
R28564 VSS.n8112 VSS.n7859 0.00318571
R28565 VSS.n8132 VSS.n7854 0.00318571
R28566 VSS.n8579 VSS.n242 0.00318571
R28567 VSS.n8589 VSS.n219 0.00318571
R28568 VSS.n8656 VSS.n8648 0.00318571
R28569 VSS.n8664 VSS.n8657 0.00318571
R28570 VSS.n1261 VSS.n1188 0.00318571
R28571 VSS.n1271 VSS.n1165 0.00318571
R28572 VSS.n1338 VSS.n1330 0.00318571
R28573 VSS.n1346 VSS.n1339 0.00318571
R28574 VSS.n1834 VSS.n1761 0.00318571
R28575 VSS.n1844 VSS.n1738 0.00318571
R28576 VSS.n1911 VSS.n1903 0.00318571
R28577 VSS.n1919 VSS.n1912 0.00318571
R28578 VSS.n3628 VSS.n3555 0.00318571
R28579 VSS.n3638 VSS.n3532 0.00318571
R28580 VSS.n3722 VSS.n3469 0.00318571
R28581 VSS.n3742 VSS.n3464 0.00318571
R28582 VSS.n4220 VSS.n4147 0.00318571
R28583 VSS.n4230 VSS.n4124 0.00318571
R28584 VSS.n4314 VSS.n4061 0.00318571
R28585 VSS.n4334 VSS.n4056 0.00318571
R28586 VSS.n4812 VSS.n4739 0.00318571
R28587 VSS.n4822 VSS.n4716 0.00318571
R28588 VSS.n4906 VSS.n4653 0.00318571
R28589 VSS.n4926 VSS.n4648 0.00318571
R28590 VSS.n5404 VSS.n5331 0.00318571
R28591 VSS.n5414 VSS.n5308 0.00318571
R28592 VSS.n5498 VSS.n5245 0.00318571
R28593 VSS.n5518 VSS.n5240 0.00318571
R28594 VSS.n5996 VSS.n5923 0.00318571
R28595 VSS.n6006 VSS.n5900 0.00318571
R28596 VSS.n6090 VSS.n5837 0.00318571
R28597 VSS.n6110 VSS.n5832 0.00318571
R28598 VSS.n6588 VSS.n6515 0.00318571
R28599 VSS.n6598 VSS.n6492 0.00318571
R28600 VSS.n6682 VSS.n6429 0.00318571
R28601 VSS.n6702 VSS.n6424 0.00318571
R28602 VSS.n2432 VSS.n2359 0.00318571
R28603 VSS.n2442 VSS.n2336 0.00318571
R28604 VSS.n2509 VSS.n2501 0.00318571
R28605 VSS.n2517 VSS.n2510 0.00318571
R28606 VSS.n3025 VSS.n2951 0.00318571
R28607 VSS.n3045 VSS.n2946 0.00318571
R28608 VSS.n3130 VSS.n2876 0.00318571
R28609 VSS.n3150 VSS.n2871 0.00318571
R28610 VSS.n292 VSS.n284 0.00318571
R28611 VSS.n301 VSS.n293 0.00318571
R28612 VSS.n9090 VSS.n143 0.00318571
R28613 VSS.n9110 VSS.n138 0.00318571
R28614 VSS.n458 VSS.n450 0.00318571
R28615 VSS.n467 VSS.n459 0.00318571
R28616 VSS.n498 VSS.n490 0.00318571
R28617 VSS.n506 VSS.n499 0.00318571
R28618 VSS.n7077 VSS.n7069 0.00318571
R28619 VSS.n7085 VSS.n7078 0.00318571
R28620 VSS.n7127 VSS.n7060 0.00317857
R28621 VSS.n8464 VSS.n7066 0.00317857
R28622 VSS.n8449 VSS.n8448 0.00317857
R28623 VSS.n7163 VSS.n7089 0.00317857
R28624 VSS.n8439 VSS.n7090 0.00317857
R28625 VSS.n8434 VSS.n7095 0.00317857
R28626 VSS.n7126 VSS.n7062 0.00317857
R28627 VSS.n8465 VSS.n7064 0.00317857
R28628 VSS.n8450 VSS.n7079 0.00317857
R28629 VSS.n8438 VSS.n7091 0.00317857
R28630 VSS.n8435 VSS.n7093 0.00317857
R28631 VSS.n896 VSS.n441 0.00317857
R28632 VSS.n992 VSS.n447 0.00317857
R28633 VSS.n983 VSS.n454 0.00317857
R28634 VSS.n930 VSS.n471 0.00317857
R28635 VSS.n967 VSS.n472 0.00317857
R28636 VSS.n962 VSS.n477 0.00317857
R28637 VSS.n7497 VSS.n7496 0.00317857
R28638 VSS.n7503 VSS.n7473 0.00317857
R28639 VSS.n7543 VSS.n7442 0.00317857
R28640 VSS.n7552 VSS.n7551 0.00317857
R28641 VSS.n7568 VSS.n7567 0.00317857
R28642 VSS.n7573 VSS.n7413 0.00317857
R28643 VSS.n1077 VSS.n1008 0.00317857
R28644 VSS.n8513 VSS.n1014 0.00317857
R28645 VSS.n8504 VSS.n1021 0.00317857
R28646 VSS.n1111 VSS.n1038 0.00317857
R28647 VSS.n8488 VSS.n1039 0.00317857
R28648 VSS.n8483 VSS.n1044 0.00317857
R28649 VSS.n1076 VSS.n1010 0.00317857
R28650 VSS.n8514 VSS.n1012 0.00317857
R28651 VSS.n8503 VSS.n8502 0.00317857
R28652 VSS.n8487 VSS.n1040 0.00317857
R28653 VSS.n8484 VSS.n1042 0.00317857
R28654 VSS.n7588 VSS.n7587 0.00317857
R28655 VSS.n7665 VSS.n7382 0.00317857
R28656 VSS.n7677 VSS.n7377 0.00317857
R28657 VSS.n7707 VSS.n7364 0.00317857
R28658 VSS.n7730 VSS.n7729 0.00317857
R28659 VSS.n7748 VSS.n7747 0.00317857
R28660 VSS.n7709 VSS.n7708 0.00317857
R28661 VSS.n7498 VSS.n7477 0.00317857
R28662 VSS.n7502 VSS.n7501 0.00317857
R28663 VSS.n7542 VSS.n7443 0.00317857
R28664 VSS.n7569 VSS.n7425 0.00317857
R28665 VSS.n7574 VSS.n7572 0.00317857
R28666 VSS.n8089 VSS.n8088 0.00317857
R28667 VSS.n8095 VSS.n7887 0.00317857
R28668 VSS.n8135 VSS.n7856 0.00317857
R28669 VSS.n8144 VSS.n8143 0.00317857
R28670 VSS.n8160 VSS.n8159 0.00317857
R28671 VSS.n8165 VSS.n7827 0.00317857
R28672 VSS.n7991 VSS.n7990 0.00317857
R28673 VSS.n7997 VSS.n7967 0.00317857
R28674 VSS.n8022 VSS.n7940 0.00317857
R28675 VSS.n7933 VSS.n7920 0.00317857
R28676 VSS.n8053 VSS.n7909 0.00317857
R28677 VSS.n8059 VSS.n7902 0.00317857
R28678 VSS.n7992 VSS.n7971 0.00317857
R28679 VSS.n7996 VSS.n7995 0.00317857
R28680 VSS.n8024 VSS.n8023 0.00317857
R28681 VSS.n8054 VSS.n7911 0.00317857
R28682 VSS.n8058 VSS.n8057 0.00317857
R28683 VSS.n8180 VSS.n8179 0.00317857
R28684 VSS.n8257 VSS.n7796 0.00317857
R28685 VSS.n8269 VSS.n7791 0.00317857
R28686 VSS.n8299 VSS.n7778 0.00317857
R28687 VSS.n8322 VSS.n8321 0.00317857
R28688 VSS.n8340 VSS.n8339 0.00317857
R28689 VSS.n8301 VSS.n8300 0.00317857
R28690 VSS.n8090 VSS.n7891 0.00317857
R28691 VSS.n8094 VSS.n8093 0.00317857
R28692 VSS.n8134 VSS.n7857 0.00317857
R28693 VSS.n8161 VSS.n7839 0.00317857
R28694 VSS.n8166 VSS.n8164 0.00317857
R28695 VSS.n8552 VSS.n8551 0.00317857
R28696 VSS.n8558 VSS.n264 0.00317857
R28697 VSS.n8583 VSS.n237 0.00317857
R28698 VSS.n230 VSS.n217 0.00317857
R28699 VSS.n8614 VSS.n206 0.00317857
R28700 VSS.n8620 VSS.n199 0.00317857
R28701 VSS.n8706 VSS.n196 0.00317857
R28702 VSS.n9037 VSS.n8645 0.00317857
R28703 VSS.n9022 VSS.n9021 0.00317857
R28704 VSS.n8742 VSS.n8668 0.00317857
R28705 VSS.n9012 VSS.n8669 0.00317857
R28706 VSS.n9007 VSS.n8674 0.00317857
R28707 VSS.n8705 VSS.n8641 0.00317857
R28708 VSS.n9038 VSS.n8643 0.00317857
R28709 VSS.n9023 VSS.n8658 0.00317857
R28710 VSS.n9011 VSS.n8670 0.00317857
R28711 VSS.n9008 VSS.n8672 0.00317857
R28712 VSS.n8788 VSS.n8787 0.00317857
R28713 VSS.n8839 VSS.n8818 0.00317857
R28714 VSS.n8866 VSS.n8865 0.00317857
R28715 VSS.n8946 VSS.n8881 0.00317857
R28716 VSS.n8935 VSS.n8889 0.00317857
R28717 VSS.n8928 VSS.n8927 0.00317857
R28718 VSS.n8947 VSS.n8879 0.00317857
R28719 VSS.n8553 VSS.n268 0.00317857
R28720 VSS.n8557 VSS.n8556 0.00317857
R28721 VSS.n8585 VSS.n8584 0.00317857
R28722 VSS.n8615 VSS.n208 0.00317857
R28723 VSS.n8619 VSS.n8618 0.00317857
R28724 VSS.n1234 VSS.n1233 0.00317857
R28725 VSS.n1240 VSS.n1210 0.00317857
R28726 VSS.n1265 VSS.n1183 0.00317857
R28727 VSS.n1176 VSS.n1163 0.00317857
R28728 VSS.n1296 VSS.n1152 0.00317857
R28729 VSS.n1302 VSS.n1145 0.00317857
R28730 VSS.n1388 VSS.n1142 0.00317857
R28731 VSS.n1700 VSS.n1327 0.00317857
R28732 VSS.n1685 VSS.n1684 0.00317857
R28733 VSS.n1424 VSS.n1350 0.00317857
R28734 VSS.n1675 VSS.n1351 0.00317857
R28735 VSS.n1670 VSS.n1356 0.00317857
R28736 VSS.n1387 VSS.n1323 0.00317857
R28737 VSS.n1701 VSS.n1325 0.00317857
R28738 VSS.n1686 VSS.n1340 0.00317857
R28739 VSS.n1674 VSS.n1352 0.00317857
R28740 VSS.n1671 VSS.n1354 0.00317857
R28741 VSS.n1469 VSS.n1468 0.00317857
R28742 VSS.n1526 VSS.n1513 0.00317857
R28743 VSS.n1573 VSS.n1508 0.00317857
R28744 VSS.n1603 VSS.n1602 0.00317857
R28745 VSS.n1559 VSS.n1558 0.00317857
R28746 VSS.n9348 VSS.n9347 0.00317857
R28747 VSS.n1601 VSS.n1541 0.00317857
R28748 VSS.n1235 VSS.n1214 0.00317857
R28749 VSS.n1239 VSS.n1238 0.00317857
R28750 VSS.n1267 VSS.n1266 0.00317857
R28751 VSS.n1297 VSS.n1154 0.00317857
R28752 VSS.n1301 VSS.n1300 0.00317857
R28753 VSS.n1807 VSS.n1806 0.00317857
R28754 VSS.n1813 VSS.n1783 0.00317857
R28755 VSS.n1838 VSS.n1756 0.00317857
R28756 VSS.n1749 VSS.n1736 0.00317857
R28757 VSS.n1869 VSS.n1725 0.00317857
R28758 VSS.n1875 VSS.n1718 0.00317857
R28759 VSS.n1961 VSS.n1715 0.00317857
R28760 VSS.n2292 VSS.n1900 0.00317857
R28761 VSS.n2277 VSS.n2276 0.00317857
R28762 VSS.n1997 VSS.n1923 0.00317857
R28763 VSS.n2267 VSS.n1924 0.00317857
R28764 VSS.n2262 VSS.n1929 0.00317857
R28765 VSS.n1960 VSS.n1896 0.00317857
R28766 VSS.n2293 VSS.n1898 0.00317857
R28767 VSS.n2278 VSS.n1913 0.00317857
R28768 VSS.n2266 VSS.n1925 0.00317857
R28769 VSS.n2263 VSS.n1927 0.00317857
R28770 VSS.n2042 VSS.n2041 0.00317857
R28771 VSS.n2099 VSS.n2086 0.00317857
R28772 VSS.n2133 VSS.n2081 0.00317857
R28773 VSS.n2195 VSS.n2194 0.00317857
R28774 VSS.n2167 VSS.n2166 0.00317857
R28775 VSS.n2176 VSS.n2154 0.00317857
R28776 VSS.n2193 VSS.n2114 0.00317857
R28777 VSS.n1808 VSS.n1787 0.00317857
R28778 VSS.n1812 VSS.n1811 0.00317857
R28779 VSS.n1840 VSS.n1839 0.00317857
R28780 VSS.n1870 VSS.n1727 0.00317857
R28781 VSS.n1874 VSS.n1873 0.00317857
R28782 VSS.n3601 VSS.n3600 0.00317857
R28783 VSS.n3607 VSS.n3577 0.00317857
R28784 VSS.n3632 VSS.n3550 0.00317857
R28785 VSS.n3543 VSS.n3530 0.00317857
R28786 VSS.n3663 VSS.n3519 0.00317857
R28787 VSS.n3669 VSS.n3512 0.00317857
R28788 VSS.n3699 VSS.n3698 0.00317857
R28789 VSS.n3705 VSS.n3497 0.00317857
R28790 VSS.n3745 VSS.n3466 0.00317857
R28791 VSS.n3754 VSS.n3753 0.00317857
R28792 VSS.n3770 VSS.n3769 0.00317857
R28793 VSS.n3775 VSS.n3437 0.00317857
R28794 VSS.n3700 VSS.n3501 0.00317857
R28795 VSS.n3704 VSS.n3703 0.00317857
R28796 VSS.n3744 VSS.n3467 0.00317857
R28797 VSS.n3771 VSS.n3449 0.00317857
R28798 VSS.n3776 VSS.n3774 0.00317857
R28799 VSS.n3790 VSS.n3789 0.00317857
R28800 VSS.n3867 VSS.n3406 0.00317857
R28801 VSS.n3879 VSS.n3401 0.00317857
R28802 VSS.n3909 VSS.n3388 0.00317857
R28803 VSS.n3933 VSS.n3932 0.00317857
R28804 VSS.n3951 VSS.n3950 0.00317857
R28805 VSS.n3911 VSS.n3910 0.00317857
R28806 VSS.n3602 VSS.n3581 0.00317857
R28807 VSS.n3606 VSS.n3605 0.00317857
R28808 VSS.n3634 VSS.n3633 0.00317857
R28809 VSS.n3664 VSS.n3521 0.00317857
R28810 VSS.n3668 VSS.n3667 0.00317857
R28811 VSS.n4193 VSS.n4192 0.00317857
R28812 VSS.n4199 VSS.n4169 0.00317857
R28813 VSS.n4224 VSS.n4142 0.00317857
R28814 VSS.n4135 VSS.n4122 0.00317857
R28815 VSS.n4255 VSS.n4111 0.00317857
R28816 VSS.n4261 VSS.n4104 0.00317857
R28817 VSS.n4291 VSS.n4290 0.00317857
R28818 VSS.n4297 VSS.n4089 0.00317857
R28819 VSS.n4337 VSS.n4058 0.00317857
R28820 VSS.n4346 VSS.n4345 0.00317857
R28821 VSS.n4362 VSS.n4361 0.00317857
R28822 VSS.n4367 VSS.n4029 0.00317857
R28823 VSS.n4292 VSS.n4093 0.00317857
R28824 VSS.n4296 VSS.n4295 0.00317857
R28825 VSS.n4336 VSS.n4059 0.00317857
R28826 VSS.n4363 VSS.n4041 0.00317857
R28827 VSS.n4368 VSS.n4366 0.00317857
R28828 VSS.n4382 VSS.n4381 0.00317857
R28829 VSS.n4459 VSS.n3998 0.00317857
R28830 VSS.n4471 VSS.n3993 0.00317857
R28831 VSS.n4501 VSS.n3980 0.00317857
R28832 VSS.n4525 VSS.n4524 0.00317857
R28833 VSS.n4543 VSS.n4542 0.00317857
R28834 VSS.n4503 VSS.n4502 0.00317857
R28835 VSS.n4194 VSS.n4173 0.00317857
R28836 VSS.n4198 VSS.n4197 0.00317857
R28837 VSS.n4226 VSS.n4225 0.00317857
R28838 VSS.n4256 VSS.n4113 0.00317857
R28839 VSS.n4260 VSS.n4259 0.00317857
R28840 VSS.n4785 VSS.n4784 0.00317857
R28841 VSS.n4791 VSS.n4761 0.00317857
R28842 VSS.n4816 VSS.n4734 0.00317857
R28843 VSS.n4727 VSS.n4714 0.00317857
R28844 VSS.n4847 VSS.n4703 0.00317857
R28845 VSS.n4853 VSS.n4696 0.00317857
R28846 VSS.n4883 VSS.n4882 0.00317857
R28847 VSS.n4889 VSS.n4681 0.00317857
R28848 VSS.n4929 VSS.n4650 0.00317857
R28849 VSS.n4938 VSS.n4937 0.00317857
R28850 VSS.n4954 VSS.n4953 0.00317857
R28851 VSS.n4959 VSS.n4621 0.00317857
R28852 VSS.n4884 VSS.n4685 0.00317857
R28853 VSS.n4888 VSS.n4887 0.00317857
R28854 VSS.n4928 VSS.n4651 0.00317857
R28855 VSS.n4955 VSS.n4633 0.00317857
R28856 VSS.n4960 VSS.n4958 0.00317857
R28857 VSS.n4974 VSS.n4973 0.00317857
R28858 VSS.n5051 VSS.n4590 0.00317857
R28859 VSS.n5063 VSS.n4585 0.00317857
R28860 VSS.n5093 VSS.n4572 0.00317857
R28861 VSS.n5117 VSS.n5116 0.00317857
R28862 VSS.n5135 VSS.n5134 0.00317857
R28863 VSS.n5095 VSS.n5094 0.00317857
R28864 VSS.n4786 VSS.n4765 0.00317857
R28865 VSS.n4790 VSS.n4789 0.00317857
R28866 VSS.n4818 VSS.n4817 0.00317857
R28867 VSS.n4848 VSS.n4705 0.00317857
R28868 VSS.n4852 VSS.n4851 0.00317857
R28869 VSS.n5377 VSS.n5376 0.00317857
R28870 VSS.n5383 VSS.n5353 0.00317857
R28871 VSS.n5408 VSS.n5326 0.00317857
R28872 VSS.n5319 VSS.n5306 0.00317857
R28873 VSS.n5439 VSS.n5295 0.00317857
R28874 VSS.n5445 VSS.n5288 0.00317857
R28875 VSS.n5475 VSS.n5474 0.00317857
R28876 VSS.n5481 VSS.n5273 0.00317857
R28877 VSS.n5521 VSS.n5242 0.00317857
R28878 VSS.n5530 VSS.n5529 0.00317857
R28879 VSS.n5546 VSS.n5545 0.00317857
R28880 VSS.n5551 VSS.n5213 0.00317857
R28881 VSS.n5476 VSS.n5277 0.00317857
R28882 VSS.n5480 VSS.n5479 0.00317857
R28883 VSS.n5520 VSS.n5243 0.00317857
R28884 VSS.n5547 VSS.n5225 0.00317857
R28885 VSS.n5552 VSS.n5550 0.00317857
R28886 VSS.n5566 VSS.n5565 0.00317857
R28887 VSS.n5643 VSS.n5182 0.00317857
R28888 VSS.n5655 VSS.n5177 0.00317857
R28889 VSS.n5685 VSS.n5164 0.00317857
R28890 VSS.n5709 VSS.n5708 0.00317857
R28891 VSS.n5727 VSS.n5726 0.00317857
R28892 VSS.n5687 VSS.n5686 0.00317857
R28893 VSS.n5378 VSS.n5357 0.00317857
R28894 VSS.n5382 VSS.n5381 0.00317857
R28895 VSS.n5410 VSS.n5409 0.00317857
R28896 VSS.n5440 VSS.n5297 0.00317857
R28897 VSS.n5444 VSS.n5443 0.00317857
R28898 VSS.n5969 VSS.n5968 0.00317857
R28899 VSS.n5975 VSS.n5945 0.00317857
R28900 VSS.n6000 VSS.n5918 0.00317857
R28901 VSS.n5911 VSS.n5898 0.00317857
R28902 VSS.n6031 VSS.n5887 0.00317857
R28903 VSS.n6037 VSS.n5880 0.00317857
R28904 VSS.n6067 VSS.n6066 0.00317857
R28905 VSS.n6073 VSS.n5865 0.00317857
R28906 VSS.n6113 VSS.n5834 0.00317857
R28907 VSS.n6122 VSS.n6121 0.00317857
R28908 VSS.n6138 VSS.n6137 0.00317857
R28909 VSS.n6143 VSS.n5805 0.00317857
R28910 VSS.n6068 VSS.n5869 0.00317857
R28911 VSS.n6072 VSS.n6071 0.00317857
R28912 VSS.n6112 VSS.n5835 0.00317857
R28913 VSS.n6139 VSS.n5817 0.00317857
R28914 VSS.n6144 VSS.n6142 0.00317857
R28915 VSS.n6158 VSS.n6157 0.00317857
R28916 VSS.n6235 VSS.n5774 0.00317857
R28917 VSS.n6247 VSS.n5769 0.00317857
R28918 VSS.n6277 VSS.n5756 0.00317857
R28919 VSS.n6301 VSS.n6300 0.00317857
R28920 VSS.n6319 VSS.n6318 0.00317857
R28921 VSS.n6279 VSS.n6278 0.00317857
R28922 VSS.n5970 VSS.n5949 0.00317857
R28923 VSS.n5974 VSS.n5973 0.00317857
R28924 VSS.n6002 VSS.n6001 0.00317857
R28925 VSS.n6032 VSS.n5889 0.00317857
R28926 VSS.n6036 VSS.n6035 0.00317857
R28927 VSS.n6561 VSS.n6560 0.00317857
R28928 VSS.n6567 VSS.n6537 0.00317857
R28929 VSS.n6592 VSS.n6510 0.00317857
R28930 VSS.n6503 VSS.n6490 0.00317857
R28931 VSS.n6623 VSS.n6479 0.00317857
R28932 VSS.n6629 VSS.n6472 0.00317857
R28933 VSS.n6659 VSS.n6658 0.00317857
R28934 VSS.n6665 VSS.n6457 0.00317857
R28935 VSS.n6705 VSS.n6426 0.00317857
R28936 VSS.n6714 VSS.n6713 0.00317857
R28937 VSS.n6730 VSS.n6729 0.00317857
R28938 VSS.n6735 VSS.n6397 0.00317857
R28939 VSS.n6660 VSS.n6461 0.00317857
R28940 VSS.n6664 VSS.n6663 0.00317857
R28941 VSS.n6704 VSS.n6427 0.00317857
R28942 VSS.n6731 VSS.n6409 0.00317857
R28943 VSS.n6736 VSS.n6734 0.00317857
R28944 VSS.n6750 VSS.n6749 0.00317857
R28945 VSS.n6827 VSS.n6366 0.00317857
R28946 VSS.n6839 VSS.n6361 0.00317857
R28947 VSS.n6869 VSS.n6348 0.00317857
R28948 VSS.n6893 VSS.n6892 0.00317857
R28949 VSS.n6911 VSS.n6910 0.00317857
R28950 VSS.n6871 VSS.n6870 0.00317857
R28951 VSS.n6562 VSS.n6541 0.00317857
R28952 VSS.n6566 VSS.n6565 0.00317857
R28953 VSS.n6594 VSS.n6593 0.00317857
R28954 VSS.n6624 VSS.n6481 0.00317857
R28955 VSS.n6628 VSS.n6627 0.00317857
R28956 VSS.n2405 VSS.n2404 0.00317857
R28957 VSS.n2411 VSS.n2381 0.00317857
R28958 VSS.n2436 VSS.n2354 0.00317857
R28959 VSS.n2347 VSS.n2334 0.00317857
R28960 VSS.n2467 VSS.n2323 0.00317857
R28961 VSS.n2473 VSS.n2316 0.00317857
R28962 VSS.n2559 VSS.n2313 0.00317857
R28963 VSS.n7036 VSS.n2498 0.00317857
R28964 VSS.n7021 VSS.n7020 0.00317857
R28965 VSS.n2595 VSS.n2521 0.00317857
R28966 VSS.n7011 VSS.n2522 0.00317857
R28967 VSS.n7006 VSS.n2527 0.00317857
R28968 VSS.n2558 VSS.n2494 0.00317857
R28969 VSS.n7037 VSS.n2496 0.00317857
R28970 VSS.n7022 VSS.n2511 0.00317857
R28971 VSS.n7010 VSS.n2523 0.00317857
R28972 VSS.n7007 VSS.n2525 0.00317857
R28973 VSS.n2640 VSS.n2639 0.00317857
R28974 VSS.n2697 VSS.n2684 0.00317857
R28975 VSS.n2731 VSS.n2679 0.00317857
R28976 VSS.n6939 VSS.n6938 0.00317857
R28977 VSS.n2765 VSS.n2764 0.00317857
R28978 VSS.n6920 VSS.n2752 0.00317857
R28979 VSS.n6937 VSS.n2712 0.00317857
R28980 VSS.n2406 VSS.n2385 0.00317857
R28981 VSS.n2410 VSS.n2409 0.00317857
R28982 VSS.n2438 VSS.n2437 0.00317857
R28983 VSS.n2468 VSS.n2325 0.00317857
R28984 VSS.n2472 VSS.n2471 0.00317857
R28985 VSS.n3002 VSS.n3001 0.00317857
R28986 VSS.n3008 VSS.n2979 0.00317857
R28987 VSS.n3041 VSS.n2954 0.00317857
R28988 VSS.n3057 VSS.n3056 0.00317857
R28989 VSS.n3074 VSS.n3073 0.00317857
R28990 VSS.n3079 VSS.n2919 0.00317857
R28991 VSS.n3107 VSS.n3106 0.00317857
R28992 VSS.n3113 VSS.n2904 0.00317857
R28993 VSS.n3153 VSS.n2873 0.00317857
R28994 VSS.n3162 VSS.n3161 0.00317857
R28995 VSS.n3178 VSS.n3177 0.00317857
R28996 VSS.n3183 VSS.n2844 0.00317857
R28997 VSS.n3108 VSS.n2908 0.00317857
R28998 VSS.n3112 VSS.n3111 0.00317857
R28999 VSS.n3152 VSS.n2874 0.00317857
R29000 VSS.n3179 VSS.n2856 0.00317857
R29001 VSS.n3184 VSS.n3182 0.00317857
R29002 VSS.n3198 VSS.n3197 0.00317857
R29003 VSS.n3275 VSS.n2813 0.00317857
R29004 VSS.n3287 VSS.n2808 0.00317857
R29005 VSS.n3317 VSS.n2795 0.00317857
R29006 VSS.n3341 VSS.n3340 0.00317857
R29007 VSS.n3359 VSS.n3358 0.00317857
R29008 VSS.n3319 VSS.n3318 0.00317857
R29009 VSS.n3003 VSS.n2983 0.00317857
R29010 VSS.n3007 VSS.n3006 0.00317857
R29011 VSS.n3042 VSS.n2952 0.00317857
R29012 VSS.n3075 VSS.n2931 0.00317857
R29013 VSS.n3080 VSS.n3078 0.00317857
R29014 VSS.n332 VSS.n275 0.00317857
R29015 VSS.n427 VSS.n281 0.00317857
R29016 VSS.n418 VSS.n288 0.00317857
R29017 VSS.n376 VSS.n305 0.00317857
R29018 VSS.n402 VSS.n306 0.00317857
R29019 VSS.n396 VSS.n179 0.00317857
R29020 VSS.n9067 VSS.n9066 0.00317857
R29021 VSS.n9073 VSS.n171 0.00317857
R29022 VSS.n9113 VSS.n140 0.00317857
R29023 VSS.n9122 VSS.n9121 0.00317857
R29024 VSS.n9138 VSS.n9137 0.00317857
R29025 VSS.n9143 VSS.n111 0.00317857
R29026 VSS.n9068 VSS.n175 0.00317857
R29027 VSS.n9072 VSS.n9071 0.00317857
R29028 VSS.n9112 VSS.n141 0.00317857
R29029 VSS.n9139 VSS.n123 0.00317857
R29030 VSS.n9144 VSS.n9142 0.00317857
R29031 VSS.n9158 VSS.n9157 0.00317857
R29032 VSS.n9235 VSS.n80 0.00317857
R29033 VSS.n9247 VSS.n75 0.00317857
R29034 VSS.n9277 VSS.n62 0.00317857
R29035 VSS.n9301 VSS.n9300 0.00317857
R29036 VSS.n9319 VSS.n9318 0.00317857
R29037 VSS.n9279 VSS.n9278 0.00317857
R29038 VSS.n331 VSS.n277 0.00317857
R29039 VSS.n428 VSS.n279 0.00317857
R29040 VSS.n417 VSS.n416 0.00317857
R29041 VSS.n401 VSS.n307 0.00317857
R29042 VSS.n398 VSS.n397 0.00317857
R29043 VSS.n860 VSS.n482 0.00317857
R29044 VSS.n855 VSS.n487 0.00317857
R29045 VSS.n840 VSS.n839 0.00317857
R29046 VSS.n587 VSS.n510 0.00317857
R29047 VSS.n830 VSS.n511 0.00317857
R29048 VSS.n825 VSS.n516 0.00317857
R29049 VSS.n859 VSS.n483 0.00317857
R29050 VSS.n856 VSS.n485 0.00317857
R29051 VSS.n841 VSS.n500 0.00317857
R29052 VSS.n829 VSS.n512 0.00317857
R29053 VSS.n826 VSS.n514 0.00317857
R29054 VSS.n632 VSS.n631 0.00317857
R29055 VSS.n689 VSS.n676 0.00317857
R29056 VSS.n732 VSS.n671 0.00317857
R29057 VSS.n758 VSS.n757 0.00317857
R29058 VSS.n721 VSS.n720 0.00317857
R29059 VSS.n9327 VSS.n34 0.00317857
R29060 VSS.n756 VSS.n704 0.00317857
R29061 VSS.n895 VSS.n443 0.00317857
R29062 VSS.n993 VSS.n445 0.00317857
R29063 VSS.n982 VSS.n981 0.00317857
R29064 VSS.n966 VSS.n473 0.00317857
R29065 VSS.n963 VSS.n475 0.00317857
R29066 VSS.n7208 VSS.n7207 0.00317857
R29067 VSS.n7265 VSS.n7252 0.00317857
R29068 VSS.n7299 VSS.n7247 0.00317857
R29069 VSS.n8367 VSS.n8366 0.00317857
R29070 VSS.n7333 VSS.n7332 0.00317857
R29071 VSS.n8348 VSS.n7320 0.00317857
R29072 VSS.n8365 VSS.n7280 0.00317857
R29073 VSS.n7136 VSS.n7067 0.00228571
R29074 VSS.n7141 VSS.n7136 0.00228571
R29075 VSS.n7137 VSS.n7116 0.00228571
R29076 VSS.n8455 VSS.n7073 0.00228571
R29077 VSS.n7168 VSS.n7167 0.00228571
R29078 VSS.n8454 VSS.n8453 0.00228571
R29079 VSS.n906 VSS.n885 0.00228571
R29080 VSS.n977 VSS.n976 0.00228571
R29081 VSS.n935 VSS.n934 0.00228571
R29082 VSS.n7514 VSS.n7464 0.00228571
R29083 VSS.n7514 VSS.n7513 0.00228571
R29084 VSS.n7525 VSS.n7456 0.00228571
R29085 VSS.n7536 VSS.n7448 0.00228571
R29086 VSS.n7557 VSS.n7556 0.00228571
R29087 VSS.n1087 VSS.n1066 0.00228571
R29088 VSS.n8498 VSS.n8497 0.00228571
R29089 VSS.n1116 VSS.n1115 0.00228571
R29090 VSS.n8499 VSS.n1028 0.00228571
R29091 VSS.n7403 VSS.n7400 0.00228571
R29092 VSS.n7639 VSS.n7638 0.00228571
R29093 VSS.n7390 VSS.n7384 0.00228571
R29094 VSS.n7712 VSS.n7363 0.00228571
R29095 VSS.n7722 VSS.n7721 0.00228571
R29096 VSS.n7537 VSS.n7446 0.00228571
R29097 VSS.n8106 VSS.n7878 0.00228571
R29098 VSS.n8106 VSS.n8105 0.00228571
R29099 VSS.n8117 VSS.n7870 0.00228571
R29100 VSS.n8128 VSS.n7862 0.00228571
R29101 VSS.n8149 VSS.n8148 0.00228571
R29102 VSS.n8012 VSS.n7955 0.00228571
R29103 VSS.n7943 VSS.n7942 0.00228571
R29104 VSS.n8044 VSS.n7926 0.00228571
R29105 VSS.n8030 VSS.n7944 0.00228571
R29106 VSS.n7817 VSS.n7814 0.00228571
R29107 VSS.n8231 VSS.n8230 0.00228571
R29108 VSS.n7804 VSS.n7798 0.00228571
R29109 VSS.n8304 VSS.n7777 0.00228571
R29110 VSS.n8314 VSS.n8313 0.00228571
R29111 VSS.n8129 VSS.n7860 0.00228571
R29112 VSS.n8573 VSS.n252 0.00228571
R29113 VSS.n240 VSS.n239 0.00228571
R29114 VSS.n8605 VSS.n223 0.00228571
R29115 VSS.n8715 VSS.n8646 0.00228571
R29116 VSS.n8720 VSS.n8715 0.00228571
R29117 VSS.n8716 VSS.n8695 0.00228571
R29118 VSS.n9028 VSS.n8652 0.00228571
R29119 VSS.n8747 VSS.n8746 0.00228571
R29120 VSS.n9027 VSS.n9026 0.00228571
R29121 VSS.n8826 VSS.n8779 0.00228571
R29122 VSS.n8976 VSS.n8803 0.00228571
R29123 VSS.n8970 VSS.n8969 0.00228571
R29124 VSS.n8910 VSS.n8906 0.00228571
R29125 VSS.n8885 VSS.n8882 0.00228571
R29126 VSS.n8591 VSS.n241 0.00228571
R29127 VSS.n1255 VSS.n1198 0.00228571
R29128 VSS.n1186 VSS.n1185 0.00228571
R29129 VSS.n1287 VSS.n1169 0.00228571
R29130 VSS.n1397 VSS.n1328 0.00228571
R29131 VSS.n1402 VSS.n1397 0.00228571
R29132 VSS.n1398 VSS.n1377 0.00228571
R29133 VSS.n1691 VSS.n1334 0.00228571
R29134 VSS.n1429 VSS.n1428 0.00228571
R29135 VSS.n1690 VSS.n1689 0.00228571
R29136 VSS.n1648 VSS.n1647 0.00228571
R29137 VSS.n1637 VSS.n1636 0.00228571
R29138 VSS.n1514 VSS.n1500 0.00228571
R29139 VSS.n1542 VSS.n1539 0.00228571
R29140 VSS.n1596 VSS.n1551 0.00228571
R29141 VSS.n1273 VSS.n1187 0.00228571
R29142 VSS.n1828 VSS.n1771 0.00228571
R29143 VSS.n1759 VSS.n1758 0.00228571
R29144 VSS.n1860 VSS.n1742 0.00228571
R29145 VSS.n1970 VSS.n1901 0.00228571
R29146 VSS.n1975 VSS.n1970 0.00228571
R29147 VSS.n1971 VSS.n1950 0.00228571
R29148 VSS.n2283 VSS.n1907 0.00228571
R29149 VSS.n2002 VSS.n2001 0.00228571
R29150 VSS.n2282 VSS.n2281 0.00228571
R29151 VSS.n2240 VSS.n2239 0.00228571
R29152 VSS.n2229 VSS.n2228 0.00228571
R29153 VSS.n2087 VSS.n2073 0.00228571
R29154 VSS.n2115 VSS.n2112 0.00228571
R29155 VSS.n2188 VSS.n2124 0.00228571
R29156 VSS.n1846 VSS.n1760 0.00228571
R29157 VSS.n3622 VSS.n3565 0.00228571
R29158 VSS.n3553 VSS.n3552 0.00228571
R29159 VSS.n3654 VSS.n3536 0.00228571
R29160 VSS.n3716 VSS.n3488 0.00228571
R29161 VSS.n3716 VSS.n3715 0.00228571
R29162 VSS.n3727 VSS.n3480 0.00228571
R29163 VSS.n3738 VSS.n3472 0.00228571
R29164 VSS.n3759 VSS.n3758 0.00228571
R29165 VSS.n3739 VSS.n3470 0.00228571
R29166 VSS.n3427 VSS.n3424 0.00228571
R29167 VSS.n3841 VSS.n3840 0.00228571
R29168 VSS.n3414 VSS.n3408 0.00228571
R29169 VSS.n3914 VSS.n3387 0.00228571
R29170 VSS.n3924 VSS.n3923 0.00228571
R29171 VSS.n3640 VSS.n3554 0.00228571
R29172 VSS.n4214 VSS.n4157 0.00228571
R29173 VSS.n4145 VSS.n4144 0.00228571
R29174 VSS.n4246 VSS.n4128 0.00228571
R29175 VSS.n4308 VSS.n4080 0.00228571
R29176 VSS.n4308 VSS.n4307 0.00228571
R29177 VSS.n4319 VSS.n4072 0.00228571
R29178 VSS.n4330 VSS.n4064 0.00228571
R29179 VSS.n4351 VSS.n4350 0.00228571
R29180 VSS.n4331 VSS.n4062 0.00228571
R29181 VSS.n4019 VSS.n4016 0.00228571
R29182 VSS.n4433 VSS.n4432 0.00228571
R29183 VSS.n4006 VSS.n4000 0.00228571
R29184 VSS.n4506 VSS.n3979 0.00228571
R29185 VSS.n4516 VSS.n4515 0.00228571
R29186 VSS.n4232 VSS.n4146 0.00228571
R29187 VSS.n4806 VSS.n4749 0.00228571
R29188 VSS.n4737 VSS.n4736 0.00228571
R29189 VSS.n4838 VSS.n4720 0.00228571
R29190 VSS.n4900 VSS.n4672 0.00228571
R29191 VSS.n4900 VSS.n4899 0.00228571
R29192 VSS.n4911 VSS.n4664 0.00228571
R29193 VSS.n4922 VSS.n4656 0.00228571
R29194 VSS.n4943 VSS.n4942 0.00228571
R29195 VSS.n4923 VSS.n4654 0.00228571
R29196 VSS.n4611 VSS.n4608 0.00228571
R29197 VSS.n5025 VSS.n5024 0.00228571
R29198 VSS.n4598 VSS.n4592 0.00228571
R29199 VSS.n5098 VSS.n4571 0.00228571
R29200 VSS.n5108 VSS.n5107 0.00228571
R29201 VSS.n4824 VSS.n4738 0.00228571
R29202 VSS.n5398 VSS.n5341 0.00228571
R29203 VSS.n5329 VSS.n5328 0.00228571
R29204 VSS.n5430 VSS.n5312 0.00228571
R29205 VSS.n5492 VSS.n5264 0.00228571
R29206 VSS.n5492 VSS.n5491 0.00228571
R29207 VSS.n5503 VSS.n5256 0.00228571
R29208 VSS.n5514 VSS.n5248 0.00228571
R29209 VSS.n5535 VSS.n5534 0.00228571
R29210 VSS.n5515 VSS.n5246 0.00228571
R29211 VSS.n5203 VSS.n5200 0.00228571
R29212 VSS.n5617 VSS.n5616 0.00228571
R29213 VSS.n5190 VSS.n5184 0.00228571
R29214 VSS.n5690 VSS.n5163 0.00228571
R29215 VSS.n5700 VSS.n5699 0.00228571
R29216 VSS.n5416 VSS.n5330 0.00228571
R29217 VSS.n5990 VSS.n5933 0.00228571
R29218 VSS.n5921 VSS.n5920 0.00228571
R29219 VSS.n6022 VSS.n5904 0.00228571
R29220 VSS.n6084 VSS.n5856 0.00228571
R29221 VSS.n6084 VSS.n6083 0.00228571
R29222 VSS.n6095 VSS.n5848 0.00228571
R29223 VSS.n6106 VSS.n5840 0.00228571
R29224 VSS.n6127 VSS.n6126 0.00228571
R29225 VSS.n6107 VSS.n5838 0.00228571
R29226 VSS.n5795 VSS.n5792 0.00228571
R29227 VSS.n6209 VSS.n6208 0.00228571
R29228 VSS.n5782 VSS.n5776 0.00228571
R29229 VSS.n6282 VSS.n5755 0.00228571
R29230 VSS.n6292 VSS.n6291 0.00228571
R29231 VSS.n6008 VSS.n5922 0.00228571
R29232 VSS.n6582 VSS.n6525 0.00228571
R29233 VSS.n6513 VSS.n6512 0.00228571
R29234 VSS.n6614 VSS.n6496 0.00228571
R29235 VSS.n6676 VSS.n6448 0.00228571
R29236 VSS.n6676 VSS.n6675 0.00228571
R29237 VSS.n6687 VSS.n6440 0.00228571
R29238 VSS.n6698 VSS.n6432 0.00228571
R29239 VSS.n6719 VSS.n6718 0.00228571
R29240 VSS.n6699 VSS.n6430 0.00228571
R29241 VSS.n6387 VSS.n6384 0.00228571
R29242 VSS.n6801 VSS.n6800 0.00228571
R29243 VSS.n6374 VSS.n6368 0.00228571
R29244 VSS.n6874 VSS.n6347 0.00228571
R29245 VSS.n6884 VSS.n6883 0.00228571
R29246 VSS.n6600 VSS.n6514 0.00228571
R29247 VSS.n2426 VSS.n2369 0.00228571
R29248 VSS.n2357 VSS.n2356 0.00228571
R29249 VSS.n2458 VSS.n2340 0.00228571
R29250 VSS.n2568 VSS.n2499 0.00228571
R29251 VSS.n2573 VSS.n2568 0.00228571
R29252 VSS.n2569 VSS.n2548 0.00228571
R29253 VSS.n7027 VSS.n2505 0.00228571
R29254 VSS.n2600 VSS.n2599 0.00228571
R29255 VSS.n7026 VSS.n7025 0.00228571
R29256 VSS.n6984 VSS.n6983 0.00228571
R29257 VSS.n6973 VSS.n6972 0.00228571
R29258 VSS.n2685 VSS.n2671 0.00228571
R29259 VSS.n2713 VSS.n2710 0.00228571
R29260 VSS.n6932 VSS.n2722 0.00228571
R29261 VSS.n2444 VSS.n2358 0.00228571
R29262 VSS.n3030 VSS.n2964 0.00228571
R29263 VSS.n3048 VSS.n2948 0.00228571
R29264 VSS.n3062 VSS.n3061 0.00228571
R29265 VSS.n3124 VSS.n2895 0.00228571
R29266 VSS.n3124 VSS.n3123 0.00228571
R29267 VSS.n3135 VSS.n2887 0.00228571
R29268 VSS.n3146 VSS.n2879 0.00228571
R29269 VSS.n3167 VSS.n3166 0.00228571
R29270 VSS.n3147 VSS.n2877 0.00228571
R29271 VSS.n2834 VSS.n2831 0.00228571
R29272 VSS.n3249 VSS.n3248 0.00228571
R29273 VSS.n2821 VSS.n2815 0.00228571
R29274 VSS.n3322 VSS.n2794 0.00228571
R29275 VSS.n3332 VSS.n3331 0.00228571
R29276 VSS.n3047 VSS.n2949 0.00228571
R29277 VSS.n354 VSS.n353 0.00228571
R29278 VSS.n412 VSS.n411 0.00228571
R29279 VSS.n372 VSS.n371 0.00228571
R29280 VSS.n9084 VSS.n162 0.00228571
R29281 VSS.n9084 VSS.n9083 0.00228571
R29282 VSS.n9095 VSS.n154 0.00228571
R29283 VSS.n9106 VSS.n146 0.00228571
R29284 VSS.n9127 VSS.n9126 0.00228571
R29285 VSS.n9107 VSS.n144 0.00228571
R29286 VSS.n101 VSS.n98 0.00228571
R29287 VSS.n9209 VSS.n9208 0.00228571
R29288 VSS.n88 VSS.n82 0.00228571
R29289 VSS.n9282 VSS.n61 0.00228571
R29290 VSS.n9292 VSS.n9291 0.00228571
R29291 VSS.n413 VSS.n295 0.00228571
R29292 VSS.n560 VSS.n488 0.00228571
R29293 VSS.n565 VSS.n560 0.00228571
R29294 VSS.n561 VSS.n537 0.00228571
R29295 VSS.n846 VSS.n494 0.00228571
R29296 VSS.n592 VSS.n591 0.00228571
R29297 VSS.n845 VSS.n844 0.00228571
R29298 VSS.n803 VSS.n802 0.00228571
R29299 VSS.n792 VSS.n791 0.00228571
R29300 VSS.n677 VSS.n663 0.00228571
R29301 VSS.n705 VSS.n702 0.00228571
R29302 VSS.n751 VSS.n714 0.00228571
R29303 VSS.n978 VSS.n461 0.00228571
R29304 VSS.n8412 VSS.n8411 0.00228571
R29305 VSS.n8401 VSS.n8400 0.00228571
R29306 VSS.n7253 VSS.n7239 0.00228571
R29307 VSS.n7281 VSS.n7278 0.00228571
R29308 VSS.n8360 VSS.n7290 0.00228571
R29309 VSS.n8517 VSS.n8516 0.00217857
R29310 VSS.n8515 VSS.n1011 0.00217857
R29311 VSS.n8486 VSS.n1035 0.00217857
R29312 VSS.n8485 VSS.n1041 0.00217857
R29313 VSS.n7499 VSS.n7475 0.00217857
R29314 VSS.n7500 VSS.n7461 0.00217857
R29315 VSS.n7570 VSS.n7423 0.00217857
R29316 VSS.n7571 VSS.n7411 0.00217857
R29317 VSS.n7993 VSS.n7969 0.00217857
R29318 VSS.n7994 VSS.n7949 0.00217857
R29319 VSS.n8055 VSS.n7918 0.00217857
R29320 VSS.n8056 VSS.n7900 0.00217857
R29321 VSS.n8091 VSS.n7889 0.00217857
R29322 VSS.n8092 VSS.n7875 0.00217857
R29323 VSS.n8162 VSS.n7837 0.00217857
R29324 VSS.n8163 VSS.n7825 0.00217857
R29325 VSS.n8554 VSS.n266 0.00217857
R29326 VSS.n8555 VSS.n246 0.00217857
R29327 VSS.n8616 VSS.n215 0.00217857
R29328 VSS.n8617 VSS.n197 0.00217857
R29329 VSS.n9041 VSS.n9040 0.00217857
R29330 VSS.n9039 VSS.n8642 0.00217857
R29331 VSS.n9010 VSS.n8665 0.00217857
R29332 VSS.n9009 VSS.n8671 0.00217857
R29333 VSS.n1236 VSS.n1212 0.00217857
R29334 VSS.n1237 VSS.n1192 0.00217857
R29335 VSS.n1298 VSS.n1161 0.00217857
R29336 VSS.n1299 VSS.n1143 0.00217857
R29337 VSS.n1704 VSS.n1703 0.00217857
R29338 VSS.n1702 VSS.n1324 0.00217857
R29339 VSS.n1673 VSS.n1347 0.00217857
R29340 VSS.n1672 VSS.n1353 0.00217857
R29341 VSS.n1809 VSS.n1785 0.00217857
R29342 VSS.n1810 VSS.n1765 0.00217857
R29343 VSS.n1871 VSS.n1734 0.00217857
R29344 VSS.n1872 VSS.n1716 0.00217857
R29345 VSS.n2296 VSS.n2295 0.00217857
R29346 VSS.n2294 VSS.n1897 0.00217857
R29347 VSS.n2265 VSS.n1920 0.00217857
R29348 VSS.n2264 VSS.n1926 0.00217857
R29349 VSS.n3603 VSS.n3579 0.00217857
R29350 VSS.n3604 VSS.n3559 0.00217857
R29351 VSS.n3665 VSS.n3528 0.00217857
R29352 VSS.n3666 VSS.n3510 0.00217857
R29353 VSS.n3701 VSS.n3499 0.00217857
R29354 VSS.n3702 VSS.n3485 0.00217857
R29355 VSS.n3772 VSS.n3447 0.00217857
R29356 VSS.n3773 VSS.n3435 0.00217857
R29357 VSS.n4195 VSS.n4171 0.00217857
R29358 VSS.n4196 VSS.n4151 0.00217857
R29359 VSS.n4257 VSS.n4120 0.00217857
R29360 VSS.n4258 VSS.n4102 0.00217857
R29361 VSS.n4293 VSS.n4091 0.00217857
R29362 VSS.n4294 VSS.n4077 0.00217857
R29363 VSS.n4364 VSS.n4039 0.00217857
R29364 VSS.n4365 VSS.n4027 0.00217857
R29365 VSS.n4787 VSS.n4763 0.00217857
R29366 VSS.n4788 VSS.n4743 0.00217857
R29367 VSS.n4849 VSS.n4712 0.00217857
R29368 VSS.n4850 VSS.n4694 0.00217857
R29369 VSS.n4885 VSS.n4683 0.00217857
R29370 VSS.n4886 VSS.n4669 0.00217857
R29371 VSS.n4956 VSS.n4631 0.00217857
R29372 VSS.n4957 VSS.n4619 0.00217857
R29373 VSS.n5379 VSS.n5355 0.00217857
R29374 VSS.n5380 VSS.n5335 0.00217857
R29375 VSS.n5441 VSS.n5304 0.00217857
R29376 VSS.n5442 VSS.n5286 0.00217857
R29377 VSS.n5477 VSS.n5275 0.00217857
R29378 VSS.n5478 VSS.n5261 0.00217857
R29379 VSS.n5548 VSS.n5223 0.00217857
R29380 VSS.n5549 VSS.n5211 0.00217857
R29381 VSS.n5971 VSS.n5947 0.00217857
R29382 VSS.n5972 VSS.n5927 0.00217857
R29383 VSS.n6033 VSS.n5896 0.00217857
R29384 VSS.n6034 VSS.n5878 0.00217857
R29385 VSS.n6069 VSS.n5867 0.00217857
R29386 VSS.n6070 VSS.n5853 0.00217857
R29387 VSS.n6140 VSS.n5815 0.00217857
R29388 VSS.n6141 VSS.n5803 0.00217857
R29389 VSS.n6563 VSS.n6539 0.00217857
R29390 VSS.n6564 VSS.n6519 0.00217857
R29391 VSS.n6625 VSS.n6488 0.00217857
R29392 VSS.n6626 VSS.n6470 0.00217857
R29393 VSS.n6661 VSS.n6459 0.00217857
R29394 VSS.n6662 VSS.n6445 0.00217857
R29395 VSS.n6732 VSS.n6407 0.00217857
R29396 VSS.n6733 VSS.n6395 0.00217857
R29397 VSS.n2407 VSS.n2383 0.00217857
R29398 VSS.n2408 VSS.n2363 0.00217857
R29399 VSS.n2469 VSS.n2332 0.00217857
R29400 VSS.n2470 VSS.n2314 0.00217857
R29401 VSS.n7040 VSS.n7039 0.00217857
R29402 VSS.n7038 VSS.n2495 0.00217857
R29403 VSS.n7009 VSS.n2518 0.00217857
R29404 VSS.n7008 VSS.n2524 0.00217857
R29405 VSS.n3004 VSS.n2981 0.00217857
R29406 VSS.n3005 VSS.n2969 0.00217857
R29407 VSS.n3076 VSS.n2929 0.00217857
R29408 VSS.n3077 VSS.n2917 0.00217857
R29409 VSS.n3109 VSS.n2906 0.00217857
R29410 VSS.n3110 VSS.n2892 0.00217857
R29411 VSS.n3180 VSS.n2854 0.00217857
R29412 VSS.n3181 VSS.n2842 0.00217857
R29413 VSS.n431 VSS.n430 0.00217857
R29414 VSS.n429 VSS.n278 0.00217857
R29415 VSS.n400 VSS.n302 0.00217857
R29416 VSS.n399 VSS.n177 0.00217857
R29417 VSS.n9069 VSS.n173 0.00217857
R29418 VSS.n9070 VSS.n159 0.00217857
R29419 VSS.n9140 VSS.n121 0.00217857
R29420 VSS.n9141 VSS.n109 0.00217857
R29421 VSS.n996 VSS.n995 0.00217857
R29422 VSS.n994 VSS.n444 0.00217857
R29423 VSS.n965 VSS.n468 0.00217857
R29424 VSS.n964 VSS.n474 0.00217857
R29425 VSS.n858 VSS.n479 0.00217857
R29426 VSS.n857 VSS.n484 0.00217857
R29427 VSS.n828 VSS.n507 0.00217857
R29428 VSS.n827 VSS.n513 0.00217857
R29429 VSS.n8468 VSS.n8467 0.00217857
R29430 VSS.n8466 VSS.n7063 0.00217857
R29431 VSS.n8437 VSS.n7086 0.00217857
R29432 VSS.n8436 VSS.n7092 0.00217857
R29433 VSS.n7177 VSS.n7106 0.00139286
R29434 VSS.n7183 VSS.n7103 0.00139286
R29435 VSS.n879 VSS.n462 0.00139286
R29436 VSS.n945 VSS.n874 0.00139286
R29437 VSS.n951 VSS.n871 0.00139286
R29438 VSS.n7566 VSS.n7429 0.00139286
R29439 VSS.n7578 VSS.n7420 0.00139286
R29440 VSS.n1060 VSS.n1029 0.00139286
R29441 VSS.n1126 VSS.n1055 0.00139286
R29442 VSS.n1132 VSS.n1052 0.00139286
R29443 VSS.n1027 VSS.n1024 0.00139286
R29444 VSS.n7680 VSS.n7675 0.00139286
R29445 VSS.n7684 VSS.n7683 0.00139286
R29446 VSS.n7676 VSS.n7379 0.00139286
R29447 VSS.n7685 VSS.n7674 0.00139286
R29448 VSS.n8158 VSS.n7843 0.00139286
R29449 VSS.n8170 VSS.n7834 0.00139286
R29450 VSS.n8033 VSS.n8032 0.00139286
R29451 VSS.n8066 VSS.n8065 0.00139286
R29452 VSS.n7917 VSS.n7913 0.00139286
R29453 VSS.n8031 VSS.n7941 0.00139286
R29454 VSS.n8272 VSS.n8267 0.00139286
R29455 VSS.n8276 VSS.n8275 0.00139286
R29456 VSS.n8268 VSS.n7793 0.00139286
R29457 VSS.n8277 VSS.n8266 0.00139286
R29458 VSS.n8594 VSS.n8593 0.00139286
R29459 VSS.n8627 VSS.n8626 0.00139286
R29460 VSS.n214 VSS.n210 0.00139286
R29461 VSS.n8756 VSS.n8685 0.00139286
R29462 VSS.n8762 VSS.n8682 0.00139286
R29463 VSS.n8869 VSS.n8857 0.00139286
R29464 VSS.n8872 VSS.n8851 0.00139286
R29465 VSS.n8860 VSS.n8858 0.00139286
R29466 VSS.n8874 VSS.n8873 0.00139286
R29467 VSS.n8592 VSS.n238 0.00139286
R29468 VSS.n1276 VSS.n1275 0.00139286
R29469 VSS.n1309 VSS.n1308 0.00139286
R29470 VSS.n1160 VSS.n1156 0.00139286
R29471 VSS.n1438 VSS.n1367 0.00139286
R29472 VSS.n1444 VSS.n1364 0.00139286
R29473 VSS.n1576 VSS.n1574 0.00139286
R29474 VSS.n1614 VSS.n1613 0.00139286
R29475 VSS.n1575 VSS.n1510 0.00139286
R29476 VSS.n1615 VSS.n1534 0.00139286
R29477 VSS.n1274 VSS.n1184 0.00139286
R29478 VSS.n1849 VSS.n1848 0.00139286
R29479 VSS.n1882 VSS.n1881 0.00139286
R29480 VSS.n1733 VSS.n1729 0.00139286
R29481 VSS.n2011 VSS.n1940 0.00139286
R29482 VSS.n2017 VSS.n1937 0.00139286
R29483 VSS.n2136 VSS.n2134 0.00139286
R29484 VSS.n2206 VSS.n2205 0.00139286
R29485 VSS.n2135 VSS.n2083 0.00139286
R29486 VSS.n2207 VSS.n2107 0.00139286
R29487 VSS.n1847 VSS.n1757 0.00139286
R29488 VSS.n3643 VSS.n3642 0.00139286
R29489 VSS.n3676 VSS.n3675 0.00139286
R29490 VSS.n3527 VSS.n3523 0.00139286
R29491 VSS.n3768 VSS.n3453 0.00139286
R29492 VSS.n3780 VSS.n3444 0.00139286
R29493 VSS.n3882 VSS.n3877 0.00139286
R29494 VSS.n3886 VSS.n3885 0.00139286
R29495 VSS.n3878 VSS.n3403 0.00139286
R29496 VSS.n3887 VSS.n3876 0.00139286
R29497 VSS.n3641 VSS.n3551 0.00139286
R29498 VSS.n4235 VSS.n4234 0.00139286
R29499 VSS.n4268 VSS.n4267 0.00139286
R29500 VSS.n4119 VSS.n4115 0.00139286
R29501 VSS.n4360 VSS.n4045 0.00139286
R29502 VSS.n4372 VSS.n4036 0.00139286
R29503 VSS.n4474 VSS.n4469 0.00139286
R29504 VSS.n4478 VSS.n4477 0.00139286
R29505 VSS.n4470 VSS.n3995 0.00139286
R29506 VSS.n4479 VSS.n4468 0.00139286
R29507 VSS.n4233 VSS.n4143 0.00139286
R29508 VSS.n4827 VSS.n4826 0.00139286
R29509 VSS.n4860 VSS.n4859 0.00139286
R29510 VSS.n4711 VSS.n4707 0.00139286
R29511 VSS.n4952 VSS.n4637 0.00139286
R29512 VSS.n4964 VSS.n4628 0.00139286
R29513 VSS.n5066 VSS.n5061 0.00139286
R29514 VSS.n5070 VSS.n5069 0.00139286
R29515 VSS.n5062 VSS.n4587 0.00139286
R29516 VSS.n5071 VSS.n5060 0.00139286
R29517 VSS.n4825 VSS.n4735 0.00139286
R29518 VSS.n5419 VSS.n5418 0.00139286
R29519 VSS.n5452 VSS.n5451 0.00139286
R29520 VSS.n5303 VSS.n5299 0.00139286
R29521 VSS.n5544 VSS.n5229 0.00139286
R29522 VSS.n5556 VSS.n5220 0.00139286
R29523 VSS.n5658 VSS.n5653 0.00139286
R29524 VSS.n5662 VSS.n5661 0.00139286
R29525 VSS.n5654 VSS.n5179 0.00139286
R29526 VSS.n5663 VSS.n5652 0.00139286
R29527 VSS.n5417 VSS.n5327 0.00139286
R29528 VSS.n6011 VSS.n6010 0.00139286
R29529 VSS.n6044 VSS.n6043 0.00139286
R29530 VSS.n5895 VSS.n5891 0.00139286
R29531 VSS.n6136 VSS.n5821 0.00139286
R29532 VSS.n6148 VSS.n5812 0.00139286
R29533 VSS.n6250 VSS.n6245 0.00139286
R29534 VSS.n6254 VSS.n6253 0.00139286
R29535 VSS.n6246 VSS.n5771 0.00139286
R29536 VSS.n6255 VSS.n6244 0.00139286
R29537 VSS.n6009 VSS.n5919 0.00139286
R29538 VSS.n6603 VSS.n6602 0.00139286
R29539 VSS.n6636 VSS.n6635 0.00139286
R29540 VSS.n6487 VSS.n6483 0.00139286
R29541 VSS.n6728 VSS.n6413 0.00139286
R29542 VSS.n6740 VSS.n6404 0.00139286
R29543 VSS.n6842 VSS.n6837 0.00139286
R29544 VSS.n6846 VSS.n6845 0.00139286
R29545 VSS.n6838 VSS.n6363 0.00139286
R29546 VSS.n6847 VSS.n6836 0.00139286
R29547 VSS.n6601 VSS.n6511 0.00139286
R29548 VSS.n2447 VSS.n2446 0.00139286
R29549 VSS.n2480 VSS.n2479 0.00139286
R29550 VSS.n2331 VSS.n2327 0.00139286
R29551 VSS.n2609 VSS.n2538 0.00139286
R29552 VSS.n2615 VSS.n2535 0.00139286
R29553 VSS.n2734 VSS.n2732 0.00139286
R29554 VSS.n6950 VSS.n6949 0.00139286
R29555 VSS.n2733 VSS.n2681 0.00139286
R29556 VSS.n6951 VSS.n2705 0.00139286
R29557 VSS.n2445 VSS.n2355 0.00139286
R29558 VSS.n3040 VSS.n2956 0.00139286
R29559 VSS.n3072 VSS.n2935 0.00139286
R29560 VSS.n3084 VSS.n2926 0.00139286
R29561 VSS.n3176 VSS.n2860 0.00139286
R29562 VSS.n3188 VSS.n2851 0.00139286
R29563 VSS.n3290 VSS.n3285 0.00139286
R29564 VSS.n3294 VSS.n3293 0.00139286
R29565 VSS.n3286 VSS.n2810 0.00139286
R29566 VSS.n3295 VSS.n3284 0.00139286
R29567 VSS.n2955 VSS.n2953 0.00139286
R29568 VSS.n362 VSS.n296 0.00139286
R29569 VSS.n379 VSS.n311 0.00139286
R29570 VSS.n390 VSS.n309 0.00139286
R29571 VSS.n9136 VSS.n127 0.00139286
R29572 VSS.n9148 VSS.n118 0.00139286
R29573 VSS.n9250 VSS.n9245 0.00139286
R29574 VSS.n9254 VSS.n9253 0.00139286
R29575 VSS.n9246 VSS.n77 0.00139286
R29576 VSS.n9255 VSS.n9244 0.00139286
R29577 VSS.n294 VSS.n291 0.00139286
R29578 VSS.n601 VSS.n527 0.00139286
R29579 VSS.n607 VSS.n524 0.00139286
R29580 VSS.n735 VSS.n733 0.00139286
R29581 VSS.n769 VSS.n768 0.00139286
R29582 VSS.n734 VSS.n673 0.00139286
R29583 VSS.n770 VSS.n697 0.00139286
R29584 VSS.n460 VSS.n457 0.00139286
R29585 VSS.n7302 VSS.n7300 0.00139286
R29586 VSS.n8378 VSS.n8377 0.00139286
R29587 VSS.n7301 VSS.n7249 0.00139286
R29588 VSS.n8379 VSS.n7273 0.00139286
R29589 VSS.n8344 VSS.n8343 0.00054824
R29590 VSS.n7752 VSS.n7751 0.00054824
R29591 VSS.n9352 VSS.n9351 0.00054824
R29592 VSS.n2173 VSS.n0 0.00054824
R29593 VSS.n3955 VSS.n3954 0.00054824
R29594 VSS.n4547 VSS.n4546 0.00054824
R29595 VSS.n5139 VSS.n5138 0.00054824
R29596 VSS.n5731 VSS.n5730 0.00054824
R29597 VSS.n6323 VSS.n6322 0.00054824
R29598 VSS.n6915 VSS.n6914 0.00054824
R29599 VSS.n6917 VSS.n6916 0.00054824
R29600 VSS.n3363 VSS.n3362 0.00054824
R29601 VSS.n8892 VSS.n37 0.00054824
R29602 VSS.n9323 VSS.n9322 0.00054824
R29603 D2_BUF.n2 D2_BUF.n1 173.293
R29604 D2_BUF.n1 D2_BUF.t3 84.3505
R29605 D2_BUF.n1 D2_BUF.t2 53.5025
R29606 D2_BUF.n0 D2_BUF.t0 46.9077
R29607 D2_BUF.n0 D2_BUF.t1 35.0239
R29608 D2_BUF D2_BUF.n2 3.75226
R29609 D2_BUF.n2 D2_BUF.n0 0.204238
R29610 switch_n_3v3_0.D4.n0 switch_n_3v3_0.D4.n1 173.293
R29611 switch_n_3v3_0.D4 switch_n_3v3_0.D4.n2 125.046
R29612 switch_n_3v3_0.D4.n1 switch_n_3v3_0.D4.t5 84.3505
R29613 switch_n_3v3_0.D4.n2 switch_n_3v3_0.D4.t4 77.1205
R29614 switch_n_3v3_0.D4.n2 switch_n_3v3_0.D4.t3 61.6965
R29615 switch_n_3v3_0.D4.n1 switch_n_3v3_0.D4.t2 53.5025
R29616 switch_n_3v3_0.D4.n0 switch_n_3v3_0.D4.t0 46.9077
R29617 switch_n_3v3_0.D4.n0 switch_n_3v3_0.D4.t1 35.0239
R29618 switch_n_3v3_0.D4 switch_n_3v3_0.D4.n0 3.95498
R29619 D5_BUF.n2 D5_BUF.n1 173.293
R29620 D5_BUF.n1 D5_BUF.t2 84.3505
R29621 D5_BUF.n1 D5_BUF.t3 53.5025
R29622 D5_BUF.n0 D5_BUF.t0 46.9077
R29623 D5_BUF.n0 D5_BUF.t1 35.0239
R29624 D5_BUF D5_BUF.n2 3.74964
R29625 D5_BUF.n2 D5_BUF.n0 0.204238
R29626 VOUT.n0 VOUT.t2 46.8495
R29627 VOUT.n0 VOUT.t1 46.5654
R29628 VOUT.n5 VOUT.t3 34.887
R29629 VOUT.n10 VOUT.t0 27.6955
R29630 VOUT.n4 VOUT.n3 13.362
R29631 VOUT.n2 VOUT.n1 9.3005
R29632 VOUT.n7 VOUT.n6 9.3005
R29633 VOUT.n9 VOUT.n8 9.3005
R29634 VOUT.n12 VOUT.n11 9.3005
R29635 VOUT.n11 VOUT.n10 9.02061
R29636 VOUT.n5 VOUT.n4 4.55875
R29637 VOUT.n0 VOUT 3.09322
R29638 VOUT VOUT.n12 0.815717
R29639 VOUT.n2 VOUT.n0 0.613
R29640 VOUT.n12 VOUT.n9 0.0439783
R29641 VOUT.n7 VOUT.n5 0.0439783
R29642 VOUT.n5 VOUT.n2 0.014087
R29643 VOUT.n9 VOUT.n7 0.00321739
R29644 switch_n_3v3_0.D3.n0 switch_n_3v3_0.D3.n1 173.293
R29645 switch_n_3v3_0.D3 switch_n_3v3_0.D3.n2 125.046
R29646 switch_n_3v3_0.D3.n1 switch_n_3v3_0.D3.t3 84.3505
R29647 switch_n_3v3_0.D3.n2 switch_n_3v3_0.D3.t2 77.1205
R29648 switch_n_3v3_0.D3.n2 switch_n_3v3_0.D3.t5 61.6965
R29649 switch_n_3v3_0.D3.n1 switch_n_3v3_0.D3.t4 53.5025
R29650 switch_n_3v3_0.D3.n0 switch_n_3v3_0.D3.t0 46.9077
R29651 switch_n_3v3_0.D3.n0 switch_n_3v3_0.D3.t1 35.0239
R29652 switch_n_3v3_0.D3 switch_n_3v3_0.D3.n0 3.95473
R29653 D4_BUF.n2 D4_BUF.n1 173.293
R29654 D4_BUF.n1 D4_BUF.t3 84.3505
R29655 D4_BUF.n1 D4_BUF.t2 53.5025
R29656 D4_BUF.n0 D4_BUF.t0 46.9077
R29657 D4_BUF.n0 D4_BUF.t1 35.0239
R29658 D4_BUF D4_BUF.n2 3.75124
R29659 D4_BUF.n2 D4_BUF.n0 0.204238
R29660 D3_BUF.n2 D3_BUF.n1 173.293
R29661 D3_BUF.n1 D3_BUF.t2 84.3505
R29662 D3_BUF.n1 D3_BUF.t3 53.5025
R29663 D3_BUF.n0 D3_BUF.t0 46.9077
R29664 D3_BUF.n0 D3_BUF.t1 35.0239
R29665 D3_BUF D3_BUF.n2 3.75099
R29666 D3_BUF.n2 D3_BUF.n0 0.204238
R29667 D3 D3.n0 125.046
R29668 D3.n0 D3.t1 77.1205
R29669 D3.n0 D3.t0 61.6965
R29670 VREFL.n1 VREFL.t0 99.7169
R29671 VREFL.n0 VREFL.t1 44.9543
R29672 VREFL.n0 VREFL.t2 37.5373
R29673 VREFL.n1 VREFL.n0 2.88557
R29674 VREFL VREFL.n1 1.84958
R29675 D4 D4.n0 125.046
R29676 D4.n0 D4.t1 77.1205
R29677 D4.n0 D4.t0 61.6965
R29678 D0 D0.n0 115.853
R29679 D0.n0 D0.t1 81.9405
R29680 D0.n0 D0.t0 56.8765
R29681 D1.n1 D1.n0 127.099
R29682 D1.n0 D1.t1 77.6025
R29683 D1.n0 D1.t0 61.2145
R29684 D1.n1 D1 0.0485769
R29685 D1 D1.n1 0.0365577
R29686 D1_BUF.n2 D1_BUF.n1 169.566
R29687 D1_BUF.n1 D1_BUF.t2 84.8325
R29688 D1_BUF.n1 D1_BUF.t3 53.0205
R29689 D1_BUF.n0 D1_BUF.t0 46.9158
R29690 D1_BUF.n0 D1_BUF.t1 35.0302
R29691 D1_BUF.n3 D1_BUF.n2 3.65455
R29692 D1_BUF D1_BUF.n3 2.58512
R29693 D1_BUF.n2 D1_BUF.n0 0.199588
R29694 D1_BUF.n3 D1_BUF 0.0389615
R29695 D2 D2.n0 125.046
R29696 D2.n0 D2.t0 77.1205
R29697 D2.n0 D2.t1 61.6965
R29698 VREFH VREFH.t0 98.0324
R29699 D5 D5.n0 125.046
R29700 D5.n0 D5.t1 77.1205
R29701 D5.n0 D5.t0 61.6965
C3488 switch_n_3v3_0.D7 VSS 3.4f
C3489 switch_n_3v3_0.D6 VSS 1.41f
C3490 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS 0.667f 
C3491 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS 1.53f 
C3492 D1_BUF VSS 1.17f
C3493 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS 1.13f 
C3494 D0_BUF VSS 2.53f
C3495 a_1556_406# VSS 1.22f 
C3496 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS 0.676f 
C3497 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS 0.519f 
C3498 VREFH VSS 0.29f
C3499 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH VSS 0.544f 
C3500 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS 1.32f 
C3501 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VSS 1.08f 
C3502 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS 0.627f 
C3503 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS 1.07f 
C3504 D2_BUF VSS 1.14f
C3505 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ VSS 1.14f 
C3506 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 VSS 1.63f 
C3507 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS 1.06f 
C3508 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 VSS 3.26f 
C3509 a_1556_1634# VSS 1.16f 
C3510 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS 0.663f 
C3511 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS 0.467f 
C3512 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS 1.5f 
C3513 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH VSS 0.543f 
C3514 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].VOUT VSS 0.95f 
C3515 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS 0.633f 
C3516 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS 1.07f 
C3517 D3_BUF VSS 1.17f
C3518 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.DX_ VSS 1.09f 
C3519 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D1 VSS 1.61f 
C3520 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS 1.06f 
C3521 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[0].D0 VSS 3.25f 
C3522 a_1556_2862# VSS 1.16f 
C3523 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS 0.663f 
C3524 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS 0.467f 
C3525 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VREFH VSS 1.42f 
C3526 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH VSS 0.543f 
C3527 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VSS 0.982f 
C3528 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].VOUT VSS 0.875f 
C3529 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VSS 0.984f 
C3530 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS 0.627f 
C3531 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS 1.07f 
C3532 5_bit_dac_0[0].4_bit_dac_0[0].switch_n_3v3_0.D2 VSS 1.87f 
C3533 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ VSS 1.08f 
C3534 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 VSS 1.61f 
C3535 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS 1.06f 
C3536 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 VSS 3.25f 
C3537 a_1556_4090# VSS 1.16f 
C3538 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS 0.663f 
C3539 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS 0.467f 
C3540 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS 1.42f 
C3541 5_bit_dac_0[0].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH VSS 0.543f 
C3542 5_bit_dac_0[0].4_bit_dac_0[0].VOUT VSS 1.46f 
C3543 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS 0.633f 
C3544 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS 1.08f 
C3545 D4_BUF VSS 2.68f
C3546 5_bit_dac_0[0].switch_n_3v3_0.DX_ VSS 1.08f 
C3547 5_bit_dac_0[0].4_bit_dac_0[0].D1 VSS 1.61f 
C3548 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS 1.06f 
C3549 5_bit_dac_0[0].4_bit_dac_0[0].D0 VSS 3.25f 
C3550 a_1556_5318# VSS 1.16f 
C3551 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS 0.663f 
C3552 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS 0.467f 
C3553 5_bit_dac_0[0].4_bit_dac_0[1].VREFH VSS 1.42f 
C3554 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH VSS 0.543f 
C3555 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS 1.02f 
C3556 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VSS 1.02f 
C3557 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS 0.627f 
C3558 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS 1.07f 
C3559 5_bit_dac_0[0].switch_n_3v3_0.D2 VSS 1.86f 
C3560 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ VSS 1.08f 
C3561 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 VSS 1.61f 
C3562 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS 1.06f 
C3563 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 VSS 3.25f 
C3564 a_1556_6546# VSS 1.16f 
C3565 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS 0.663f 
C3566 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS 0.467f 
C3567 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS 1.42f 
C3568 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH VSS 0.543f 
C3569 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].VOUT VSS 0.863f 
C3570 5_bit_dac_0[0].4_bit_dac_0[1].VOUT VSS 1.24f 
C3571 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS 0.633f 
C3572 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS 1.07f 
C3573 5_bit_dac_0[0].switch_n_3v3_0.D3 VSS 1.89f 
C3574 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.DX_ VSS 1.08f 
C3575 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D1 VSS 1.61f 
C3576 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS 1.06f 
C3577 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[0].D0 VSS 3.25f 
C3578 a_1556_7774# VSS 1.16f 
C3579 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS 0.663f 
C3580 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS 0.467f 
C3581 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VREFH VSS 1.42f 
C3582 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH VSS 0.543f 
C3583 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VSS 0.982f 
C3584 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].VOUT VSS 0.862f 
C3585 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VSS 1.04f 
C3586 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS 0.627f 
C3587 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS 1.07f 
C3588 5_bit_dac_0[0].4_bit_dac_0[1].switch_n_3v3_0.D2 VSS 1.86f 
C3589 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ VSS 1.08f 
C3590 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 VSS 1.61f 
C3591 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS 1.06f 
C3592 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 VSS 3.25f 
C3593 a_1556_9002# VSS 1.16f 
C3594 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS 0.663f 
C3595 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS 0.467f 
C3596 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS 1.42f 
C3597 5_bit_dac_0[0].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH VSS 0.543f 
C3598 5_bit_dac_0[0].VOUT VSS 2.63f 
C3599 VOUT VSS 0.442f
C3600 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS 0.633f 
C3601 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS 1.08f 
C3602 D5_BUF VSS 8.89f
C3603 switch_n_3v3_0.DX_ VSS 1.09f 
C3604 D5 VSS 9.87f
C3605 5_bit_dac_0[0].D1 VSS 1.61f 
C3606 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS 1.06f 
C3607 5_bit_dac_0[0].D0 VSS 3.25f 
C3608 a_1556_10230# VSS 1.16f 
C3609 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS 0.663f 
C3610 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS 0.467f 
C3611 5_bit_dac_0[1].VREFH VSS 1.42f 
C3612 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH VSS 0.543f 
C3613 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS 1.02f 
C3614 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VSS 1.02f 
C3615 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS 0.627f 
C3616 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS 1.07f 
C3617 switch_n_3v3_0.D2 VSS 1.86f 
C3618 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].switch_n_3v3_1.DX_ VSS 1.08f 
C3619 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D1 VSS 1.61f 
C3620 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS 1.06f 
C3621 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[0].D0 VSS 3.25f 
C3622 a_1556_11458# VSS 1.16f 
C3623 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS 0.663f 
C3624 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS 0.467f 
C3625 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS 1.42f 
C3626 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH VSS 0.543f 
C3627 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].VOUT VSS 0.872f 
C3628 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS 0.633f 
C3629 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS 1.07f 
C3630 switch_n_3v3_0.D3 VSS 3.39f 
C3631 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.DX_ VSS 1.08f 
C3632 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D1 VSS 1.61f 
C3633 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS 1.06f 
C3634 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[0].D0 VSS 3.25f 
C3635 a_1556_12686# VSS 1.16f 
C3636 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS 0.663f 
C3637 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS 0.467f 
C3638 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VREFH VSS 1.42f 
C3639 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH VSS 0.543f 
C3640 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VSS 0.981f 
C3641 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].VOUT VSS 0.848f 
C3642 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VSS 0.984f 
C3643 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS 0.627f 
C3644 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS 1.07f 
C3645 5_bit_dac_0[1].4_bit_dac_0[0].switch_n_3v3_0.D2 VSS 1.86f 
C3646 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].switch_n_3v3_1.DX_ VSS 1.08f 
C3647 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D1 VSS 1.61f 
C3648 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS 1.06f 
C3649 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[0].D0 VSS 3.25f 
C3650 a_1556_13914# VSS 1.16f 
C3651 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS 0.663f 
C3652 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS 0.467f 
C3653 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS 1.42f 
C3654 5_bit_dac_0[1].4_bit_dac_0[0].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH VSS 0.543f 
C3655 5_bit_dac_0[1].4_bit_dac_0[0].VOUT VSS 1.22f 
C3656 5_bit_dac_0[1].VOUT VSS 2.38f 
C3657 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS 0.633f 
C3658 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS 1.08f 
C3659 switch_n_3v3_0.D4 VSS 7.7f 
C3660 5_bit_dac_0[1].switch_n_3v3_0.DX_ VSS 1.09f 
C3661 D4 VSS 2.71f
C3662 5_bit_dac_0[1].4_bit_dac_0[0].D1 VSS 1.61f 
C3663 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS 1.06f 
C3664 5_bit_dac_0[1].4_bit_dac_0[0].D0 VSS 3.25f 
C3665 a_1556_15142# VSS 1.16f 
C3666 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS 0.663f 
C3667 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS 0.467f 
C3668 5_bit_dac_0[1].4_bit_dac_0[1].VREFH VSS 1.42f 
C3669 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].switch2n_3v3_0.VREFH VSS 0.543f 
C3670 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].VOUT VSS 1.02f 
C3671 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VOUT VSS 1.02f 
C3672 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS 0.627f 
C3673 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS 1.07f 
C3674 5_bit_dac_0[1].switch_n_3v3_0.D2 VSS 1.86f 
C3675 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].switch_n_3v3_1.DX_ VSS 1.08f 
C3676 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D1 VSS 1.61f 
C3677 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS 1.06f 
C3678 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[0].D0 VSS 3.25f 
C3679 a_1556_16370# VSS 1.16f 
C3680 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS 0.663f 
C3681 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS 0.467f 
C3682 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].VREFH VSS 1.42f 
C3683 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].2_bit_dac_0[1].switch2n_3v3_0.VREFH VSS 0.543f 
C3684 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].VOUT VSS 0.864f 
C3685 5_bit_dac_0[1].4_bit_dac_0[1].VOUT VSS 1.73f 
C3686 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTH VSS 0.633f 
C3687 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VOUTL VSS 1.07f 
C3688 5_bit_dac_0[1].switch_n_3v3_0.D3 VSS 1.89f 
C3689 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.DX_ VSS 1.08f 
C3690 D3 VSS 0.641f
C3691 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D1 VSS 1.61f 
C3692 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch_n_3v3_v2_0.DX_ VSS 1.06f 
C3693 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[0].D0 VSS 3.25f 
C3694 a_1556_17598# VSS 1.16f 
C3695 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_L VSS 0.663f 
C3696 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.R_H VSS 0.467f 
C3697 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VREFH VSS 1.42f 
C3698 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].switch2n_3v3_0.VREFH VSS 0.543f 
C3699 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].VOUT VSS 0.984f 
C3700 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].VOUT VSS 0.923f 
C3701 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VOUT VSS 1.36f 
C3702 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTH VSS 0.905f 
C3703 VREFL VSS 1.15f
C3704 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VOUTL VSS 1.11f 
C3705 5_bit_dac_0[1].4_bit_dac_0[1].switch_n_3v3_0.D2 VSS 1.86f 
C3706 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].switch_n_3v3_1.DX_ VSS 1.1f 
C3707 D2 VSS 0.59f
C3708 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D1 VSS 1.61f 
C3709 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch_n_3v3_v2_0.DX_ VSS 1.08f 
C3710 D1 VSS 0.48f
C3711 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[0].D0 VSS 3.35f 
C3712 a_1556_18826# VSS 1.18f 
C3713 D0 VSS 0.729f
C3714 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_L VSS 0.68f 
C3715 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.R_H VSS 0.521f 
C3716 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].VREFH VSS 1.42f 
C3717 5_bit_dac_0[1].4_bit_dac_0[1].3_bit_dac_0[1].2_bit_dac_0[1].switch2n_3v3_0.VREFH VSS 0.714f 
C3718 VCC VSS 0.185p
C3719 D5.t1 VSS 0.33f 
C3720 D5.t0 VSS 0.189f 
C3721 D5.n0 VSS 0.362f 
C3722 D4.t1 VSS 0.145f 
C3723 D4.t0 VSS 0.0828f 
C3724 D4.n0 VSS 0.159f 
C3725 D4_BUF.t1 VSS 0.038f 
C3726 D4_BUF.t0 VSS 0.0226f 
C3727 D4_BUF.n0 VSS 0.283f 
C3728 D4_BUF.t3 VSS 0.115f 
C3729 D4_BUF.t2 VSS 0.0568f 
C3730 D4_BUF.n1 VSS 0.119f 
C3731 D4_BUF.n2 VSS 0.221f 
C3732 switch_n_3v3_0.D3.n0 VSS 0.44f 
C3733 switch_n_3v3_0.D3.t1 VSS 0.0332f 
C3734 switch_n_3v3_0.D3.t0 VSS 0.0197f 
C3735 switch_n_3v3_0.D3.t3 VSS 0.101f 
C3736 switch_n_3v3_0.D3.t4 VSS 0.0496f 
C3737 switch_n_3v3_0.D3.n1 VSS 0.104f 
C3738 switch_n_3v3_0.D3.t2 VSS 0.0961f 
C3739 switch_n_3v3_0.D3.t5 VSS 0.0549f 
C3740 switch_n_3v3_0.D3.n2 VSS 0.105f 
C3741 D5_BUF.t1 VSS 0.0979f 
C3742 D5_BUF.t0 VSS 0.0581f 
C3743 D5_BUF.n0 VSS 0.728f 
C3744 D5_BUF.t2 VSS 0.297f 
C3745 D5_BUF.t3 VSS 0.146f 
C3746 D5_BUF.n1 VSS 0.307f 
C3747 D5_BUF.n2 VSS 0.568f 
C3748 switch_n_3v3_0.D4.n0 VSS 0.881f 
C3749 switch_n_3v3_0.D4.t1 VSS 0.0665f 
C3750 switch_n_3v3_0.D4.t0 VSS 0.0395f 
C3751 switch_n_3v3_0.D4.t5 VSS 0.202f 
C3752 switch_n_3v3_0.D4.t2 VSS 0.0994f 
C3753 switch_n_3v3_0.D4.n1 VSS 0.209f 
C3754 switch_n_3v3_0.D4.t4 VSS 0.192f 
C3755 switch_n_3v3_0.D4.t3 VSS 0.11f 
C3756 switch_n_3v3_0.D4.n2 VSS 0.211f 
C3757 VCC.n0 VSS 5.76e-20 
C3758 VCC.n1 VSS 2.88e-20 
C3759 VCC.n2 VSS 3.5e-20 
C3760 VCC.n3 VSS 3.42e-20 
C3761 VCC.n4 VSS 3.5e-20 
C3762 VCC.n5 VSS 4.53e-19 
C3763 VCC.n6 VSS 1.17e-19 
C3764 VCC.n7 VSS 3.5e-20 
C3765 VCC.n8 VSS 1.44e-20 
C3766 VCC.n9 VSS 4.12e-20 
C3767 VCC.n10 VSS 5.76e-20 
C3768 VCC.t36 VSS 1.56e-19 
C3769 VCC.n11 VSS 7.62e-19 
C3770 VCC.n12 VSS 1.23e-20 
C3771 VCC.n13 VSS 5.76e-20 
C3772 VCC.n14 VSS 2.06e-20 
C3773 VCC.n15 VSS 3.29e-20 
C3774 VCC.n16 VSS 7.2e-20 
C3775 VCC.n17 VSS 3.29e-20 
C3776 VCC.n18 VSS 4.73e-20 
C3777 VCC.n19 VSS 2.26e-20 
C3778 VCC.n20 VSS 1.01e-19 
C3779 VCC.n21 VSS 1.36e-19 
C3780 VCC.n22 VSS 1.35e-19 
C3781 VCC.n23 VSS 3.5e-20 
C3782 VCC.n24 VSS 3.5e-20 
C3783 VCC.n25 VSS 3.5e-20 
C3784 VCC.n26 VSS 3.5e-20 
C3785 VCC.n27 VSS 3.09e-20 
C3786 VCC.n28 VSS 3.91e-20 
C3787 VCC.n29 VSS 4.73e-20 
C3788 VCC.n30 VSS 4.32e-20 
C3789 VCC.n31 VSS 2.68e-20 
C3790 VCC.n32 VSS 4.53e-20 
C3791 VCC.n33 VSS 4.53e-20 
C3792 VCC.n34 VSS 3.09e-20 
C3793 VCC.n35 VSS 4.32e-20 
C3794 VCC.n36 VSS 2.68e-20 
C3795 VCC.n37 VSS 7.82e-20 
C3796 VCC.n38 VSS 5.56e-20 
C3797 VCC.n39 VSS 1.4e-19 
C3798 VCC.n40 VSS 2.18e-19 
C3799 VCC.n41 VSS 1.35e-19 
C3800 VCC.n42 VSS 1.13e-19 
C3801 VCC.n43 VSS 3.5e-20 
C3802 VCC.n44 VSS 1.85e-20 
C3803 VCC.n45 VSS 3.7e-20 
C3804 VCC.n46 VSS 3.09e-20 
C3805 VCC.n47 VSS 6.59e-20 
C3806 VCC.n48 VSS 2.68e-20 
C3807 VCC.n49 VSS 5.76e-20 
C3808 VCC.n50 VSS 4.73e-20 
C3809 VCC.n51 VSS 3.5e-20 
C3810 VCC.t253 VSS 1.56e-19 
C3811 VCC.n52 VSS 7.97e-19 
C3812 VCC.n53 VSS 3.09e-20 
C3813 VCC.n54 VSS 3.5e-20 
C3814 VCC.n55 VSS 3.5e-20 
C3815 VCC.t252 VSS 4.21e-19 
C3816 VCC.n56 VSS 1.32e-19 
C3817 VCC.n57 VSS 1.09e-19 
C3818 VCC.n58 VSS 3.5e-20 
C3819 VCC.n59 VSS 3.09e-20 
C3820 VCC.n60 VSS 5.97e-20 
C3821 VCC.n61 VSS 2.26e-20 
C3822 VCC.n62 VSS 5.76e-20 
C3823 VCC.n63 VSS 2.68e-20 
C3824 VCC.n64 VSS 2.68e-20 
C3825 VCC.n65 VSS 1.9e-19 
C3826 VCC.n66 VSS 5.76e-20 
C3827 VCC.n67 VSS 2.68e-20 
C3828 VCC.n68 VSS 2.68e-20 
C3829 VCC.n69 VSS 2.68e-20 
C3830 VCC.n70 VSS 5.76e-20 
C3831 VCC.n71 VSS 2.26e-20 
C3832 VCC.n72 VSS 3.09e-20 
C3833 VCC.n73 VSS 2.26e-20 
C3834 VCC.n74 VSS 5.15e-20 
C3835 VCC.n75 VSS 4.73e-20 
C3836 VCC.n76 VSS 3.7e-20 
C3837 VCC.n77 VSS 3.5e-20 
C3838 VCC.n78 VSS 7.41e-20 
C3839 VCC.n79 VSS 1.91e-19 
C3840 VCC.n80 VSS 9.88e-20 
C3841 VCC.n81 VSS 3e-20 
C3842 VCC.n82 VSS 5.12e-19 
C3843 VCC.n83 VSS 1.18e-19 
C3844 VCC.n84 VSS 3.5e-20 
C3845 VCC.n85 VSS 3.5e-20 
C3846 VCC.n86 VSS 5.15e-20 
C3847 VCC.n87 VSS 4.32e-20 
C3848 VCC.n88 VSS 2.68e-20 
C3849 VCC.n89 VSS 3.91e-20 
C3850 VCC.n90 VSS 1.44e-20 
C3851 VCC.n91 VSS 3.5e-20 
C3852 VCC.n92 VSS 3e-20 
C3853 VCC.n93 VSS 7.95e-19 
C3854 VCC.n94 VSS 1.83e-19 
C3855 VCC.n95 VSS 2.88e-20 
C3856 VCC.n96 VSS 2.68e-20 
C3857 VCC.n97 VSS 2.68e-20 
C3858 VCC.n98 VSS 2.68e-20 
C3859 VCC.n99 VSS 4.53e-20 
C3860 VCC.n100 VSS 3.7e-20 
C3861 VCC.n101 VSS 7.82e-20 
C3862 VCC.n102 VSS 1.17e-19 
C3863 VCC.n103 VSS 3.91e-20 
C3864 VCC.n104 VSS 1.65e-20 
C3865 VCC.n105 VSS 2.68e-20 
C3866 VCC.n106 VSS 3.5e-20 
C3867 VCC.n107 VSS 3e-20 
C3868 VCC.n108 VSS 5.12e-19 
C3869 VCC.n109 VSS 1.18e-19 
C3870 VCC.n110 VSS 3.5e-20 
C3871 VCC.n111 VSS 3.5e-20 
C3872 VCC.t249 VSS 1.55e-19 
C3873 VCC.n112 VSS 7.57e-19 
C3874 VCC.n113 VSS 4.73e-20 
C3875 VCC.n114 VSS 1.54e-19 
C3876 VCC.n115 VSS 2.88e-20 
C3877 VCC.n116 VSS 2.88e-20 
C3878 VCC.n117 VSS 3.5e-20 
C3879 VCC.n118 VSS 5.76e-20 
C3880 VCC.n119 VSS 9.88e-20 
C3881 VCC.n120 VSS 1.3e-19 
C3882 VCC.n121 VSS 3e-20 
C3883 VCC.t250 VSS 0.005f 
C3884 VCC.t211 VSS 0.00453f 
C3885 VCC.n122 VSS 0.00229f 
C3886 VCC.n123 VSS 1.91e-19 
C3887 VCC.n124 VSS 3.5e-20 
C3888 VCC.n125 VSS 3.14e-19 
C3889 VCC.n126 VSS 2.47e-20 
C3890 VCC.n127 VSS 5.76e-20 
C3891 VCC.n128 VSS 2.47e-20 
C3892 VCC.n129 VSS 8.23e-21 
C3893 VCC.n130 VSS 2.88e-20 
C3894 VCC.n131 VSS 5.76e-20 
C3895 VCC.n132 VSS 2.47e-20 
C3896 VCC.n133 VSS 2.88e-20 
C3897 VCC.n134 VSS 2.47e-20 
C3898 VCC.n135 VSS 5.15e-20 
C3899 VCC.n136 VSS 4.73e-20 
C3900 VCC.n137 VSS 3.7e-20 
C3901 VCC.n138 VSS 3.5e-20 
C3902 VCC.n139 VSS 7.41e-20 
C3903 VCC.t289 VSS 6.42e-19 
C3904 VCC.n140 VSS 3e-20 
C3905 VCC.n141 VSS 5.97e-20 
C3906 VCC.n142 VSS 4.13e-19 
C3907 VCC.n143 VSS 9.53e-20 
C3908 VCC.n144 VSS 3.5e-20 
C3909 VCC.n145 VSS 3.5e-20 
C3910 VCC.n146 VSS 5.35e-20 
C3911 VCC.n147 VSS 4.32e-20 
C3912 VCC.n148 VSS 2.68e-20 
C3913 VCC.n149 VSS 3.7e-20 
C3914 VCC.n150 VSS 1.65e-20 
C3915 VCC.n151 VSS 4.53e-20 
C3916 VCC.n152 VSS 1.2e-19 
C3917 VCC.n153 VSS 5.2e-19 
C3918 VCC.n154 VSS 1.2e-19 
C3919 VCC.n155 VSS 6.38e-20 
C3920 VCC.n156 VSS 2.47e-20 
C3921 VCC.n157 VSS 4.53e-20 
C3922 VCC.n158 VSS 3.5e-20 
C3923 VCC.n159 VSS 3.5e-20 
C3924 VCC.n160 VSS 2.68e-20 
C3925 VCC.n161 VSS 2.68e-20 
C3926 VCC.n162 VSS 2.47e-20 
C3927 VCC.n163 VSS 4.53e-20 
C3928 VCC.n164 VSS 2.68e-20 
C3929 VCC.n165 VSS 4.32e-20 
C3930 VCC.n166 VSS 2.68e-20 
C3931 VCC.n167 VSS 3.91e-20 
C3932 VCC.n168 VSS 2.88e-20 
C3933 VCC.n169 VSS 4.73e-20 
C3934 VCC.n170 VSS 3.7e-20 
C3935 VCC.n171 VSS 3.7e-20 
C3936 VCC.n172 VSS 3.5e-20 
C3937 VCC.n173 VSS 5.76e-20 
C3938 VCC.n174 VSS 4.73e-20 
C3939 VCC.n175 VSS 3.09e-20 
C3940 VCC.n176 VSS 3.5e-20 
C3941 VCC.n177 VSS 3.5e-20 
C3942 VCC.n178 VSS 3.5e-20 
C3943 VCC.n179 VSS 1.18e-19 
C3944 VCC.n180 VSS 3e-20 
C3945 VCC.n181 VSS 1.15e-19 
C3946 VCC.n182 VSS 9.88e-20 
C3947 VCC.n183 VSS 5.76e-20 
C3948 VCC.n184 VSS 3.5e-20 
C3949 VCC.n185 VSS 3.09e-20 
C3950 VCC.n186 VSS 3.09e-20 
C3951 VCC.n187 VSS 2.26e-20 
C3952 VCC.n188 VSS 5.76e-20 
C3953 VCC.n189 VSS 2.68e-20 
C3954 VCC.n190 VSS 2.68e-20 
C3955 VCC.n191 VSS 0.00185f 
C3956 VCC.n192 VSS 2.72e-19 
C3957 VCC.n193 VSS 2.26e-20 
C3958 VCC.n194 VSS 1.87e-19 
C3959 VCC.n195 VSS 3.5e-20 
C3960 VCC.n196 VSS 2.68e-20 
C3961 VCC.n197 VSS 5.97e-20 
C3962 VCC.n198 VSS 4.73e-20 
C3963 VCC.n199 VSS 4.73e-20 
C3964 VCC.n200 VSS 5.15e-20 
C3965 VCC.n201 VSS 7.41e-20 
C3966 VCC.n202 VSS 3.7e-20 
C3967 VCC.n203 VSS 2.26e-20 
C3968 VCC.n204 VSS 6.38e-20 
C3969 VCC.n205 VSS 4.73e-20 
C3970 VCC.n206 VSS 3.29e-20 
C3971 VCC.n207 VSS 3.5e-20 
C3972 VCC.n208 VSS 3e-20 
C3973 VCC.t261 VSS 0.005f 
C3974 VCC.t151 VSS 0.00453f 
C3975 VCC.n209 VSS 0.00228f 
C3976 VCC.n210 VSS 1.3e-19 
C3977 VCC.t262 VSS 4.05e-19 
C3978 VCC.n211 VSS 4.05e-19 
C3979 VCC.n212 VSS 1.15e-19 
C3980 VCC.n213 VSS 3.36e-19 
C3981 VCC.n214 VSS 6.17e-21 
C3982 VCC.n215 VSS 3.12e-19 
C3983 VCC.n216 VSS 1.65e-20 
C3984 VCC.n217 VSS 1.54e-19 
C3985 VCC.n218 VSS 1.54e-19 
C3986 VCC.n219 VSS 1.65e-20 
C3987 VCC.n220 VSS 1.03e-20 
C3988 VCC.n221 VSS 3.5e-20 
C3989 VCC.n222 VSS 2.26e-20 
C3990 VCC.n223 VSS 4.73e-20 
C3991 VCC.n224 VSS 3.5e-20 
C3992 VCC.n225 VSS 3e-20 
C3993 VCC.n226 VSS 1.3e-19 
C3994 VCC.n227 VSS 5.12e-19 
C3995 VCC.n228 VSS 1.3e-19 
C3996 VCC.n229 VSS 4.13e-19 
C3997 VCC.n230 VSS 9.53e-20 
C3998 VCC.n231 VSS 5.76e-20 
C3999 VCC.n232 VSS 7.41e-20 
C4000 VCC.n233 VSS 5.56e-20 
C4001 VCC.t263 VSS 1.55e-19 
C4002 VCC.n234 VSS 3.91e-20 
C4003 VCC.n235 VSS 3.91e-20 
C4004 VCC.n236 VSS 1.85e-20 
C4005 VCC.n237 VSS 7.55e-19 
C4006 VCC.n238 VSS 4.94e-20 
C4007 VCC.n239 VSS 5.15e-20 
C4008 VCC.n240 VSS 7.2e-20 
C4009 VCC.n241 VSS 1.38e-19 
C4010 VCC.n242 VSS 1.17e-19 
C4011 VCC.n243 VSS 4.32e-20 
C4012 VCC.n244 VSS 2.88e-20 
C4013 VCC.n245 VSS 2.68e-20 
C4014 VCC.n246 VSS 3.5e-20 
C4015 VCC.n247 VSS 3.5e-20 
C4016 VCC.n248 VSS 2.88e-20 
C4017 VCC.n249 VSS 2.68e-20 
C4018 VCC.n250 VSS 2.68e-20 
C4019 VCC.n251 VSS 2.68e-20 
C4020 VCC.n252 VSS 4.12e-20 
C4021 VCC.n253 VSS 4.12e-20 
C4022 VCC.n254 VSS 3.91e-20 
C4023 VCC.n255 VSS 4.53e-20 
C4024 VCC.n256 VSS 4.53e-20 
C4025 VCC.n257 VSS 1.05e-19 
C4026 VCC.n258 VSS 1.05e-19 
C4027 VCC.n259 VSS 4.32e-20 
C4028 VCC.n260 VSS 3.7e-20 
C4029 VCC.n261 VSS 2.68e-20 
C4030 VCC.n262 VSS 2.68e-20 
C4031 VCC.n263 VSS 6.79e-20 
C4032 VCC.n264 VSS 9.26e-20 
C4033 VCC.n265 VSS 1.83e-19 
C4034 VCC.n266 VSS 7.95e-19 
C4035 VCC.n267 VSS 5.2e-19 
C4036 VCC.n268 VSS 1.3e-19 
C4037 VCC.n269 VSS 3e-20 
C4038 VCC.n270 VSS 3.5e-20 
C4039 VCC.n271 VSS 5.97e-20 
C4040 VCC.n272 VSS 7.41e-20 
C4041 VCC.n273 VSS 5.15e-20 
C4042 VCC.n274 VSS 5.15e-20 
C4043 VCC.n275 VSS 3.09e-20 
C4044 VCC.n276 VSS 3.09e-20 
C4045 VCC.n277 VSS 3.7e-20 
C4046 VCC.n278 VSS 2.68e-20 
C4047 VCC.n279 VSS 3.91e-20 
C4048 VCC.n280 VSS 1.17e-19 
C4049 VCC.n281 VSS 1.38e-19 
C4050 VCC.n282 VSS 7e-20 
C4051 VCC.n283 VSS 4.73e-20 
C4052 VCC.n284 VSS 3.5e-20 
C4053 VCC.n285 VSS 3.5e-20 
C4054 VCC.n286 VSS 3.5e-20 
C4055 VCC.n287 VSS 4.53e-20 
C4056 VCC.n288 VSS 1.18e-19 
C4057 VCC.n289 VSS 5.12e-19 
C4058 VCC.n290 VSS 1.3e-19 
C4059 VCC.n291 VSS 1.61e-19 
C4060 VCC.n292 VSS 9.9e-20 
C4061 VCC.n293 VSS 0.00243f 
C4062 VCC.n294 VSS 2.26e-20 
C4063 VCC.n295 VSS 4.13e-19 
C4064 VCC.n296 VSS 3.5e-20 
C4065 VCC.n297 VSS 3.5e-20 
C4066 VCC.n298 VSS 2.47e-20 
C4067 VCC.n299 VSS 2.06e-20 
C4068 VCC.n300 VSS 6.17e-20 
C4069 VCC.n301 VSS 6.17e-20 
C4070 VCC.n302 VSS 4.73e-20 
C4071 VCC.n303 VSS 4.73e-20 
C4072 VCC.n304 VSS 2.88e-20 
C4073 VCC.n305 VSS 1.44e-20 
C4074 VCC.n306 VSS 1.65e-20 
C4075 VCC.n307 VSS 1.54e-19 
C4076 VCC.n308 VSS 1.54e-19 
C4077 VCC.n309 VSS 1.65e-20 
C4078 VCC.n310 VSS 3.09e-20 
C4079 VCC.t290 VSS 1.55e-19 
C4080 VCC.n311 VSS 0.00102f 
C4081 VCC.n312 VSS 2.73e-19 
C4082 VCC.n313 VSS 0.00136f 
C4083 VCC.n314 VSS 2.73e-19 
C4084 VCC.n315 VSS 0.00181f 
C4085 VCC.n316 VSS 5.76e-20 
C4086 VCC.n317 VSS 1.54e-19 
C4087 VCC.n318 VSS 1.65e-20 
C4088 VCC.n319 VSS 2.88e-20 
C4089 VCC.n320 VSS 2.47e-20 
C4090 VCC.n321 VSS 6.17e-20 
C4091 VCC.n322 VSS 4.73e-20 
C4092 VCC.n323 VSS 4.73e-20 
C4093 VCC.n324 VSS 5.15e-20 
C4094 VCC.n325 VSS 3.5e-20 
C4095 VCC.n326 VSS 7.41e-20 
C4096 VCC.n327 VSS 3.7e-20 
C4097 VCC.n328 VSS 2.26e-20 
C4098 VCC.n329 VSS 6.17e-20 
C4099 VCC.n330 VSS 4.73e-20 
C4100 VCC.n331 VSS 3.5e-20 
C4101 VCC.n332 VSS 2.88e-20 
C4102 VCC.n333 VSS 3.4e-19 
C4103 VCC.n334 VSS 1.15e-19 
C4104 VCC.n335 VSS 3.98e-19 
C4105 VCC.t248 VSS 4.05e-19 
C4106 VCC.n336 VSS 1.22e-19 
C4107 VCC.n337 VSS 1.3e-19 
C4108 VCC.n338 VSS 3e-20 
C4109 VCC.n339 VSS 3.5e-20 
C4110 VCC.n340 VSS 3.5e-20 
C4111 VCC.n341 VSS 4.73e-20 
C4112 VCC.n342 VSS 2.47e-20 
C4113 VCC.n343 VSS 1.23e-20 
C4114 VCC.n344 VSS 1.65e-20 
C4115 VCC.n345 VSS 2.47e-20 
C4116 VCC.n346 VSS 5.76e-20 
C4117 VCC.n347 VSS 1.38e-19 
C4118 VCC.n348 VSS 7e-20 
C4119 VCC.n349 VSS 3.7e-20 
C4120 VCC.n350 VSS 2.47e-20 
C4121 VCC.n351 VSS 3.7e-20 
C4122 VCC.n352 VSS 1.85e-20 
C4123 VCC.n353 VSS 3.09e-20 
C4124 VCC.n354 VSS 5.35e-20 
C4125 VCC.n355 VSS 4.73e-20 
C4126 VCC.n356 VSS 5.35e-20 
C4127 VCC.n357 VSS 7.41e-20 
C4128 VCC.n358 VSS 5.76e-20 
C4129 VCC.n359 VSS 9.53e-20 
C4130 VCC.n360 VSS 4.13e-19 
C4131 VCC.n361 VSS 1.3e-19 
C4132 VCC.n362 VSS 5.2e-19 
C4133 VCC.n363 VSS 1.2e-19 
C4134 VCC.n364 VSS 4.73e-20 
C4135 VCC.n365 VSS 2.68e-20 
C4136 VCC.n366 VSS 3.5e-20 
C4137 VCC.n367 VSS 3.5e-20 
C4138 VCC.n368 VSS 2.68e-20 
C4139 VCC.n369 VSS 2.68e-20 
C4140 VCC.n370 VSS 4.32e-20 
C4141 VCC.n371 VSS 4.32e-20 
C4142 VCC.n372 VSS 4.32e-20 
C4143 VCC.n373 VSS 2.88e-20 
C4144 VCC.n374 VSS 3.5e-20 
C4145 VCC.n375 VSS 2.68e-20 
C4146 VCC.n376 VSS 7.82e-20 
C4147 VCC.n377 VSS 4.73e-20 
C4148 VCC.n378 VSS 4.73e-20 
C4149 VCC.n379 VSS 1.05e-19 
C4150 VCC.n380 VSS 1.05e-19 
C4151 VCC.n381 VSS 4.53e-20 
C4152 VCC.n382 VSS 2.68e-20 
C4153 VCC.n383 VSS 2.68e-20 
C4154 VCC.n384 VSS 6.59e-20 
C4155 VCC.n385 VSS 9.26e-20 
C4156 VCC.n386 VSS 6.59e-20 
C4157 VCC.n387 VSS 2.47e-20 
C4158 VCC.n388 VSS 2.47e-20 
C4159 VCC.n389 VSS 2.88e-20 
C4160 VCC.n390 VSS 3.5e-20 
C4161 VCC.n391 VSS 3.5e-20 
C4162 VCC.n392 VSS 4.53e-20 
C4163 VCC.n393 VSS 1.2e-19 
C4164 VCC.n394 VSS 5.2e-19 
C4165 VCC.n395 VSS 1.3e-19 
C4166 VCC.n396 VSS 4.13e-19 
C4167 VCC.n397 VSS 9.53e-20 
C4168 VCC.n398 VSS 5.97e-20 
C4169 VCC.n399 VSS 7.41e-20 
C4170 VCC.n400 VSS 5.35e-20 
C4171 VCC.n401 VSS 5.15e-20 
C4172 VCC.n402 VSS 3.09e-20 
C4173 VCC.n403 VSS 3.09e-20 
C4174 VCC.n404 VSS 3.91e-20 
C4175 VCC.n405 VSS 2.47e-20 
C4176 VCC.n406 VSS 3.7e-20 
C4177 VCC.n407 VSS 1.17e-19 
C4178 VCC.n408 VSS 1.38e-19 
C4179 VCC.n409 VSS 7.2e-20 
C4180 VCC.n410 VSS 4.73e-20 
C4181 VCC.n411 VSS 3.5e-20 
C4182 VCC.n412 VSS 3.5e-20 
C4183 VCC.n413 VSS 4.53e-20 
C4184 VCC.n414 VSS 5.97e-20 
C4185 VCC.n415 VSS 3.5e-20 
C4186 VCC.n416 VSS 3e-20 
C4187 VCC.n417 VSS 1.3e-19 
C4188 VCC.n418 VSS 1.53e-19 
C4189 VCC.t102 VSS 4.05e-19 
C4190 VCC.n419 VSS 2.06e-19 
C4191 VCC.n420 VSS 1.35e-19 
C4192 VCC.n421 VSS 9.67e-20 
C4193 VCC.n422 VSS 3.35e-20 
C4194 VCC.n423 VSS 3.5e-20 
C4195 VCC.n424 VSS 2.36e-19 
C4196 VCC.n425 VSS 0.0023f 
C4197 VCC.t251 VSS 0.0031f 
C4198 VCC.t283 VSS 0.00366f 
C4199 VCC.t254 VSS 0.00365f 
C4200 VCC.t282 VSS 0.00386f 
C4201 VCC.n426 VSS 0.00569f 
C4202 VCC.n427 VSS 1.3e-19 
C4203 VCC.n428 VSS 3.67e-19 
C4204 VCC.n429 VSS 1.15e-19 
C4205 VCC.n430 VSS 3.38e-19 
C4206 VCC.n431 VSS 3.5e-20 
C4207 VCC.n432 VSS 3.5e-20 
C4208 VCC.n433 VSS 2.68e-20 
C4209 VCC.n434 VSS 2.06e-20 
C4210 VCC.n435 VSS 6.38e-20 
C4211 VCC.n436 VSS 5.97e-20 
C4212 VCC.n437 VSS 4.73e-20 
C4213 VCC.n438 VSS 4.73e-20 
C4214 VCC.n439 VSS 3.09e-20 
C4215 VCC.n440 VSS 1.23e-20 
C4216 VCC.n441 VSS 1.65e-20 
C4217 VCC.n442 VSS 1.54e-19 
C4218 VCC.n443 VSS 1.54e-19 
C4219 VCC.n444 VSS 1.65e-20 
C4220 VCC.n445 VSS 3.29e-20 
C4221 VCC.t103 VSS 1.67e-19 
C4222 VCC.n446 VSS 0.00101f 
C4223 VCC.n447 VSS 2.71e-19 
C4224 VCC.n448 VSS 7.46e-19 
C4225 VCC.n449 VSS 0.00333f 
C4226 VCC.n450 VSS 2.46e-19 
C4227 VCC.n451 VSS 3.02e-19 
C4228 VCC.n452 VSS 3.7e-20 
C4229 VCC.n453 VSS 5.15e-20 
C4230 VCC.n454 VSS 6.38e-20 
C4231 VCC.n455 VSS 4.73e-20 
C4232 VCC.n456 VSS 4.73e-20 
C4233 VCC.n457 VSS 2.68e-20 
C4234 VCC.n458 VSS 3.29e-20 
C4235 VCC.n459 VSS 1.65e-20 
C4236 VCC.n460 VSS 1.54e-19 
C4237 VCC.n461 VSS 1.54e-19 
C4238 VCC.n462 VSS 5.56e-20 
C4239 VCC.n463 VSS 2.88e-20 
C4240 VCC.n464 VSS 1.65e-20 
C4241 VCC.n465 VSS 3.09e-20 
C4242 VCC.n466 VSS 4.73e-20 
C4243 VCC.n467 VSS 4.73e-20 
C4244 VCC.n468 VSS 4.32e-20 
C4245 VCC.n469 VSS 1.17e-19 
C4246 VCC.n470 VSS 3.33e-19 
C4247 VCC.n471 VSS 1.35e-19 
C4248 VCC.n472 VSS 4.37e-19 
C4249 VCC.n473 VSS 5.24e-19 
C4250 VCC.n474 VSS 1.36e-19 
C4251 VCC.n475 VSS 1.01e-19 
C4252 VCC.n476 VSS 1.05e-19 
C4253 VCC.n477 VSS 2.06e-20 
C4254 VCC.n478 VSS 2.26e-20 
C4255 VCC.n479 VSS 3.7e-20 
C4256 VCC.n480 VSS 5.15e-20 
C4257 VCC.n481 VSS 1.38e-19 
C4258 VCC.n482 VSS 3.91e-20 
C4259 VCC.n483 VSS 2.88e-20 
C4260 VCC.n484 VSS 4.32e-20 
C4261 VCC.n485 VSS 1.17e-19 
C4262 VCC.n486 VSS 3.7e-20 
C4263 VCC.n487 VSS 3.91e-20 
C4264 VCC.n488 VSS 3.5e-20 
C4265 VCC.n489 VSS 1.65e-20 
C4266 VCC.n490 VSS 8.23e-21 
C4267 VCC.n491 VSS 3.5e-20 
C4268 VCC.n492 VSS 3.5e-20 
C4269 VCC.n493 VSS 1.4e-19 
C4270 VCC.n494 VSS 5.4e-19 
C4271 VCC.n495 VSS 8.42e-19 
C4272 VCC.n496 VSS 5.4e-19 
C4273 VCC.n497 VSS 1.4e-19 
C4274 VCC.n498 VSS 1.4e-19 
C4275 VCC.n499 VSS 2.18e-19 
C4276 VCC.n500 VSS 7.82e-20 
C4277 VCC.n501 VSS 4.32e-20 
C4278 VCC.n502 VSS 4.32e-20 
C4279 VCC.n503 VSS 1.05e-19 
C4280 VCC.n504 VSS 1.05e-19 
C4281 VCC.n505 VSS 4.32e-20 
C4282 VCC.n506 VSS 3.7e-20 
C4283 VCC.n507 VSS 2.68e-20 
C4284 VCC.n508 VSS 5.76e-20 
C4285 VCC.n509 VSS 6.38e-20 
C4286 VCC.n510 VSS 3.5e-20 
C4287 VCC.n511 VSS 3.5e-20 
C4288 VCC.n512 VSS 1.17e-19 
C4289 VCC.n513 VSS 1.38e-19 
C4290 VCC.n514 VSS 5.15e-20 
C4291 VCC.n515 VSS 1.05e-19 
C4292 VCC.n516 VSS 2.26e-20 
C4293 VCC.n517 VSS 5.76e-20 
C4294 VCC.n518 VSS 3.7e-20 
C4295 VCC.n519 VSS 3.7e-20 
C4296 VCC.n520 VSS 3.09e-20 
C4297 VCC.n521 VSS 1.85e-20 
C4298 VCC.n522 VSS 1.65e-20 
C4299 VCC.n523 VSS 8.23e-21 
C4300 VCC.n524 VSS 1.13e-19 
C4301 VCC.n525 VSS 3.33e-19 
C4302 VCC.t35 VSS 4.21e-19 
C4303 VCC.n526 VSS 2.06e-19 
C4304 VCC.n527 VSS 1.35e-19 
C4305 VCC.n528 VSS 3.5e-20 
C4306 VCC.n529 VSS 3.5e-20 
C4307 VCC.n530 VSS 3.5e-20 
C4308 VCC.n531 VSS 1.03e-20 
C4309 VCC.n532 VSS 2.68e-20 
C4310 VCC.n533 VSS 3.09e-20 
C4311 VCC.n534 VSS 2.68e-20 
C4312 VCC.n535 VSS 1.65e-20 
C4313 VCC.n536 VSS 1.54e-19 
C4314 VCC.n537 VSS 1.54e-19 
C4315 VCC.n538 VSS 1.65e-20 
C4316 VCC.n539 VSS 2.47e-20 
C4317 VCC.n540 VSS 4.73e-20 
C4318 VCC.n541 VSS 6.59e-20 
C4319 VCC.n542 VSS 5.15e-20 
C4320 VCC.n543 VSS 2.47e-20 
C4321 VCC.n544 VSS 7.41e-20 
C4322 VCC.n545 VSS 9.47e-20 
C4323 VCC.n546 VSS 1.32e-19 
C4324 VCC.n547 VSS 7.71e-19 
C4325 VCC.n548 VSS 9.83e-19 
C4326 VCC.n549 VSS 2.36e-19 
C4327 VCC.n550 VSS 3.21e-19 
C4328 VCC.n551 VSS 2.61e-19 
C4329 VCC.n552 VSS 0.00189f 
C4330 VCC.n553 VSS 5.37e-19 
C4331 VCC.n554 VSS 5.76e-20 
C4332 VCC.n555 VSS 2.88e-20 
C4333 VCC.n556 VSS 3.5e-20 
C4334 VCC.n557 VSS 3.42e-20 
C4335 VCC.n558 VSS 3.5e-20 
C4336 VCC.n559 VSS 4.53e-19 
C4337 VCC.n560 VSS 1.17e-19 
C4338 VCC.n561 VSS 3.5e-20 
C4339 VCC.n562 VSS 1.44e-20 
C4340 VCC.n563 VSS 4.12e-20 
C4341 VCC.n564 VSS 5.76e-20 
C4342 VCC.n565 VSS 5.76e-20 
C4343 VCC.n566 VSS 2.06e-20 
C4344 VCC.n567 VSS 3.29e-20 
C4345 VCC.n568 VSS 7.2e-20 
C4346 VCC.n569 VSS 3.29e-20 
C4347 VCC.n570 VSS 4.73e-20 
C4348 VCC.n571 VSS 2.26e-20 
C4349 VCC.n572 VSS 1.01e-19 
C4350 VCC.n573 VSS 1.36e-19 
C4351 VCC.n574 VSS 1.35e-19 
C4352 VCC.n575 VSS 3.5e-20 
C4353 VCC.n576 VSS 3.5e-20 
C4354 VCC.n577 VSS 3.5e-20 
C4355 VCC.n578 VSS 3.5e-20 
C4356 VCC.n579 VSS 3.09e-20 
C4357 VCC.n580 VSS 3.91e-20 
C4358 VCC.n581 VSS 4.73e-20 
C4359 VCC.n582 VSS 4.32e-20 
C4360 VCC.n583 VSS 2.68e-20 
C4361 VCC.n584 VSS 4.53e-20 
C4362 VCC.n585 VSS 4.53e-20 
C4363 VCC.n586 VSS 3.09e-20 
C4364 VCC.n587 VSS 4.32e-20 
C4365 VCC.n588 VSS 2.68e-20 
C4366 VCC.n589 VSS 7.82e-20 
C4367 VCC.n590 VSS 5.56e-20 
C4368 VCC.n591 VSS 1.4e-19 
C4369 VCC.n592 VSS 2.18e-19 
C4370 VCC.n593 VSS 1.35e-19 
C4371 VCC.n594 VSS 1.13e-19 
C4372 VCC.n595 VSS 3.5e-20 
C4373 VCC.n596 VSS 1.85e-20 
C4374 VCC.n597 VSS 3.7e-20 
C4375 VCC.n598 VSS 3.09e-20 
C4376 VCC.n599 VSS 6.59e-20 
C4377 VCC.n600 VSS 2.68e-20 
C4378 VCC.n601 VSS 5.76e-20 
C4379 VCC.n602 VSS 4.73e-20 
C4380 VCC.n603 VSS 3.5e-20 
C4381 VCC.t30 VSS 1.56e-19 
C4382 VCC.n604 VSS 7.97e-19 
C4383 VCC.n605 VSS 3.09e-20 
C4384 VCC.n606 VSS 3.5e-20 
C4385 VCC.n607 VSS 3.5e-20 
C4386 VCC.t29 VSS 4.21e-19 
C4387 VCC.n608 VSS 1.32e-19 
C4388 VCC.n609 VSS 1.09e-19 
C4389 VCC.n610 VSS 3.5e-20 
C4390 VCC.n611 VSS 3.09e-20 
C4391 VCC.n612 VSS 5.97e-20 
C4392 VCC.n613 VSS 2.26e-20 
C4393 VCC.n614 VSS 5.76e-20 
C4394 VCC.n615 VSS 2.68e-20 
C4395 VCC.n616 VSS 2.68e-20 
C4396 VCC.n617 VSS 1.9e-19 
C4397 VCC.n618 VSS 5.76e-20 
C4398 VCC.n619 VSS 2.68e-20 
C4399 VCC.n620 VSS 2.68e-20 
C4400 VCC.n621 VSS 2.68e-20 
C4401 VCC.n622 VSS 5.76e-20 
C4402 VCC.n623 VSS 2.26e-20 
C4403 VCC.n624 VSS 3.09e-20 
C4404 VCC.n625 VSS 2.26e-20 
C4405 VCC.n626 VSS 5.15e-20 
C4406 VCC.n627 VSS 4.73e-20 
C4407 VCC.n628 VSS 3.7e-20 
C4408 VCC.n629 VSS 3.5e-20 
C4409 VCC.n630 VSS 7.41e-20 
C4410 VCC.n631 VSS 1.91e-19 
C4411 VCC.n632 VSS 9.88e-20 
C4412 VCC.n633 VSS 3e-20 
C4413 VCC.n634 VSS 5.12e-19 
C4414 VCC.n635 VSS 1.18e-19 
C4415 VCC.n636 VSS 3.5e-20 
C4416 VCC.n637 VSS 3.5e-20 
C4417 VCC.n638 VSS 5.15e-20 
C4418 VCC.n639 VSS 4.32e-20 
C4419 VCC.n640 VSS 2.68e-20 
C4420 VCC.n641 VSS 3.91e-20 
C4421 VCC.n642 VSS 1.44e-20 
C4422 VCC.n643 VSS 3.5e-20 
C4423 VCC.n644 VSS 3e-20 
C4424 VCC.n645 VSS 7.95e-19 
C4425 VCC.n646 VSS 1.83e-19 
C4426 VCC.n647 VSS 2.88e-20 
C4427 VCC.n648 VSS 2.68e-20 
C4428 VCC.n649 VSS 2.68e-20 
C4429 VCC.n650 VSS 2.68e-20 
C4430 VCC.n651 VSS 4.53e-20 
C4431 VCC.n652 VSS 3.7e-20 
C4432 VCC.n653 VSS 7.82e-20 
C4433 VCC.n654 VSS 1.17e-19 
C4434 VCC.n655 VSS 3.91e-20 
C4435 VCC.n656 VSS 1.65e-20 
C4436 VCC.n657 VSS 2.68e-20 
C4437 VCC.n658 VSS 3.5e-20 
C4438 VCC.n659 VSS 3e-20 
C4439 VCC.n660 VSS 5.12e-19 
C4440 VCC.n661 VSS 1.18e-19 
C4441 VCC.n662 VSS 3.5e-20 
C4442 VCC.n663 VSS 3.5e-20 
C4443 VCC.t106 VSS 1.55e-19 
C4444 VCC.n664 VSS 7.57e-19 
C4445 VCC.n665 VSS 4.73e-20 
C4446 VCC.n666 VSS 1.54e-19 
C4447 VCC.n667 VSS 2.88e-20 
C4448 VCC.n668 VSS 2.88e-20 
C4449 VCC.n669 VSS 3.5e-20 
C4450 VCC.n670 VSS 5.76e-20 
C4451 VCC.n671 VSS 9.88e-20 
C4452 VCC.n672 VSS 1.3e-19 
C4453 VCC.n673 VSS 3e-20 
C4454 VCC.t104 VSS 0.005f 
C4455 VCC.t257 VSS 0.00453f 
C4456 VCC.n674 VSS 0.00229f 
C4457 VCC.n675 VSS 1.91e-19 
C4458 VCC.n676 VSS 3.5e-20 
C4459 VCC.n677 VSS 3.14e-19 
C4460 VCC.n678 VSS 2.47e-20 
C4461 VCC.n679 VSS 5.76e-20 
C4462 VCC.n680 VSS 2.47e-20 
C4463 VCC.n681 VSS 8.23e-21 
C4464 VCC.n682 VSS 2.88e-20 
C4465 VCC.n683 VSS 5.76e-20 
C4466 VCC.n684 VSS 2.47e-20 
C4467 VCC.n685 VSS 2.88e-20 
C4468 VCC.n686 VSS 2.47e-20 
C4469 VCC.n687 VSS 5.15e-20 
C4470 VCC.n688 VSS 4.73e-20 
C4471 VCC.n689 VSS 3.7e-20 
C4472 VCC.n690 VSS 3.5e-20 
C4473 VCC.n691 VSS 7.41e-20 
C4474 VCC.t235 VSS 6.42e-19 
C4475 VCC.n692 VSS 3e-20 
C4476 VCC.n693 VSS 5.97e-20 
C4477 VCC.n694 VSS 4.13e-19 
C4478 VCC.n695 VSS 9.53e-20 
C4479 VCC.n696 VSS 3.5e-20 
C4480 VCC.n697 VSS 3.5e-20 
C4481 VCC.n698 VSS 5.35e-20 
C4482 VCC.n699 VSS 4.32e-20 
C4483 VCC.n700 VSS 2.68e-20 
C4484 VCC.n701 VSS 3.7e-20 
C4485 VCC.n702 VSS 1.65e-20 
C4486 VCC.n703 VSS 4.53e-20 
C4487 VCC.n704 VSS 1.2e-19 
C4488 VCC.n705 VSS 5.2e-19 
C4489 VCC.n706 VSS 1.2e-19 
C4490 VCC.n707 VSS 6.38e-20 
C4491 VCC.n708 VSS 2.47e-20 
C4492 VCC.n709 VSS 4.53e-20 
C4493 VCC.n710 VSS 3.5e-20 
C4494 VCC.n711 VSS 3.5e-20 
C4495 VCC.n712 VSS 2.68e-20 
C4496 VCC.n713 VSS 2.68e-20 
C4497 VCC.n714 VSS 2.47e-20 
C4498 VCC.n715 VSS 4.53e-20 
C4499 VCC.n716 VSS 2.68e-20 
C4500 VCC.n717 VSS 4.32e-20 
C4501 VCC.n718 VSS 2.68e-20 
C4502 VCC.n719 VSS 3.91e-20 
C4503 VCC.n720 VSS 2.88e-20 
C4504 VCC.n721 VSS 4.73e-20 
C4505 VCC.n722 VSS 3.7e-20 
C4506 VCC.n723 VSS 3.7e-20 
C4507 VCC.n724 VSS 3.5e-20 
C4508 VCC.n725 VSS 5.76e-20 
C4509 VCC.n726 VSS 4.73e-20 
C4510 VCC.n727 VSS 3.09e-20 
C4511 VCC.n728 VSS 3.5e-20 
C4512 VCC.n729 VSS 3.5e-20 
C4513 VCC.n730 VSS 3.5e-20 
C4514 VCC.n731 VSS 1.18e-19 
C4515 VCC.n732 VSS 3e-20 
C4516 VCC.n733 VSS 1.15e-19 
C4517 VCC.n734 VSS 9.88e-20 
C4518 VCC.n735 VSS 5.76e-20 
C4519 VCC.n736 VSS 3.5e-20 
C4520 VCC.n737 VSS 3.09e-20 
C4521 VCC.n738 VSS 3.09e-20 
C4522 VCC.n739 VSS 2.26e-20 
C4523 VCC.n740 VSS 5.76e-20 
C4524 VCC.n741 VSS 2.68e-20 
C4525 VCC.n742 VSS 2.68e-20 
C4526 VCC.n743 VSS 0.00185f 
C4527 VCC.n744 VSS 2.72e-19 
C4528 VCC.n745 VSS 2.26e-20 
C4529 VCC.n746 VSS 1.87e-19 
C4530 VCC.n747 VSS 3.5e-20 
C4531 VCC.n748 VSS 2.68e-20 
C4532 VCC.n749 VSS 5.97e-20 
C4533 VCC.n750 VSS 4.73e-20 
C4534 VCC.n751 VSS 4.73e-20 
C4535 VCC.n752 VSS 5.15e-20 
C4536 VCC.n753 VSS 7.41e-20 
C4537 VCC.n754 VSS 3.7e-20 
C4538 VCC.n755 VSS 2.26e-20 
C4539 VCC.n756 VSS 6.38e-20 
C4540 VCC.n757 VSS 4.73e-20 
C4541 VCC.n758 VSS 3.29e-20 
C4542 VCC.n759 VSS 3.5e-20 
C4543 VCC.n760 VSS 3e-20 
C4544 VCC.t304 VSS 0.005f 
C4545 VCC.t146 VSS 0.00453f 
C4546 VCC.n761 VSS 0.00228f 
C4547 VCC.n762 VSS 1.3e-19 
C4548 VCC.t305 VSS 4.05e-19 
C4549 VCC.n763 VSS 4.05e-19 
C4550 VCC.n764 VSS 1.15e-19 
C4551 VCC.n765 VSS 3.36e-19 
C4552 VCC.n766 VSS 6.17e-21 
C4553 VCC.n767 VSS 3.12e-19 
C4554 VCC.n768 VSS 1.65e-20 
C4555 VCC.n769 VSS 1.54e-19 
C4556 VCC.n770 VSS 1.54e-19 
C4557 VCC.n771 VSS 1.65e-20 
C4558 VCC.n772 VSS 1.03e-20 
C4559 VCC.n773 VSS 3.5e-20 
C4560 VCC.n774 VSS 2.26e-20 
C4561 VCC.n775 VSS 4.73e-20 
C4562 VCC.n776 VSS 3.5e-20 
C4563 VCC.n777 VSS 3e-20 
C4564 VCC.n778 VSS 1.3e-19 
C4565 VCC.n779 VSS 5.12e-19 
C4566 VCC.n780 VSS 1.3e-19 
C4567 VCC.n781 VSS 4.13e-19 
C4568 VCC.n782 VSS 9.53e-20 
C4569 VCC.n783 VSS 5.76e-20 
C4570 VCC.n784 VSS 7.41e-20 
C4571 VCC.n785 VSS 5.56e-20 
C4572 VCC.t306 VSS 1.55e-19 
C4573 VCC.n786 VSS 3.91e-20 
C4574 VCC.n787 VSS 3.91e-20 
C4575 VCC.n788 VSS 1.85e-20 
C4576 VCC.n789 VSS 7.55e-19 
C4577 VCC.n790 VSS 4.94e-20 
C4578 VCC.n791 VSS 5.15e-20 
C4579 VCC.n792 VSS 7.2e-20 
C4580 VCC.n793 VSS 1.38e-19 
C4581 VCC.n794 VSS 1.17e-19 
C4582 VCC.n795 VSS 4.32e-20 
C4583 VCC.n796 VSS 2.88e-20 
C4584 VCC.n797 VSS 2.68e-20 
C4585 VCC.n798 VSS 3.5e-20 
C4586 VCC.n799 VSS 3.5e-20 
C4587 VCC.n800 VSS 2.88e-20 
C4588 VCC.n801 VSS 2.68e-20 
C4589 VCC.n802 VSS 2.68e-20 
C4590 VCC.n803 VSS 2.68e-20 
C4591 VCC.n804 VSS 4.12e-20 
C4592 VCC.n805 VSS 4.12e-20 
C4593 VCC.n806 VSS 3.91e-20 
C4594 VCC.n807 VSS 4.53e-20 
C4595 VCC.n808 VSS 4.53e-20 
C4596 VCC.n809 VSS 1.05e-19 
C4597 VCC.n810 VSS 1.05e-19 
C4598 VCC.n811 VSS 4.32e-20 
C4599 VCC.n812 VSS 3.7e-20 
C4600 VCC.n813 VSS 2.68e-20 
C4601 VCC.n814 VSS 2.68e-20 
C4602 VCC.n815 VSS 6.79e-20 
C4603 VCC.n816 VSS 9.26e-20 
C4604 VCC.n817 VSS 1.83e-19 
C4605 VCC.n818 VSS 7.95e-19 
C4606 VCC.n819 VSS 5.2e-19 
C4607 VCC.n820 VSS 1.3e-19 
C4608 VCC.n821 VSS 3e-20 
C4609 VCC.n822 VSS 3.5e-20 
C4610 VCC.n823 VSS 5.97e-20 
C4611 VCC.n824 VSS 7.41e-20 
C4612 VCC.n825 VSS 5.15e-20 
C4613 VCC.n826 VSS 5.15e-20 
C4614 VCC.n827 VSS 3.09e-20 
C4615 VCC.n828 VSS 3.09e-20 
C4616 VCC.n829 VSS 3.7e-20 
C4617 VCC.n830 VSS 2.68e-20 
C4618 VCC.n831 VSS 3.91e-20 
C4619 VCC.n832 VSS 1.17e-19 
C4620 VCC.n833 VSS 1.38e-19 
C4621 VCC.n834 VSS 7e-20 
C4622 VCC.n835 VSS 4.73e-20 
C4623 VCC.n836 VSS 3.5e-20 
C4624 VCC.n837 VSS 3.5e-20 
C4625 VCC.n838 VSS 3.5e-20 
C4626 VCC.n839 VSS 4.53e-20 
C4627 VCC.n840 VSS 1.18e-19 
C4628 VCC.n841 VSS 5.12e-19 
C4629 VCC.n842 VSS 1.3e-19 
C4630 VCC.n843 VSS 1.61e-19 
C4631 VCC.n844 VSS 9.9e-20 
C4632 VCC.n845 VSS 0.00243f 
C4633 VCC.n846 VSS 2.26e-20 
C4634 VCC.n847 VSS 4.13e-19 
C4635 VCC.n848 VSS 3.5e-20 
C4636 VCC.n849 VSS 3.5e-20 
C4637 VCC.n850 VSS 2.47e-20 
C4638 VCC.n851 VSS 2.06e-20 
C4639 VCC.n852 VSS 6.17e-20 
C4640 VCC.n853 VSS 6.17e-20 
C4641 VCC.n854 VSS 4.73e-20 
C4642 VCC.n855 VSS 4.73e-20 
C4643 VCC.n856 VSS 2.88e-20 
C4644 VCC.n857 VSS 1.44e-20 
C4645 VCC.n858 VSS 1.65e-20 
C4646 VCC.n859 VSS 1.54e-19 
C4647 VCC.n860 VSS 1.54e-19 
C4648 VCC.n861 VSS 1.65e-20 
C4649 VCC.n862 VSS 3.09e-20 
C4650 VCC.t236 VSS 1.55e-19 
C4651 VCC.n863 VSS 0.00102f 
C4652 VCC.n864 VSS 2.73e-19 
C4653 VCC.n865 VSS 0.00136f 
C4654 VCC.n866 VSS 2.73e-19 
C4655 VCC.n867 VSS 0.00181f 
C4656 VCC.n868 VSS 5.76e-20 
C4657 VCC.n869 VSS 1.54e-19 
C4658 VCC.n870 VSS 1.65e-20 
C4659 VCC.n871 VSS 2.88e-20 
C4660 VCC.n872 VSS 2.47e-20 
C4661 VCC.n873 VSS 6.17e-20 
C4662 VCC.n874 VSS 4.73e-20 
C4663 VCC.n875 VSS 4.73e-20 
C4664 VCC.n876 VSS 5.15e-20 
C4665 VCC.n877 VSS 3.5e-20 
C4666 VCC.n878 VSS 7.41e-20 
C4667 VCC.n879 VSS 3.7e-20 
C4668 VCC.n880 VSS 2.26e-20 
C4669 VCC.n881 VSS 6.17e-20 
C4670 VCC.n882 VSS 4.73e-20 
C4671 VCC.n883 VSS 3.5e-20 
C4672 VCC.n884 VSS 2.88e-20 
C4673 VCC.n885 VSS 3.4e-19 
C4674 VCC.n886 VSS 1.15e-19 
C4675 VCC.n887 VSS 3.98e-19 
C4676 VCC.t105 VSS 4.05e-19 
C4677 VCC.n888 VSS 1.22e-19 
C4678 VCC.n889 VSS 1.3e-19 
C4679 VCC.n890 VSS 3e-20 
C4680 VCC.n891 VSS 3.5e-20 
C4681 VCC.n892 VSS 3.5e-20 
C4682 VCC.n893 VSS 4.73e-20 
C4683 VCC.n894 VSS 2.47e-20 
C4684 VCC.n895 VSS 1.23e-20 
C4685 VCC.n896 VSS 1.65e-20 
C4686 VCC.n897 VSS 2.47e-20 
C4687 VCC.n898 VSS 5.76e-20 
C4688 VCC.n899 VSS 1.38e-19 
C4689 VCC.n900 VSS 7e-20 
C4690 VCC.n901 VSS 3.7e-20 
C4691 VCC.n902 VSS 2.47e-20 
C4692 VCC.n903 VSS 3.7e-20 
C4693 VCC.n904 VSS 1.85e-20 
C4694 VCC.n905 VSS 3.09e-20 
C4695 VCC.n906 VSS 5.35e-20 
C4696 VCC.n907 VSS 4.73e-20 
C4697 VCC.n908 VSS 5.35e-20 
C4698 VCC.n909 VSS 7.41e-20 
C4699 VCC.n910 VSS 5.76e-20 
C4700 VCC.n911 VSS 9.53e-20 
C4701 VCC.n912 VSS 4.13e-19 
C4702 VCC.n913 VSS 1.3e-19 
C4703 VCC.n914 VSS 5.2e-19 
C4704 VCC.n915 VSS 1.2e-19 
C4705 VCC.n916 VSS 4.73e-20 
C4706 VCC.n917 VSS 2.68e-20 
C4707 VCC.n918 VSS 3.5e-20 
C4708 VCC.n919 VSS 3.5e-20 
C4709 VCC.n920 VSS 2.68e-20 
C4710 VCC.n921 VSS 2.68e-20 
C4711 VCC.n922 VSS 4.32e-20 
C4712 VCC.n923 VSS 4.32e-20 
C4713 VCC.n924 VSS 4.32e-20 
C4714 VCC.n925 VSS 2.88e-20 
C4715 VCC.n926 VSS 3.5e-20 
C4716 VCC.n927 VSS 2.68e-20 
C4717 VCC.n928 VSS 7.82e-20 
C4718 VCC.n929 VSS 4.73e-20 
C4719 VCC.n930 VSS 4.73e-20 
C4720 VCC.n931 VSS 1.05e-19 
C4721 VCC.n932 VSS 1.05e-19 
C4722 VCC.n933 VSS 4.53e-20 
C4723 VCC.n934 VSS 2.68e-20 
C4724 VCC.n935 VSS 2.68e-20 
C4725 VCC.n936 VSS 6.59e-20 
C4726 VCC.n937 VSS 9.26e-20 
C4727 VCC.n938 VSS 6.59e-20 
C4728 VCC.n939 VSS 2.47e-20 
C4729 VCC.n940 VSS 2.47e-20 
C4730 VCC.n941 VSS 2.88e-20 
C4731 VCC.n942 VSS 3.5e-20 
C4732 VCC.n943 VSS 3.5e-20 
C4733 VCC.n944 VSS 4.53e-20 
C4734 VCC.n945 VSS 1.2e-19 
C4735 VCC.n946 VSS 5.2e-19 
C4736 VCC.n947 VSS 1.3e-19 
C4737 VCC.n948 VSS 4.13e-19 
C4738 VCC.n949 VSS 9.53e-20 
C4739 VCC.n950 VSS 5.97e-20 
C4740 VCC.n951 VSS 7.41e-20 
C4741 VCC.n952 VSS 5.35e-20 
C4742 VCC.n953 VSS 5.15e-20 
C4743 VCC.n954 VSS 3.09e-20 
C4744 VCC.n955 VSS 3.09e-20 
C4745 VCC.n956 VSS 3.91e-20 
C4746 VCC.n957 VSS 2.47e-20 
C4747 VCC.n958 VSS 3.7e-20 
C4748 VCC.n959 VSS 1.17e-19 
C4749 VCC.n960 VSS 1.38e-19 
C4750 VCC.n961 VSS 7.2e-20 
C4751 VCC.n962 VSS 4.73e-20 
C4752 VCC.n963 VSS 3.5e-20 
C4753 VCC.n964 VSS 3.5e-20 
C4754 VCC.n965 VSS 4.53e-20 
C4755 VCC.n966 VSS 5.97e-20 
C4756 VCC.n967 VSS 3.5e-20 
C4757 VCC.n968 VSS 3e-20 
C4758 VCC.n969 VSS 1.3e-19 
C4759 VCC.n970 VSS 1.53e-19 
C4760 VCC.t212 VSS 4.05e-19 
C4761 VCC.n971 VSS 2.06e-19 
C4762 VCC.n972 VSS 1.35e-19 
C4763 VCC.n973 VSS 9.67e-20 
C4764 VCC.n974 VSS 3.35e-20 
C4765 VCC.n975 VSS 3.5e-20 
C4766 VCC.n976 VSS 2.36e-19 
C4767 VCC.n977 VSS 0.0023f 
C4768 VCC.t28 VSS 0.0031f 
C4769 VCC.t133 VSS 0.00366f 
C4770 VCC.t31 VSS 0.00365f 
C4771 VCC.t136 VSS 0.00386f 
C4772 VCC.n978 VSS 0.00569f 
C4773 VCC.n979 VSS 1.3e-19 
C4774 VCC.n980 VSS 3.67e-19 
C4775 VCC.n981 VSS 1.15e-19 
C4776 VCC.n982 VSS 3.38e-19 
C4777 VCC.n983 VSS 3.5e-20 
C4778 VCC.n984 VSS 3.5e-20 
C4779 VCC.n985 VSS 2.68e-20 
C4780 VCC.n986 VSS 2.06e-20 
C4781 VCC.n987 VSS 6.38e-20 
C4782 VCC.n988 VSS 5.97e-20 
C4783 VCC.n989 VSS 4.73e-20 
C4784 VCC.n990 VSS 4.73e-20 
C4785 VCC.n991 VSS 3.09e-20 
C4786 VCC.n992 VSS 1.23e-20 
C4787 VCC.n993 VSS 1.65e-20 
C4788 VCC.n994 VSS 1.54e-19 
C4789 VCC.n995 VSS 1.54e-19 
C4790 VCC.n996 VSS 1.65e-20 
C4791 VCC.n997 VSS 3.29e-20 
C4792 VCC.t213 VSS 1.67e-19 
C4793 VCC.n998 VSS 0.00101f 
C4794 VCC.n999 VSS 2.71e-19 
C4795 VCC.n1000 VSS 7.46e-19 
C4796 VCC.n1001 VSS 0.00333f 
C4797 VCC.n1002 VSS 2.46e-19 
C4798 VCC.n1003 VSS 3.02e-19 
C4799 VCC.n1004 VSS 3.7e-20 
C4800 VCC.n1005 VSS 5.15e-20 
C4801 VCC.n1006 VSS 6.38e-20 
C4802 VCC.n1007 VSS 4.73e-20 
C4803 VCC.n1008 VSS 4.73e-20 
C4804 VCC.n1009 VSS 2.68e-20 
C4805 VCC.n1010 VSS 3.29e-20 
C4806 VCC.n1011 VSS 1.65e-20 
C4807 VCC.n1012 VSS 1.54e-19 
C4808 VCC.n1013 VSS 1.54e-19 
C4809 VCC.n1014 VSS 5.56e-20 
C4810 VCC.n1015 VSS 2.88e-20 
C4811 VCC.n1016 VSS 1.65e-20 
C4812 VCC.n1017 VSS 3.09e-20 
C4813 VCC.n1018 VSS 4.73e-20 
C4814 VCC.n1019 VSS 4.73e-20 
C4815 VCC.n1020 VSS 4.32e-20 
C4816 VCC.n1021 VSS 1.17e-19 
C4817 VCC.n1022 VSS 3.33e-19 
C4818 VCC.n1023 VSS 1.35e-19 
C4819 VCC.n1024 VSS 4.37e-19 
C4820 VCC.n1025 VSS 5.24e-19 
C4821 VCC.n1026 VSS 1.36e-19 
C4822 VCC.n1027 VSS 1.01e-19 
C4823 VCC.n1028 VSS 1.05e-19 
C4824 VCC.n1029 VSS 2.06e-20 
C4825 VCC.n1030 VSS 2.26e-20 
C4826 VCC.n1031 VSS 3.7e-20 
C4827 VCC.n1032 VSS 5.15e-20 
C4828 VCC.n1033 VSS 1.38e-19 
C4829 VCC.n1034 VSS 3.91e-20 
C4830 VCC.n1035 VSS 2.88e-20 
C4831 VCC.n1036 VSS 4.32e-20 
C4832 VCC.n1037 VSS 1.17e-19 
C4833 VCC.n1038 VSS 3.7e-20 
C4834 VCC.n1039 VSS 3.91e-20 
C4835 VCC.n1040 VSS 3.5e-20 
C4836 VCC.n1041 VSS 1.65e-20 
C4837 VCC.n1042 VSS 8.23e-21 
C4838 VCC.n1043 VSS 3.5e-20 
C4839 VCC.n1044 VSS 3.5e-20 
C4840 VCC.n1045 VSS 1.4e-19 
C4841 VCC.n1046 VSS 5.4e-19 
C4842 VCC.n1047 VSS 8.42e-19 
C4843 VCC.n1048 VSS 5.4e-19 
C4844 VCC.n1049 VSS 1.4e-19 
C4845 VCC.n1050 VSS 1.4e-19 
C4846 VCC.n1051 VSS 2.18e-19 
C4847 VCC.n1052 VSS 7.82e-20 
C4848 VCC.n1053 VSS 4.32e-20 
C4849 VCC.n1054 VSS 4.32e-20 
C4850 VCC.n1055 VSS 1.05e-19 
C4851 VCC.n1056 VSS 1.05e-19 
C4852 VCC.n1057 VSS 4.32e-20 
C4853 VCC.n1058 VSS 3.7e-20 
C4854 VCC.n1059 VSS 2.68e-20 
C4855 VCC.n1060 VSS 5.76e-20 
C4856 VCC.n1061 VSS 6.38e-20 
C4857 VCC.n1062 VSS 3.5e-20 
C4858 VCC.n1063 VSS 3.5e-20 
C4859 VCC.n1064 VSS 1.17e-19 
C4860 VCC.n1065 VSS 1.38e-19 
C4861 VCC.n1066 VSS 5.15e-20 
C4862 VCC.n1067 VSS 1.05e-19 
C4863 VCC.n1068 VSS 2.26e-20 
C4864 VCC.n1069 VSS 5.76e-20 
C4865 VCC.n1070 VSS 3.7e-20 
C4866 VCC.n1071 VSS 3.7e-20 
C4867 VCC.n1072 VSS 3.09e-20 
C4868 VCC.n1073 VSS 1.85e-20 
C4869 VCC.n1074 VSS 1.65e-20 
C4870 VCC.n1075 VSS 8.23e-21 
C4871 VCC.n1076 VSS 1.13e-19 
C4872 VCC.n1077 VSS 3.33e-19 
C4873 VCC.t284 VSS 4.21e-19 
C4874 VCC.n1078 VSS 2.06e-19 
C4875 VCC.n1079 VSS 1.35e-19 
C4876 VCC.n1080 VSS 3.5e-20 
C4877 VCC.n1081 VSS 3.5e-20 
C4878 VCC.n1082 VSS 3.5e-20 
C4879 VCC.n1083 VSS 1.03e-20 
C4880 VCC.n1084 VSS 2.68e-20 
C4881 VCC.n1085 VSS 3.09e-20 
C4882 VCC.n1086 VSS 2.68e-20 
C4883 VCC.n1087 VSS 1.65e-20 
C4884 VCC.n1088 VSS 1.54e-19 
C4885 VCC.n1089 VSS 1.54e-19 
C4886 VCC.n1090 VSS 1.65e-20 
C4887 VCC.t285 VSS 1.56e-19 
C4888 VCC.n1091 VSS 7.62e-19 
C4889 VCC.n1092 VSS 1.23e-20 
C4890 VCC.n1093 VSS 2.47e-20 
C4891 VCC.n1094 VSS 4.73e-20 
C4892 VCC.n1095 VSS 6.59e-20 
C4893 VCC.n1096 VSS 5.15e-20 
C4894 VCC.n1097 VSS 2.47e-20 
C4895 VCC.n1098 VSS 7.41e-20 
C4896 VCC.n1099 VSS 9.47e-20 
C4897 VCC.n1100 VSS 1.32e-19 
C4898 VCC.n1101 VSS 7.71e-19 
C4899 VCC.n1102 VSS 9.83e-19 
C4900 VCC.n1103 VSS 2.36e-19 
C4901 VCC.n1104 VSS 3.21e-19 
C4902 VCC.n1105 VSS 2.61e-19 
C4903 VCC.n1106 VSS 0.00189f 
C4904 VCC.n1107 VSS 0.00274f 
C4905 VCC.n1108 VSS 5.76e-20 
C4906 VCC.n1109 VSS 2.88e-20 
C4907 VCC.n1110 VSS 3.5e-20 
C4908 VCC.n1111 VSS 9.83e-19 
C4909 VCC.n1112 VSS 9.47e-20 
C4910 VCC.n1113 VSS 1.17e-19 
C4911 VCC.n1114 VSS 2.06e-19 
C4912 VCC.n1115 VSS 1.36e-19 
C4913 VCC.n1116 VSS 1.01e-19 
C4914 VCC.n1117 VSS 3.5e-20 
C4915 VCC.n1118 VSS 3.09e-20 
C4916 VCC.n1119 VSS 3.29e-20 
C4917 VCC.n1120 VSS 3.29e-20 
C4918 VCC.n1121 VSS 4.73e-20 
C4919 VCC.n1122 VSS 1.44e-20 
C4920 VCC.n1123 VSS 3.5e-20 
C4921 VCC.n1124 VSS 7.41e-20 
C4922 VCC.n1125 VSS 2.47e-20 
C4923 VCC.t135 VSS 1.56e-19 
C4924 VCC.n1126 VSS 5.76e-20 
C4925 VCC.n1127 VSS 2.06e-20 
C4926 VCC.n1128 VSS 5.76e-20 
C4927 VCC.n1129 VSS 3.7e-20 
C4928 VCC.n1130 VSS 4.32e-20 
C4929 VCC.n1131 VSS 2.68e-20 
C4930 VCC.n1132 VSS 3.91e-20 
C4931 VCC.n1133 VSS 6.38e-20 
C4932 VCC.n1134 VSS 1.85e-20 
C4933 VCC.n1135 VSS 3.5e-20 
C4934 VCC.n1136 VSS 3.09e-20 
C4935 VCC.n1137 VSS 3.7e-20 
C4936 VCC.n1138 VSS 3.09e-20 
C4937 VCC.n1139 VSS 2.26e-20 
C4938 VCC.n1140 VSS 1.05e-19 
C4939 VCC.n1141 VSS 3.5e-20 
C4940 VCC.n1142 VSS 3.5e-20 
C4941 VCC.n1143 VSS 8.42e-19 
C4942 VCC.n1144 VSS 2.18e-19 
C4943 VCC.n1145 VSS 1.4e-19 
C4944 VCC.n1146 VSS 4.32e-20 
C4945 VCC.n1147 VSS 7.82e-20 
C4946 VCC.n1148 VSS 5.76e-20 
C4947 VCC.n1149 VSS 2.68e-20 
C4948 VCC.n1150 VSS 4.32e-20 
C4949 VCC.n1151 VSS 3.91e-20 
C4950 VCC.n1152 VSS 3.7e-20 
C4951 VCC.n1153 VSS 3.7e-20 
C4952 VCC.n1154 VSS 5.76e-20 
C4953 VCC.n1155 VSS 4.73e-20 
C4954 VCC.n1156 VSS 3.5e-20 
C4955 VCC.t25 VSS 1.56e-19 
C4956 VCC.n1157 VSS 7.97e-19 
C4957 VCC.n1158 VSS 3.09e-20 
C4958 VCC.n1159 VSS 1.01e-19 
C4959 VCC.n1160 VSS 3.5e-20 
C4960 VCC.n1161 VSS 1.36e-19 
C4961 VCC.n1162 VSS 3.5e-20 
C4962 VCC.n1163 VSS 3.33e-19 
C4963 VCC.n1164 VSS 1.17e-19 
C4964 VCC.n1165 VSS 1.09e-19 
C4965 VCC.n1166 VSS 3.5e-20 
C4966 VCC.n1167 VSS 4.73e-20 
C4967 VCC.n1168 VSS 5.56e-20 
C4968 VCC.n1169 VSS 2.88e-20 
C4969 VCC.n1170 VSS 2.26e-20 
C4970 VCC.n1171 VSS 5.76e-20 
C4971 VCC.n1172 VSS 2.68e-20 
C4972 VCC.n1173 VSS 2.68e-20 
C4973 VCC.n1174 VSS 1.9e-19 
C4974 VCC.n1175 VSS 5.76e-20 
C4975 VCC.n1176 VSS 2.68e-20 
C4976 VCC.n1177 VSS 2.68e-20 
C4977 VCC.n1178 VSS 2.68e-20 
C4978 VCC.n1179 VSS 5.76e-20 
C4979 VCC.n1180 VSS 2.26e-20 
C4980 VCC.n1181 VSS 3.09e-20 
C4981 VCC.n1182 VSS 2.26e-20 
C4982 VCC.n1183 VSS 5.15e-20 
C4983 VCC.n1184 VSS 4.73e-20 
C4984 VCC.n1185 VSS 3.7e-20 
C4985 VCC.n1186 VSS 3.5e-20 
C4986 VCC.n1187 VSS 7.41e-20 
C4987 VCC.n1188 VSS 1.91e-19 
C4988 VCC.n1189 VSS 9.88e-20 
C4989 VCC.n1190 VSS 3e-20 
C4990 VCC.n1191 VSS 5.12e-19 
C4991 VCC.n1192 VSS 1.18e-19 
C4992 VCC.n1193 VSS 3.5e-20 
C4993 VCC.n1194 VSS 3.5e-20 
C4994 VCC.n1195 VSS 5.15e-20 
C4995 VCC.n1196 VSS 4.32e-20 
C4996 VCC.n1197 VSS 2.68e-20 
C4997 VCC.n1198 VSS 3.91e-20 
C4998 VCC.n1199 VSS 1.44e-20 
C4999 VCC.n1200 VSS 3.5e-20 
C5000 VCC.n1201 VSS 3e-20 
C5001 VCC.n1202 VSS 7.95e-19 
C5002 VCC.n1203 VSS 1.83e-19 
C5003 VCC.n1204 VSS 2.88e-20 
C5004 VCC.n1205 VSS 2.68e-20 
C5005 VCC.n1206 VSS 2.68e-20 
C5006 VCC.n1207 VSS 2.68e-20 
C5007 VCC.n1208 VSS 4.53e-20 
C5008 VCC.n1209 VSS 3.7e-20 
C5009 VCC.n1210 VSS 7.82e-20 
C5010 VCC.n1211 VSS 1.17e-19 
C5011 VCC.n1212 VSS 3.91e-20 
C5012 VCC.n1213 VSS 1.65e-20 
C5013 VCC.n1214 VSS 2.68e-20 
C5014 VCC.n1215 VSS 3.5e-20 
C5015 VCC.n1216 VSS 3e-20 
C5016 VCC.n1217 VSS 5.12e-19 
C5017 VCC.n1218 VSS 1.18e-19 
C5018 VCC.n1219 VSS 3.5e-20 
C5019 VCC.n1220 VSS 3.5e-20 
C5020 VCC.t139 VSS 1.55e-19 
C5021 VCC.n1221 VSS 7.57e-19 
C5022 VCC.n1222 VSS 4.73e-20 
C5023 VCC.n1223 VSS 1.54e-19 
C5024 VCC.n1224 VSS 2.88e-20 
C5025 VCC.n1225 VSS 2.88e-20 
C5026 VCC.n1226 VSS 3.5e-20 
C5027 VCC.n1227 VSS 5.76e-20 
C5028 VCC.n1228 VSS 9.88e-20 
C5029 VCC.n1229 VSS 1.3e-19 
C5030 VCC.n1230 VSS 3e-20 
C5031 VCC.t137 VSS 0.005f 
C5032 VCC.t17 VSS 0.00453f 
C5033 VCC.n1231 VSS 0.00229f 
C5034 VCC.n1232 VSS 1.91e-19 
C5035 VCC.n1233 VSS 3.5e-20 
C5036 VCC.n1234 VSS 3.14e-19 
C5037 VCC.n1235 VSS 3.5e-20 
C5038 VCC.n1236 VSS 2.47e-20 
C5039 VCC.n1237 VSS 5.76e-20 
C5040 VCC.n1238 VSS 2.47e-20 
C5041 VCC.n1239 VSS 8.23e-21 
C5042 VCC.n1240 VSS 2.88e-20 
C5043 VCC.n1241 VSS 5.76e-20 
C5044 VCC.n1242 VSS 2.47e-20 
C5045 VCC.n1243 VSS 2.88e-20 
C5046 VCC.n1244 VSS 2.47e-20 
C5047 VCC.n1245 VSS 5.15e-20 
C5048 VCC.n1246 VSS 4.73e-20 
C5049 VCC.n1247 VSS 3.7e-20 
C5050 VCC.n1248 VSS 3.5e-20 
C5051 VCC.n1249 VSS 7.41e-20 
C5052 VCC.t149 VSS 6.42e-19 
C5053 VCC.n1250 VSS 3e-20 
C5054 VCC.n1251 VSS 5.97e-20 
C5055 VCC.n1252 VSS 4.13e-19 
C5056 VCC.n1253 VSS 9.53e-20 
C5057 VCC.n1254 VSS 3.5e-20 
C5058 VCC.n1255 VSS 3.5e-20 
C5059 VCC.n1256 VSS 5.35e-20 
C5060 VCC.n1257 VSS 4.32e-20 
C5061 VCC.n1258 VSS 2.68e-20 
C5062 VCC.n1259 VSS 3.7e-20 
C5063 VCC.n1260 VSS 1.65e-20 
C5064 VCC.n1261 VSS 4.53e-20 
C5065 VCC.n1262 VSS 1.2e-19 
C5066 VCC.n1263 VSS 5.2e-19 
C5067 VCC.n1264 VSS 1.2e-19 
C5068 VCC.n1265 VSS 6.38e-20 
C5069 VCC.n1266 VSS 2.47e-20 
C5070 VCC.n1267 VSS 4.53e-20 
C5071 VCC.n1268 VSS 3.5e-20 
C5072 VCC.n1269 VSS 3.5e-20 
C5073 VCC.n1270 VSS 2.68e-20 
C5074 VCC.n1271 VSS 2.68e-20 
C5075 VCC.n1272 VSS 2.47e-20 
C5076 VCC.n1273 VSS 4.53e-20 
C5077 VCC.n1274 VSS 2.68e-20 
C5078 VCC.n1275 VSS 4.32e-20 
C5079 VCC.n1276 VSS 2.68e-20 
C5080 VCC.n1277 VSS 3.91e-20 
C5081 VCC.n1278 VSS 2.88e-20 
C5082 VCC.n1279 VSS 4.73e-20 
C5083 VCC.n1280 VSS 3.7e-20 
C5084 VCC.n1281 VSS 3.7e-20 
C5085 VCC.n1282 VSS 3.5e-20 
C5086 VCC.n1283 VSS 5.76e-20 
C5087 VCC.n1284 VSS 4.73e-20 
C5088 VCC.n1285 VSS 3.09e-20 
C5089 VCC.n1286 VSS 3.5e-20 
C5090 VCC.n1287 VSS 3.5e-20 
C5091 VCC.n1288 VSS 3.5e-20 
C5092 VCC.n1289 VSS 1.18e-19 
C5093 VCC.n1290 VSS 3e-20 
C5094 VCC.n1291 VSS 1.15e-19 
C5095 VCC.n1292 VSS 9.88e-20 
C5096 VCC.n1293 VSS 5.76e-20 
C5097 VCC.n1294 VSS 3.5e-20 
C5098 VCC.n1295 VSS 3.09e-20 
C5099 VCC.n1296 VSS 3.09e-20 
C5100 VCC.n1297 VSS 2.26e-20 
C5101 VCC.n1298 VSS 5.76e-20 
C5102 VCC.n1299 VSS 2.68e-20 
C5103 VCC.n1300 VSS 2.68e-20 
C5104 VCC.n1301 VSS 0.00185f 
C5105 VCC.n1302 VSS 2.72e-19 
C5106 VCC.n1303 VSS 2.26e-20 
C5107 VCC.n1304 VSS 1.87e-19 
C5108 VCC.n1305 VSS 3.5e-20 
C5109 VCC.n1306 VSS 2.68e-20 
C5110 VCC.n1307 VSS 5.97e-20 
C5111 VCC.n1308 VSS 4.73e-20 
C5112 VCC.n1309 VSS 4.73e-20 
C5113 VCC.n1310 VSS 5.15e-20 
C5114 VCC.n1311 VSS 7.41e-20 
C5115 VCC.n1312 VSS 3.7e-20 
C5116 VCC.n1313 VSS 2.26e-20 
C5117 VCC.n1314 VSS 6.38e-20 
C5118 VCC.n1315 VSS 4.73e-20 
C5119 VCC.n1316 VSS 3.29e-20 
C5120 VCC.n1317 VSS 3.5e-20 
C5121 VCC.n1318 VSS 3e-20 
C5122 VCC.t6 VSS 0.005f 
C5123 VCC.t34 VSS 0.00453f 
C5124 VCC.n1319 VSS 0.00228f 
C5125 VCC.n1320 VSS 1.3e-19 
C5126 VCC.t4 VSS 4.05e-19 
C5127 VCC.n1321 VSS 4.05e-19 
C5128 VCC.n1322 VSS 1.15e-19 
C5129 VCC.n1323 VSS 3.36e-19 
C5130 VCC.n1324 VSS 6.17e-21 
C5131 VCC.n1325 VSS 3.12e-19 
C5132 VCC.n1326 VSS 1.65e-20 
C5133 VCC.n1327 VSS 1.54e-19 
C5134 VCC.n1328 VSS 1.54e-19 
C5135 VCC.n1329 VSS 1.65e-20 
C5136 VCC.n1330 VSS 1.03e-20 
C5137 VCC.n1331 VSS 3.5e-20 
C5138 VCC.n1332 VSS 2.26e-20 
C5139 VCC.n1333 VSS 4.73e-20 
C5140 VCC.n1334 VSS 3.5e-20 
C5141 VCC.n1335 VSS 3e-20 
C5142 VCC.n1336 VSS 1.3e-19 
C5143 VCC.n1337 VSS 5.12e-19 
C5144 VCC.n1338 VSS 1.3e-19 
C5145 VCC.n1339 VSS 4.13e-19 
C5146 VCC.n1340 VSS 9.53e-20 
C5147 VCC.n1341 VSS 5.76e-20 
C5148 VCC.n1342 VSS 7.41e-20 
C5149 VCC.n1343 VSS 5.56e-20 
C5150 VCC.t5 VSS 1.55e-19 
C5151 VCC.n1344 VSS 3.91e-20 
C5152 VCC.n1345 VSS 3.91e-20 
C5153 VCC.n1346 VSS 1.85e-20 
C5154 VCC.n1347 VSS 7.55e-19 
C5155 VCC.n1348 VSS 4.94e-20 
C5156 VCC.n1349 VSS 5.15e-20 
C5157 VCC.n1350 VSS 7.2e-20 
C5158 VCC.n1351 VSS 1.38e-19 
C5159 VCC.n1352 VSS 1.17e-19 
C5160 VCC.n1353 VSS 4.32e-20 
C5161 VCC.n1354 VSS 2.88e-20 
C5162 VCC.n1355 VSS 2.68e-20 
C5163 VCC.n1356 VSS 3.5e-20 
C5164 VCC.n1357 VSS 3.5e-20 
C5165 VCC.n1358 VSS 2.88e-20 
C5166 VCC.n1359 VSS 2.68e-20 
C5167 VCC.n1360 VSS 2.68e-20 
C5168 VCC.n1361 VSS 2.68e-20 
C5169 VCC.n1362 VSS 4.12e-20 
C5170 VCC.n1363 VSS 4.12e-20 
C5171 VCC.n1364 VSS 3.91e-20 
C5172 VCC.n1365 VSS 4.53e-20 
C5173 VCC.n1366 VSS 4.53e-20 
C5174 VCC.n1367 VSS 1.05e-19 
C5175 VCC.n1368 VSS 1.05e-19 
C5176 VCC.n1369 VSS 4.32e-20 
C5177 VCC.n1370 VSS 3.7e-20 
C5178 VCC.n1371 VSS 2.68e-20 
C5179 VCC.n1372 VSS 2.68e-20 
C5180 VCC.n1373 VSS 6.79e-20 
C5181 VCC.n1374 VSS 9.26e-20 
C5182 VCC.n1375 VSS 1.83e-19 
C5183 VCC.n1376 VSS 7.95e-19 
C5184 VCC.n1377 VSS 5.2e-19 
C5185 VCC.n1378 VSS 1.3e-19 
C5186 VCC.n1379 VSS 3e-20 
C5187 VCC.n1380 VSS 3.5e-20 
C5188 VCC.n1381 VSS 5.97e-20 
C5189 VCC.n1382 VSS 7.41e-20 
C5190 VCC.n1383 VSS 5.15e-20 
C5191 VCC.n1384 VSS 5.15e-20 
C5192 VCC.n1385 VSS 3.09e-20 
C5193 VCC.n1386 VSS 3.09e-20 
C5194 VCC.n1387 VSS 3.7e-20 
C5195 VCC.n1388 VSS 2.68e-20 
C5196 VCC.n1389 VSS 3.91e-20 
C5197 VCC.n1390 VSS 1.17e-19 
C5198 VCC.n1391 VSS 1.38e-19 
C5199 VCC.n1392 VSS 7e-20 
C5200 VCC.n1393 VSS 4.73e-20 
C5201 VCC.n1394 VSS 3.5e-20 
C5202 VCC.n1395 VSS 3.5e-20 
C5203 VCC.n1396 VSS 3.5e-20 
C5204 VCC.n1397 VSS 4.53e-20 
C5205 VCC.n1398 VSS 1.18e-19 
C5206 VCC.n1399 VSS 5.12e-19 
C5207 VCC.n1400 VSS 1.3e-19 
C5208 VCC.n1401 VSS 1.61e-19 
C5209 VCC.n1402 VSS 9.9e-20 
C5210 VCC.n1403 VSS 0.00243f 
C5211 VCC.n1404 VSS 2.26e-20 
C5212 VCC.n1405 VSS 4.13e-19 
C5213 VCC.n1406 VSS 3.5e-20 
C5214 VCC.n1407 VSS 3.5e-20 
C5215 VCC.n1408 VSS 2.47e-20 
C5216 VCC.n1409 VSS 2.06e-20 
C5217 VCC.n1410 VSS 6.17e-20 
C5218 VCC.n1411 VSS 6.17e-20 
C5219 VCC.n1412 VSS 4.73e-20 
C5220 VCC.n1413 VSS 4.73e-20 
C5221 VCC.n1414 VSS 2.88e-20 
C5222 VCC.n1415 VSS 1.44e-20 
C5223 VCC.n1416 VSS 1.65e-20 
C5224 VCC.n1417 VSS 1.54e-19 
C5225 VCC.n1418 VSS 1.54e-19 
C5226 VCC.n1419 VSS 1.65e-20 
C5227 VCC.n1420 VSS 3.09e-20 
C5228 VCC.t150 VSS 1.55e-19 
C5229 VCC.n1421 VSS 0.00102f 
C5230 VCC.n1422 VSS 2.73e-19 
C5231 VCC.n1423 VSS 0.00136f 
C5232 VCC.n1424 VSS 2.73e-19 
C5233 VCC.n1425 VSS 0.00181f 
C5234 VCC.n1426 VSS 5.76e-20 
C5235 VCC.n1427 VSS 1.54e-19 
C5236 VCC.n1428 VSS 1.65e-20 
C5237 VCC.n1429 VSS 6.17e-20 
C5238 VCC.n1430 VSS 2.47e-20 
C5239 VCC.n1431 VSS 4.73e-20 
C5240 VCC.n1432 VSS 4.73e-20 
C5241 VCC.n1433 VSS 5.15e-20 
C5242 VCC.n1434 VSS 3.5e-20 
C5243 VCC.n1435 VSS 7.41e-20 
C5244 VCC.n1436 VSS 3.7e-20 
C5245 VCC.n1437 VSS 2.26e-20 
C5246 VCC.n1438 VSS 6.17e-20 
C5247 VCC.n1439 VSS 4.73e-20 
C5248 VCC.n1440 VSS 2.88e-20 
C5249 VCC.n1441 VSS 2.88e-20 
C5250 VCC.n1442 VSS 3.4e-19 
C5251 VCC.n1443 VSS 1.15e-19 
C5252 VCC.n1444 VSS 3.98e-19 
C5253 VCC.t138 VSS 4.05e-19 
C5254 VCC.n1445 VSS 1.22e-19 
C5255 VCC.n1446 VSS 1.3e-19 
C5256 VCC.n1447 VSS 3e-20 
C5257 VCC.n1448 VSS 3.5e-20 
C5258 VCC.n1449 VSS 3.5e-20 
C5259 VCC.n1450 VSS 4.73e-20 
C5260 VCC.n1451 VSS 2.47e-20 
C5261 VCC.n1452 VSS 1.23e-20 
C5262 VCC.n1453 VSS 1.65e-20 
C5263 VCC.n1454 VSS 2.47e-20 
C5264 VCC.n1455 VSS 5.76e-20 
C5265 VCC.n1456 VSS 1.38e-19 
C5266 VCC.n1457 VSS 7e-20 
C5267 VCC.n1458 VSS 3.7e-20 
C5268 VCC.n1459 VSS 2.47e-20 
C5269 VCC.n1460 VSS 3.7e-20 
C5270 VCC.n1461 VSS 1.85e-20 
C5271 VCC.n1462 VSS 3.09e-20 
C5272 VCC.n1463 VSS 5.35e-20 
C5273 VCC.n1464 VSS 4.73e-20 
C5274 VCC.n1465 VSS 5.35e-20 
C5275 VCC.n1466 VSS 7.41e-20 
C5276 VCC.n1467 VSS 5.76e-20 
C5277 VCC.n1468 VSS 9.53e-20 
C5278 VCC.n1469 VSS 4.13e-19 
C5279 VCC.n1470 VSS 1.3e-19 
C5280 VCC.n1471 VSS 5.2e-19 
C5281 VCC.n1472 VSS 1.2e-19 
C5282 VCC.n1473 VSS 4.73e-20 
C5283 VCC.n1474 VSS 2.68e-20 
C5284 VCC.n1475 VSS 3.5e-20 
C5285 VCC.n1476 VSS 3.5e-20 
C5286 VCC.n1477 VSS 2.68e-20 
C5287 VCC.n1478 VSS 2.68e-20 
C5288 VCC.n1479 VSS 4.32e-20 
C5289 VCC.n1480 VSS 4.32e-20 
C5290 VCC.n1481 VSS 4.32e-20 
C5291 VCC.n1482 VSS 2.88e-20 
C5292 VCC.n1483 VSS 3.5e-20 
C5293 VCC.n1484 VSS 2.68e-20 
C5294 VCC.n1485 VSS 7.82e-20 
C5295 VCC.n1486 VSS 4.73e-20 
C5296 VCC.n1487 VSS 4.73e-20 
C5297 VCC.n1488 VSS 1.05e-19 
C5298 VCC.n1489 VSS 1.05e-19 
C5299 VCC.n1490 VSS 4.53e-20 
C5300 VCC.n1491 VSS 2.68e-20 
C5301 VCC.n1492 VSS 2.68e-20 
C5302 VCC.n1493 VSS 6.59e-20 
C5303 VCC.n1494 VSS 9.26e-20 
C5304 VCC.n1495 VSS 6.59e-20 
C5305 VCC.n1496 VSS 2.47e-20 
C5306 VCC.n1497 VSS 2.47e-20 
C5307 VCC.n1498 VSS 2.88e-20 
C5308 VCC.n1499 VSS 3.5e-20 
C5309 VCC.n1500 VSS 3.5e-20 
C5310 VCC.n1501 VSS 4.53e-20 
C5311 VCC.n1502 VSS 1.2e-19 
C5312 VCC.n1503 VSS 5.2e-19 
C5313 VCC.n1504 VSS 1.3e-19 
C5314 VCC.n1505 VSS 4.13e-19 
C5315 VCC.n1506 VSS 9.53e-20 
C5316 VCC.n1507 VSS 5.97e-20 
C5317 VCC.n1508 VSS 7.41e-20 
C5318 VCC.n1509 VSS 5.35e-20 
C5319 VCC.n1510 VSS 5.15e-20 
C5320 VCC.n1511 VSS 3.09e-20 
C5321 VCC.n1512 VSS 3.09e-20 
C5322 VCC.n1513 VSS 3.91e-20 
C5323 VCC.n1514 VSS 2.47e-20 
C5324 VCC.n1515 VSS 3.7e-20 
C5325 VCC.n1516 VSS 1.17e-19 
C5326 VCC.n1517 VSS 1.38e-19 
C5327 VCC.n1518 VSS 7.2e-20 
C5328 VCC.n1519 VSS 4.73e-20 
C5329 VCC.n1520 VSS 3.5e-20 
C5330 VCC.n1521 VSS 3.5e-20 
C5331 VCC.n1522 VSS 4.53e-20 
C5332 VCC.n1523 VSS 5.97e-20 
C5333 VCC.n1524 VSS 3.5e-20 
C5334 VCC.n1525 VSS 3e-20 
C5335 VCC.n1526 VSS 1.3e-19 
C5336 VCC.n1527 VSS 1.53e-19 
C5337 VCC.t255 VSS 4.05e-19 
C5338 VCC.n1528 VSS 1.35e-19 
C5339 VCC.t24 VSS 4.21e-19 
C5340 VCC.n1529 VSS 2.06e-19 
C5341 VCC.n1530 VSS 1.32e-19 
C5342 VCC.n1531 VSS 9.67e-20 
C5343 VCC.n1532 VSS 3.35e-20 
C5344 VCC.n1533 VSS 3.5e-20 
C5345 VCC.n1534 VSS 2.36e-19 
C5346 VCC.n1535 VSS 0.0023f 
C5347 VCC.t27 VSS 0.0031f 
C5348 VCC.t0 VSS 0.00366f 
C5349 VCC.t26 VSS 0.00365f 
C5350 VCC.t1 VSS 0.00386f 
C5351 VCC.n1536 VSS 0.00569f 
C5352 VCC.n1537 VSS 1.3e-19 
C5353 VCC.n1538 VSS 3.67e-19 
C5354 VCC.n1539 VSS 1.15e-19 
C5355 VCC.n1540 VSS 3.38e-19 
C5356 VCC.n1541 VSS 3.5e-20 
C5357 VCC.n1542 VSS 3.5e-20 
C5358 VCC.n1543 VSS 2.68e-20 
C5359 VCC.n1544 VSS 2.06e-20 
C5360 VCC.n1545 VSS 6.38e-20 
C5361 VCC.n1546 VSS 5.97e-20 
C5362 VCC.n1547 VSS 4.73e-20 
C5363 VCC.n1548 VSS 4.73e-20 
C5364 VCC.n1549 VSS 3.09e-20 
C5365 VCC.n1550 VSS 1.23e-20 
C5366 VCC.n1551 VSS 1.65e-20 
C5367 VCC.n1552 VSS 1.54e-19 
C5368 VCC.n1553 VSS 1.54e-19 
C5369 VCC.n1554 VSS 1.65e-20 
C5370 VCC.n1555 VSS 3.29e-20 
C5371 VCC.t256 VSS 1.67e-19 
C5372 VCC.n1556 VSS 0.00101f 
C5373 VCC.n1557 VSS 2.71e-19 
C5374 VCC.n1558 VSS 7.46e-19 
C5375 VCC.n1559 VSS 0.00333f 
C5376 VCC.n1560 VSS 2.46e-19 
C5377 VCC.n1561 VSS 3.02e-19 
C5378 VCC.n1562 VSS 3.7e-20 
C5379 VCC.n1563 VSS 5.15e-20 
C5380 VCC.n1564 VSS 5.97e-20 
C5381 VCC.n1565 VSS 6.38e-20 
C5382 VCC.n1566 VSS 4.73e-20 
C5383 VCC.n1567 VSS 4.73e-20 
C5384 VCC.n1568 VSS 2.68e-20 
C5385 VCC.n1569 VSS 3.29e-20 
C5386 VCC.n1570 VSS 1.65e-20 
C5387 VCC.n1571 VSS 1.54e-19 
C5388 VCC.n1572 VSS 1.54e-19 
C5389 VCC.n1573 VSS 1.65e-20 
C5390 VCC.n1574 VSS 3.09e-20 
C5391 VCC.n1575 VSS 3.09e-20 
C5392 VCC.n1576 VSS 4.73e-20 
C5393 VCC.n1577 VSS 4.32e-20 
C5394 VCC.n1578 VSS 3.5e-20 
C5395 VCC.n1579 VSS 3.5e-20 
C5396 VCC.n1580 VSS 1.35e-19 
C5397 VCC.n1581 VSS 5.24e-19 
C5398 VCC.n1582 VSS 1.4e-19 
C5399 VCC.n1583 VSS 5.4e-19 
C5400 VCC.n1584 VSS 1.35e-19 
C5401 VCC.n1585 VSS 4.37e-19 
C5402 VCC.n1586 VSS 1.13e-19 
C5403 VCC.n1587 VSS 8.23e-21 
C5404 VCC.n1588 VSS 1.65e-20 
C5405 VCC.n1589 VSS 3.5e-20 
C5406 VCC.n1590 VSS 3.91e-20 
C5407 VCC.n1591 VSS 3.09e-20 
C5408 VCC.n1592 VSS 1.85e-20 
C5409 VCC.n1593 VSS 3.5e-20 
C5410 VCC.n1594 VSS 1.05e-19 
C5411 VCC.n1595 VSS 2.06e-20 
C5412 VCC.n1596 VSS 2.26e-20 
C5413 VCC.n1597 VSS 3.7e-20 
C5414 VCC.n1598 VSS 5.15e-20 
C5415 VCC.n1599 VSS 1.38e-19 
C5416 VCC.n1600 VSS 1.17e-19 
C5417 VCC.n1601 VSS 4.32e-20 
C5418 VCC.n1602 VSS 2.88e-20 
C5419 VCC.n1603 VSS 2.68e-20 
C5420 VCC.n1604 VSS 6.59e-20 
C5421 VCC.n1605 VSS 5.56e-20 
C5422 VCC.n1606 VSS 2.68e-20 
C5423 VCC.n1607 VSS 4.32e-20 
C5424 VCC.n1608 VSS 1.05e-19 
C5425 VCC.n1609 VSS 3.09e-20 
C5426 VCC.n1610 VSS 3.7e-20 
C5427 VCC.n1611 VSS 4.32e-20 
C5428 VCC.n1612 VSS 1.05e-19 
C5429 VCC.n1613 VSS 4.53e-20 
C5430 VCC.n1614 VSS 4.53e-20 
C5431 VCC.n1615 VSS 7.82e-20 
C5432 VCC.n1616 VSS 2.18e-19 
C5433 VCC.n1617 VSS 1.4e-19 
C5434 VCC.n1618 VSS 1.4e-19 
C5435 VCC.n1619 VSS 5.4e-19 
C5436 VCC.n1620 VSS 1.35e-19 
C5437 VCC.t134 VSS 4.21e-19 
C5438 VCC.n1621 VSS 3.33e-19 
C5439 VCC.n1622 VSS 1.13e-19 
C5440 VCC.n1623 VSS 8.23e-21 
C5441 VCC.n1624 VSS 1.65e-20 
C5442 VCC.n1625 VSS 3.5e-20 
C5443 VCC.n1626 VSS 3.5e-20 
C5444 VCC.n1627 VSS 3.5e-20 
C5445 VCC.n1628 VSS 1.17e-19 
C5446 VCC.n1629 VSS 1.38e-19 
C5447 VCC.n1630 VSS 5.15e-20 
C5448 VCC.n1631 VSS 4.73e-20 
C5449 VCC.n1632 VSS 7.2e-20 
C5450 VCC.n1633 VSS 2.68e-20 
C5451 VCC.n1634 VSS 1.65e-20 
C5452 VCC.n1635 VSS 1.54e-19 
C5453 VCC.n1636 VSS 1.54e-19 
C5454 VCC.n1637 VSS 1.65e-20 
C5455 VCC.n1638 VSS 2.47e-20 
C5456 VCC.n1639 VSS 1.23e-20 
C5457 VCC.n1640 VSS 7.62e-19 
C5458 VCC.n1641 VSS 4.12e-20 
C5459 VCC.n1642 VSS 5.15e-20 
C5460 VCC.n1643 VSS 6.59e-20 
C5461 VCC.n1644 VSS 5.76e-20 
C5462 VCC.n1645 VSS 4.73e-20 
C5463 VCC.n1646 VSS 2.26e-20 
C5464 VCC.n1647 VSS 2.68e-20 
C5465 VCC.n1648 VSS 1.03e-20 
C5466 VCC.n1649 VSS 3.5e-20 
C5467 VCC.n1650 VSS 3.5e-20 
C5468 VCC.n1651 VSS 1.35e-19 
C5469 VCC.n1652 VSS 4.53e-19 
C5470 VCC.n1653 VSS 7.71e-19 
C5471 VCC.n1654 VSS 1.32e-19 
C5472 VCC.n1655 VSS 3.5e-20 
C5473 VCC.n1656 VSS 3.42e-20 
C5474 VCC.n1657 VSS 2.36e-19 
C5475 VCC.n1658 VSS 3.21e-19 
C5476 VCC.n1659 VSS 2.61e-19 
C5477 VCC.n1660 VSS 0.00189f 
C5478 VCC.n1661 VSS 2.68e-19 
C5479 VCC.n1662 VSS 0.00246f 
C5480 VCC.n1663 VSS 5.76e-20 
C5481 VCC.n1664 VSS 2.88e-20 
C5482 VCC.n1665 VSS 3.5e-20 
C5483 VCC.n1666 VSS 3.42e-20 
C5484 VCC.n1667 VSS 3.5e-20 
C5485 VCC.n1668 VSS 4.53e-19 
C5486 VCC.n1669 VSS 1.17e-19 
C5487 VCC.n1670 VSS 3.5e-20 
C5488 VCC.n1671 VSS 1.44e-20 
C5489 VCC.n1672 VSS 4.12e-20 
C5490 VCC.n1673 VSS 5.76e-20 
C5491 VCC.n1674 VSS 5.76e-20 
C5492 VCC.n1675 VSS 2.06e-20 
C5493 VCC.n1676 VSS 3.29e-20 
C5494 VCC.n1677 VSS 7.2e-20 
C5495 VCC.n1678 VSS 3.29e-20 
C5496 VCC.n1679 VSS 4.73e-20 
C5497 VCC.n1680 VSS 2.26e-20 
C5498 VCC.n1681 VSS 1.01e-19 
C5499 VCC.n1682 VSS 1.36e-19 
C5500 VCC.n1683 VSS 1.35e-19 
C5501 VCC.n1684 VSS 3.5e-20 
C5502 VCC.n1685 VSS 3.5e-20 
C5503 VCC.n1686 VSS 3.5e-20 
C5504 VCC.n1687 VSS 3.5e-20 
C5505 VCC.n1688 VSS 3.09e-20 
C5506 VCC.n1689 VSS 3.91e-20 
C5507 VCC.n1690 VSS 4.73e-20 
C5508 VCC.n1691 VSS 4.32e-20 
C5509 VCC.n1692 VSS 2.68e-20 
C5510 VCC.n1693 VSS 4.53e-20 
C5511 VCC.n1694 VSS 4.53e-20 
C5512 VCC.n1695 VSS 3.09e-20 
C5513 VCC.n1696 VSS 4.32e-20 
C5514 VCC.n1697 VSS 2.68e-20 
C5515 VCC.n1698 VSS 7.82e-20 
C5516 VCC.n1699 VSS 5.56e-20 
C5517 VCC.n1700 VSS 1.4e-19 
C5518 VCC.n1701 VSS 2.18e-19 
C5519 VCC.n1702 VSS 1.35e-19 
C5520 VCC.n1703 VSS 1.13e-19 
C5521 VCC.n1704 VSS 3.5e-20 
C5522 VCC.n1705 VSS 1.85e-20 
C5523 VCC.n1706 VSS 3.7e-20 
C5524 VCC.n1707 VSS 3.09e-20 
C5525 VCC.n1708 VSS 6.59e-20 
C5526 VCC.n1709 VSS 2.68e-20 
C5527 VCC.n1710 VSS 5.76e-20 
C5528 VCC.n1711 VSS 4.73e-20 
C5529 VCC.n1712 VSS 3.5e-20 
C5530 VCC.t22 VSS 1.56e-19 
C5531 VCC.n1713 VSS 7.97e-19 
C5532 VCC.n1714 VSS 3.09e-20 
C5533 VCC.n1715 VSS 3.5e-20 
C5534 VCC.n1716 VSS 3.5e-20 
C5535 VCC.t21 VSS 4.21e-19 
C5536 VCC.n1717 VSS 1.32e-19 
C5537 VCC.n1718 VSS 1.09e-19 
C5538 VCC.n1719 VSS 3.5e-20 
C5539 VCC.n1720 VSS 3.09e-20 
C5540 VCC.n1721 VSS 5.97e-20 
C5541 VCC.n1722 VSS 2.26e-20 
C5542 VCC.n1723 VSS 5.76e-20 
C5543 VCC.n1724 VSS 2.68e-20 
C5544 VCC.n1725 VSS 2.68e-20 
C5545 VCC.n1726 VSS 1.9e-19 
C5546 VCC.n1727 VSS 5.76e-20 
C5547 VCC.n1728 VSS 2.68e-20 
C5548 VCC.n1729 VSS 2.68e-20 
C5549 VCC.n1730 VSS 2.68e-20 
C5550 VCC.n1731 VSS 5.76e-20 
C5551 VCC.n1732 VSS 2.26e-20 
C5552 VCC.n1733 VSS 3.09e-20 
C5553 VCC.n1734 VSS 2.26e-20 
C5554 VCC.n1735 VSS 5.15e-20 
C5555 VCC.n1736 VSS 4.73e-20 
C5556 VCC.n1737 VSS 3.7e-20 
C5557 VCC.n1738 VSS 3.5e-20 
C5558 VCC.n1739 VSS 7.41e-20 
C5559 VCC.n1740 VSS 1.91e-19 
C5560 VCC.n1741 VSS 9.88e-20 
C5561 VCC.n1742 VSS 3e-20 
C5562 VCC.n1743 VSS 5.12e-19 
C5563 VCC.n1744 VSS 1.18e-19 
C5564 VCC.n1745 VSS 3.5e-20 
C5565 VCC.n1746 VSS 3.5e-20 
C5566 VCC.n1747 VSS 5.15e-20 
C5567 VCC.n1748 VSS 4.32e-20 
C5568 VCC.n1749 VSS 2.68e-20 
C5569 VCC.n1750 VSS 3.91e-20 
C5570 VCC.n1751 VSS 1.44e-20 
C5571 VCC.n1752 VSS 3.5e-20 
C5572 VCC.n1753 VSS 3e-20 
C5573 VCC.n1754 VSS 7.95e-19 
C5574 VCC.n1755 VSS 1.83e-19 
C5575 VCC.n1756 VSS 2.88e-20 
C5576 VCC.n1757 VSS 2.68e-20 
C5577 VCC.n1758 VSS 2.68e-20 
C5578 VCC.n1759 VSS 2.68e-20 
C5579 VCC.n1760 VSS 4.53e-20 
C5580 VCC.n1761 VSS 3.7e-20 
C5581 VCC.n1762 VSS 7.82e-20 
C5582 VCC.n1763 VSS 1.17e-19 
C5583 VCC.n1764 VSS 3.91e-20 
C5584 VCC.n1765 VSS 1.65e-20 
C5585 VCC.n1766 VSS 2.68e-20 
C5586 VCC.n1767 VSS 3.5e-20 
C5587 VCC.n1768 VSS 3e-20 
C5588 VCC.n1769 VSS 5.12e-19 
C5589 VCC.n1770 VSS 1.18e-19 
C5590 VCC.n1771 VSS 3.5e-20 
C5591 VCC.n1772 VSS 3.5e-20 
C5592 VCC.t51 VSS 1.55e-19 
C5593 VCC.n1773 VSS 7.57e-19 
C5594 VCC.n1774 VSS 4.73e-20 
C5595 VCC.n1775 VSS 1.54e-19 
C5596 VCC.n1776 VSS 2.88e-20 
C5597 VCC.n1777 VSS 2.88e-20 
C5598 VCC.n1778 VSS 3.5e-20 
C5599 VCC.n1779 VSS 5.76e-20 
C5600 VCC.n1780 VSS 9.88e-20 
C5601 VCC.n1781 VSS 1.3e-19 
C5602 VCC.n1782 VSS 3e-20 
C5603 VCC.t49 VSS 0.005f 
C5604 VCC.t145 VSS 0.00453f 
C5605 VCC.n1783 VSS 0.00229f 
C5606 VCC.n1784 VSS 1.91e-19 
C5607 VCC.n1785 VSS 3.5e-20 
C5608 VCC.n1786 VSS 3.14e-19 
C5609 VCC.n1787 VSS 2.47e-20 
C5610 VCC.n1788 VSS 5.76e-20 
C5611 VCC.n1789 VSS 2.47e-20 
C5612 VCC.n1790 VSS 8.23e-21 
C5613 VCC.n1791 VSS 2.88e-20 
C5614 VCC.n1792 VSS 5.76e-20 
C5615 VCC.n1793 VSS 2.47e-20 
C5616 VCC.n1794 VSS 2.88e-20 
C5617 VCC.n1795 VSS 2.47e-20 
C5618 VCC.n1796 VSS 5.15e-20 
C5619 VCC.n1797 VSS 4.73e-20 
C5620 VCC.n1798 VSS 3.7e-20 
C5621 VCC.n1799 VSS 3.5e-20 
C5622 VCC.n1800 VSS 7.41e-20 
C5623 VCC.t76 VSS 6.42e-19 
C5624 VCC.n1801 VSS 3e-20 
C5625 VCC.n1802 VSS 5.97e-20 
C5626 VCC.n1803 VSS 4.13e-19 
C5627 VCC.n1804 VSS 9.53e-20 
C5628 VCC.n1805 VSS 3.5e-20 
C5629 VCC.n1806 VSS 3.5e-20 
C5630 VCC.n1807 VSS 5.35e-20 
C5631 VCC.n1808 VSS 4.32e-20 
C5632 VCC.n1809 VSS 2.68e-20 
C5633 VCC.n1810 VSS 3.7e-20 
C5634 VCC.n1811 VSS 1.65e-20 
C5635 VCC.n1812 VSS 4.53e-20 
C5636 VCC.n1813 VSS 1.2e-19 
C5637 VCC.n1814 VSS 5.2e-19 
C5638 VCC.n1815 VSS 1.2e-19 
C5639 VCC.n1816 VSS 6.38e-20 
C5640 VCC.n1817 VSS 2.47e-20 
C5641 VCC.n1818 VSS 4.53e-20 
C5642 VCC.n1819 VSS 3.5e-20 
C5643 VCC.n1820 VSS 3.5e-20 
C5644 VCC.n1821 VSS 2.68e-20 
C5645 VCC.n1822 VSS 2.68e-20 
C5646 VCC.n1823 VSS 2.47e-20 
C5647 VCC.n1824 VSS 4.53e-20 
C5648 VCC.n1825 VSS 2.68e-20 
C5649 VCC.n1826 VSS 4.32e-20 
C5650 VCC.n1827 VSS 2.68e-20 
C5651 VCC.n1828 VSS 3.91e-20 
C5652 VCC.n1829 VSS 2.88e-20 
C5653 VCC.n1830 VSS 4.73e-20 
C5654 VCC.n1831 VSS 3.7e-20 
C5655 VCC.n1832 VSS 3.7e-20 
C5656 VCC.n1833 VSS 3.5e-20 
C5657 VCC.n1834 VSS 5.76e-20 
C5658 VCC.n1835 VSS 4.73e-20 
C5659 VCC.n1836 VSS 3.09e-20 
C5660 VCC.n1837 VSS 3.5e-20 
C5661 VCC.n1838 VSS 3.5e-20 
C5662 VCC.n1839 VSS 3.5e-20 
C5663 VCC.n1840 VSS 1.18e-19 
C5664 VCC.n1841 VSS 3e-20 
C5665 VCC.n1842 VSS 1.15e-19 
C5666 VCC.n1843 VSS 9.88e-20 
C5667 VCC.n1844 VSS 5.76e-20 
C5668 VCC.n1845 VSS 3.5e-20 
C5669 VCC.n1846 VSS 3.09e-20 
C5670 VCC.n1847 VSS 3.09e-20 
C5671 VCC.n1848 VSS 2.26e-20 
C5672 VCC.n1849 VSS 5.76e-20 
C5673 VCC.n1850 VSS 2.68e-20 
C5674 VCC.n1851 VSS 2.68e-20 
C5675 VCC.n1852 VSS 0.00185f 
C5676 VCC.n1853 VSS 2.72e-19 
C5677 VCC.n1854 VSS 2.26e-20 
C5678 VCC.n1855 VSS 1.87e-19 
C5679 VCC.n1856 VSS 3.5e-20 
C5680 VCC.n1857 VSS 2.68e-20 
C5681 VCC.n1858 VSS 5.97e-20 
C5682 VCC.n1859 VSS 4.73e-20 
C5683 VCC.n1860 VSS 4.73e-20 
C5684 VCC.n1861 VSS 5.15e-20 
C5685 VCC.n1862 VSS 7.41e-20 
C5686 VCC.n1863 VSS 3.7e-20 
C5687 VCC.n1864 VSS 2.26e-20 
C5688 VCC.n1865 VSS 6.38e-20 
C5689 VCC.n1866 VSS 4.73e-20 
C5690 VCC.n1867 VSS 3.29e-20 
C5691 VCC.n1868 VSS 3.5e-20 
C5692 VCC.n1869 VSS 3e-20 
C5693 VCC.t210 VSS 0.005f 
C5694 VCC.t90 VSS 0.00453f 
C5695 VCC.n1870 VSS 0.00228f 
C5696 VCC.n1871 VSS 1.3e-19 
C5697 VCC.t208 VSS 4.05e-19 
C5698 VCC.n1872 VSS 4.05e-19 
C5699 VCC.n1873 VSS 1.15e-19 
C5700 VCC.n1874 VSS 3.36e-19 
C5701 VCC.n1875 VSS 6.17e-21 
C5702 VCC.n1876 VSS 3.12e-19 
C5703 VCC.n1877 VSS 1.65e-20 
C5704 VCC.n1878 VSS 1.54e-19 
C5705 VCC.n1879 VSS 1.54e-19 
C5706 VCC.n1880 VSS 1.65e-20 
C5707 VCC.n1881 VSS 1.03e-20 
C5708 VCC.n1882 VSS 3.5e-20 
C5709 VCC.n1883 VSS 2.26e-20 
C5710 VCC.n1884 VSS 4.73e-20 
C5711 VCC.n1885 VSS 3.5e-20 
C5712 VCC.n1886 VSS 3e-20 
C5713 VCC.n1887 VSS 1.3e-19 
C5714 VCC.n1888 VSS 5.12e-19 
C5715 VCC.n1889 VSS 1.3e-19 
C5716 VCC.n1890 VSS 4.13e-19 
C5717 VCC.n1891 VSS 9.53e-20 
C5718 VCC.n1892 VSS 5.76e-20 
C5719 VCC.n1893 VSS 7.41e-20 
C5720 VCC.n1894 VSS 5.56e-20 
C5721 VCC.t209 VSS 1.55e-19 
C5722 VCC.n1895 VSS 3.91e-20 
C5723 VCC.n1896 VSS 3.91e-20 
C5724 VCC.n1897 VSS 1.85e-20 
C5725 VCC.n1898 VSS 7.55e-19 
C5726 VCC.n1899 VSS 4.94e-20 
C5727 VCC.n1900 VSS 5.15e-20 
C5728 VCC.n1901 VSS 7.2e-20 
C5729 VCC.n1902 VSS 1.38e-19 
C5730 VCC.n1903 VSS 1.17e-19 
C5731 VCC.n1904 VSS 4.32e-20 
C5732 VCC.n1905 VSS 2.88e-20 
C5733 VCC.n1906 VSS 2.68e-20 
C5734 VCC.n1907 VSS 3.5e-20 
C5735 VCC.n1908 VSS 3.5e-20 
C5736 VCC.n1909 VSS 2.88e-20 
C5737 VCC.n1910 VSS 2.68e-20 
C5738 VCC.n1911 VSS 2.68e-20 
C5739 VCC.n1912 VSS 2.68e-20 
C5740 VCC.n1913 VSS 4.12e-20 
C5741 VCC.n1914 VSS 4.12e-20 
C5742 VCC.n1915 VSS 3.91e-20 
C5743 VCC.n1916 VSS 4.53e-20 
C5744 VCC.n1917 VSS 4.53e-20 
C5745 VCC.n1918 VSS 1.05e-19 
C5746 VCC.n1919 VSS 1.05e-19 
C5747 VCC.n1920 VSS 4.32e-20 
C5748 VCC.n1921 VSS 3.7e-20 
C5749 VCC.n1922 VSS 2.68e-20 
C5750 VCC.n1923 VSS 2.68e-20 
C5751 VCC.n1924 VSS 6.79e-20 
C5752 VCC.n1925 VSS 9.26e-20 
C5753 VCC.n1926 VSS 1.83e-19 
C5754 VCC.n1927 VSS 7.95e-19 
C5755 VCC.n1928 VSS 5.2e-19 
C5756 VCC.n1929 VSS 1.3e-19 
C5757 VCC.n1930 VSS 3e-20 
C5758 VCC.n1931 VSS 3.5e-20 
C5759 VCC.n1932 VSS 5.97e-20 
C5760 VCC.n1933 VSS 7.41e-20 
C5761 VCC.n1934 VSS 5.15e-20 
C5762 VCC.n1935 VSS 5.15e-20 
C5763 VCC.n1936 VSS 3.09e-20 
C5764 VCC.n1937 VSS 3.09e-20 
C5765 VCC.n1938 VSS 3.7e-20 
C5766 VCC.n1939 VSS 2.68e-20 
C5767 VCC.n1940 VSS 3.91e-20 
C5768 VCC.n1941 VSS 1.17e-19 
C5769 VCC.n1942 VSS 1.38e-19 
C5770 VCC.n1943 VSS 7e-20 
C5771 VCC.n1944 VSS 4.73e-20 
C5772 VCC.n1945 VSS 3.5e-20 
C5773 VCC.n1946 VSS 3.5e-20 
C5774 VCC.n1947 VSS 3.5e-20 
C5775 VCC.n1948 VSS 4.53e-20 
C5776 VCC.n1949 VSS 1.18e-19 
C5777 VCC.n1950 VSS 5.12e-19 
C5778 VCC.n1951 VSS 1.3e-19 
C5779 VCC.n1952 VSS 1.61e-19 
C5780 VCC.n1953 VSS 9.9e-20 
C5781 VCC.n1954 VSS 0.00243f 
C5782 VCC.n1955 VSS 2.26e-20 
C5783 VCC.n1956 VSS 4.13e-19 
C5784 VCC.n1957 VSS 3.5e-20 
C5785 VCC.n1958 VSS 3.5e-20 
C5786 VCC.n1959 VSS 2.47e-20 
C5787 VCC.n1960 VSS 2.06e-20 
C5788 VCC.n1961 VSS 6.17e-20 
C5789 VCC.n1962 VSS 6.17e-20 
C5790 VCC.n1963 VSS 4.73e-20 
C5791 VCC.n1964 VSS 4.73e-20 
C5792 VCC.n1965 VSS 2.88e-20 
C5793 VCC.n1966 VSS 1.44e-20 
C5794 VCC.n1967 VSS 1.65e-20 
C5795 VCC.n1968 VSS 1.54e-19 
C5796 VCC.n1969 VSS 1.54e-19 
C5797 VCC.n1970 VSS 1.65e-20 
C5798 VCC.n1971 VSS 3.09e-20 
C5799 VCC.t77 VSS 1.55e-19 
C5800 VCC.n1972 VSS 0.00102f 
C5801 VCC.n1973 VSS 2.73e-19 
C5802 VCC.n1974 VSS 0.00136f 
C5803 VCC.n1975 VSS 2.73e-19 
C5804 VCC.n1976 VSS 0.00181f 
C5805 VCC.n1977 VSS 5.76e-20 
C5806 VCC.n1978 VSS 1.54e-19 
C5807 VCC.n1979 VSS 1.65e-20 
C5808 VCC.n1980 VSS 2.88e-20 
C5809 VCC.n1981 VSS 2.47e-20 
C5810 VCC.n1982 VSS 6.17e-20 
C5811 VCC.n1983 VSS 4.73e-20 
C5812 VCC.n1984 VSS 4.73e-20 
C5813 VCC.n1985 VSS 5.15e-20 
C5814 VCC.n1986 VSS 3.5e-20 
C5815 VCC.n1987 VSS 7.41e-20 
C5816 VCC.n1988 VSS 3.7e-20 
C5817 VCC.n1989 VSS 2.26e-20 
C5818 VCC.n1990 VSS 6.17e-20 
C5819 VCC.n1991 VSS 4.73e-20 
C5820 VCC.n1992 VSS 3.5e-20 
C5821 VCC.n1993 VSS 2.88e-20 
C5822 VCC.n1994 VSS 3.4e-19 
C5823 VCC.n1995 VSS 1.15e-19 
C5824 VCC.n1996 VSS 3.98e-19 
C5825 VCC.t50 VSS 4.05e-19 
C5826 VCC.n1997 VSS 1.22e-19 
C5827 VCC.n1998 VSS 1.3e-19 
C5828 VCC.n1999 VSS 3e-20 
C5829 VCC.n2000 VSS 3.5e-20 
C5830 VCC.n2001 VSS 3.5e-20 
C5831 VCC.n2002 VSS 4.73e-20 
C5832 VCC.n2003 VSS 2.47e-20 
C5833 VCC.n2004 VSS 1.23e-20 
C5834 VCC.n2005 VSS 1.65e-20 
C5835 VCC.n2006 VSS 2.47e-20 
C5836 VCC.n2007 VSS 5.76e-20 
C5837 VCC.n2008 VSS 1.38e-19 
C5838 VCC.n2009 VSS 7e-20 
C5839 VCC.n2010 VSS 3.7e-20 
C5840 VCC.n2011 VSS 2.47e-20 
C5841 VCC.n2012 VSS 3.7e-20 
C5842 VCC.n2013 VSS 1.85e-20 
C5843 VCC.n2014 VSS 3.09e-20 
C5844 VCC.n2015 VSS 5.35e-20 
C5845 VCC.n2016 VSS 4.73e-20 
C5846 VCC.n2017 VSS 5.35e-20 
C5847 VCC.n2018 VSS 7.41e-20 
C5848 VCC.n2019 VSS 5.76e-20 
C5849 VCC.n2020 VSS 9.53e-20 
C5850 VCC.n2021 VSS 4.13e-19 
C5851 VCC.n2022 VSS 1.3e-19 
C5852 VCC.n2023 VSS 5.2e-19 
C5853 VCC.n2024 VSS 1.2e-19 
C5854 VCC.n2025 VSS 4.73e-20 
C5855 VCC.n2026 VSS 2.68e-20 
C5856 VCC.n2027 VSS 3.5e-20 
C5857 VCC.n2028 VSS 3.5e-20 
C5858 VCC.n2029 VSS 2.68e-20 
C5859 VCC.n2030 VSS 2.68e-20 
C5860 VCC.n2031 VSS 4.32e-20 
C5861 VCC.n2032 VSS 4.32e-20 
C5862 VCC.n2033 VSS 4.32e-20 
C5863 VCC.n2034 VSS 2.88e-20 
C5864 VCC.n2035 VSS 3.5e-20 
C5865 VCC.n2036 VSS 2.68e-20 
C5866 VCC.n2037 VSS 7.82e-20 
C5867 VCC.n2038 VSS 4.73e-20 
C5868 VCC.n2039 VSS 4.73e-20 
C5869 VCC.n2040 VSS 1.05e-19 
C5870 VCC.n2041 VSS 1.05e-19 
C5871 VCC.n2042 VSS 4.53e-20 
C5872 VCC.n2043 VSS 2.68e-20 
C5873 VCC.n2044 VSS 2.68e-20 
C5874 VCC.n2045 VSS 6.59e-20 
C5875 VCC.n2046 VSS 9.26e-20 
C5876 VCC.n2047 VSS 6.59e-20 
C5877 VCC.n2048 VSS 2.47e-20 
C5878 VCC.n2049 VSS 2.47e-20 
C5879 VCC.n2050 VSS 2.88e-20 
C5880 VCC.n2051 VSS 3.5e-20 
C5881 VCC.n2052 VSS 3.5e-20 
C5882 VCC.n2053 VSS 4.53e-20 
C5883 VCC.n2054 VSS 1.2e-19 
C5884 VCC.n2055 VSS 5.2e-19 
C5885 VCC.n2056 VSS 1.3e-19 
C5886 VCC.n2057 VSS 4.13e-19 
C5887 VCC.n2058 VSS 9.53e-20 
C5888 VCC.n2059 VSS 5.97e-20 
C5889 VCC.n2060 VSS 7.41e-20 
C5890 VCC.n2061 VSS 5.35e-20 
C5891 VCC.n2062 VSS 5.15e-20 
C5892 VCC.n2063 VSS 3.09e-20 
C5893 VCC.n2064 VSS 3.09e-20 
C5894 VCC.n2065 VSS 3.91e-20 
C5895 VCC.n2066 VSS 2.47e-20 
C5896 VCC.n2067 VSS 3.7e-20 
C5897 VCC.n2068 VSS 1.17e-19 
C5898 VCC.n2069 VSS 1.38e-19 
C5899 VCC.n2070 VSS 7.2e-20 
C5900 VCC.n2071 VSS 4.73e-20 
C5901 VCC.n2072 VSS 3.5e-20 
C5902 VCC.n2073 VSS 3.5e-20 
C5903 VCC.n2074 VSS 4.53e-20 
C5904 VCC.n2075 VSS 5.97e-20 
C5905 VCC.n2076 VSS 3.5e-20 
C5906 VCC.n2077 VSS 3e-20 
C5907 VCC.n2078 VSS 1.3e-19 
C5908 VCC.n2079 VSS 1.53e-19 
C5909 VCC.t18 VSS 4.05e-19 
C5910 VCC.n2080 VSS 2.06e-19 
C5911 VCC.n2081 VSS 1.35e-19 
C5912 VCC.n2082 VSS 9.67e-20 
C5913 VCC.n2083 VSS 3.35e-20 
C5914 VCC.n2084 VSS 3.5e-20 
C5915 VCC.n2085 VSS 2.36e-19 
C5916 VCC.n2086 VSS 0.0023f 
C5917 VCC.t20 VSS 0.0031f 
C5918 VCC.t44 VSS 0.00366f 
C5919 VCC.t23 VSS 0.00365f 
C5920 VCC.t47 VSS 0.00386f 
C5921 VCC.n2087 VSS 0.00569f 
C5922 VCC.n2088 VSS 1.3e-19 
C5923 VCC.n2089 VSS 3.67e-19 
C5924 VCC.n2090 VSS 1.15e-19 
C5925 VCC.n2091 VSS 3.38e-19 
C5926 VCC.n2092 VSS 3.5e-20 
C5927 VCC.n2093 VSS 3.5e-20 
C5928 VCC.n2094 VSS 2.68e-20 
C5929 VCC.n2095 VSS 2.06e-20 
C5930 VCC.n2096 VSS 6.38e-20 
C5931 VCC.n2097 VSS 5.97e-20 
C5932 VCC.n2098 VSS 4.73e-20 
C5933 VCC.n2099 VSS 4.73e-20 
C5934 VCC.n2100 VSS 3.09e-20 
C5935 VCC.n2101 VSS 1.23e-20 
C5936 VCC.n2102 VSS 1.65e-20 
C5937 VCC.n2103 VSS 1.54e-19 
C5938 VCC.n2104 VSS 1.54e-19 
C5939 VCC.n2105 VSS 1.65e-20 
C5940 VCC.n2106 VSS 3.29e-20 
C5941 VCC.t19 VSS 1.67e-19 
C5942 VCC.n2107 VSS 0.00101f 
C5943 VCC.n2108 VSS 2.71e-19 
C5944 VCC.n2109 VSS 7.46e-19 
C5945 VCC.n2110 VSS 0.00333f 
C5946 VCC.n2111 VSS 2.46e-19 
C5947 VCC.n2112 VSS 3.02e-19 
C5948 VCC.n2113 VSS 3.7e-20 
C5949 VCC.n2114 VSS 5.15e-20 
C5950 VCC.n2115 VSS 6.38e-20 
C5951 VCC.n2116 VSS 4.73e-20 
C5952 VCC.n2117 VSS 4.73e-20 
C5953 VCC.n2118 VSS 2.68e-20 
C5954 VCC.n2119 VSS 3.29e-20 
C5955 VCC.n2120 VSS 1.65e-20 
C5956 VCC.n2121 VSS 1.54e-19 
C5957 VCC.n2122 VSS 1.54e-19 
C5958 VCC.n2123 VSS 5.56e-20 
C5959 VCC.n2124 VSS 2.88e-20 
C5960 VCC.n2125 VSS 1.65e-20 
C5961 VCC.n2126 VSS 3.09e-20 
C5962 VCC.n2127 VSS 4.73e-20 
C5963 VCC.n2128 VSS 4.73e-20 
C5964 VCC.n2129 VSS 4.32e-20 
C5965 VCC.n2130 VSS 1.17e-19 
C5966 VCC.n2131 VSS 3.33e-19 
C5967 VCC.n2132 VSS 1.35e-19 
C5968 VCC.n2133 VSS 4.37e-19 
C5969 VCC.n2134 VSS 5.24e-19 
C5970 VCC.n2135 VSS 1.36e-19 
C5971 VCC.n2136 VSS 1.01e-19 
C5972 VCC.n2137 VSS 1.05e-19 
C5973 VCC.n2138 VSS 2.06e-20 
C5974 VCC.n2139 VSS 2.26e-20 
C5975 VCC.n2140 VSS 3.7e-20 
C5976 VCC.n2141 VSS 5.15e-20 
C5977 VCC.n2142 VSS 1.38e-19 
C5978 VCC.n2143 VSS 3.91e-20 
C5979 VCC.n2144 VSS 2.88e-20 
C5980 VCC.n2145 VSS 4.32e-20 
C5981 VCC.n2146 VSS 1.17e-19 
C5982 VCC.n2147 VSS 3.7e-20 
C5983 VCC.n2148 VSS 3.91e-20 
C5984 VCC.n2149 VSS 3.5e-20 
C5985 VCC.n2150 VSS 1.65e-20 
C5986 VCC.n2151 VSS 8.23e-21 
C5987 VCC.n2152 VSS 3.5e-20 
C5988 VCC.n2153 VSS 3.5e-20 
C5989 VCC.n2154 VSS 1.4e-19 
C5990 VCC.n2155 VSS 5.4e-19 
C5991 VCC.n2156 VSS 8.42e-19 
C5992 VCC.n2157 VSS 5.4e-19 
C5993 VCC.n2158 VSS 1.4e-19 
C5994 VCC.n2159 VSS 1.4e-19 
C5995 VCC.n2160 VSS 2.18e-19 
C5996 VCC.n2161 VSS 7.82e-20 
C5997 VCC.n2162 VSS 4.32e-20 
C5998 VCC.n2163 VSS 4.32e-20 
C5999 VCC.n2164 VSS 1.05e-19 
C6000 VCC.n2165 VSS 1.05e-19 
C6001 VCC.n2166 VSS 4.32e-20 
C6002 VCC.n2167 VSS 3.7e-20 
C6003 VCC.n2168 VSS 2.68e-20 
C6004 VCC.n2169 VSS 5.76e-20 
C6005 VCC.n2170 VSS 6.38e-20 
C6006 VCC.n2171 VSS 3.5e-20 
C6007 VCC.n2172 VSS 3.5e-20 
C6008 VCC.n2173 VSS 1.17e-19 
C6009 VCC.n2174 VSS 1.38e-19 
C6010 VCC.n2175 VSS 5.15e-20 
C6011 VCC.n2176 VSS 1.05e-19 
C6012 VCC.n2177 VSS 2.26e-20 
C6013 VCC.n2178 VSS 5.76e-20 
C6014 VCC.n2179 VSS 3.7e-20 
C6015 VCC.n2180 VSS 3.7e-20 
C6016 VCC.n2181 VSS 3.09e-20 
C6017 VCC.n2182 VSS 1.85e-20 
C6018 VCC.n2183 VSS 1.65e-20 
C6019 VCC.n2184 VSS 8.23e-21 
C6020 VCC.n2185 VSS 1.13e-19 
C6021 VCC.n2186 VSS 3.33e-19 
C6022 VCC.t2 VSS 4.21e-19 
C6023 VCC.n2187 VSS 2.06e-19 
C6024 VCC.n2188 VSS 1.35e-19 
C6025 VCC.n2189 VSS 3.5e-20 
C6026 VCC.n2190 VSS 3.5e-20 
C6027 VCC.n2191 VSS 3.5e-20 
C6028 VCC.n2192 VSS 1.03e-20 
C6029 VCC.n2193 VSS 2.68e-20 
C6030 VCC.n2194 VSS 3.09e-20 
C6031 VCC.n2195 VSS 2.68e-20 
C6032 VCC.n2196 VSS 1.65e-20 
C6033 VCC.n2197 VSS 1.54e-19 
C6034 VCC.n2198 VSS 1.54e-19 
C6035 VCC.n2199 VSS 1.65e-20 
C6036 VCC.t3 VSS 1.56e-19 
C6037 VCC.n2200 VSS 7.62e-19 
C6038 VCC.n2201 VSS 1.23e-20 
C6039 VCC.n2202 VSS 2.47e-20 
C6040 VCC.n2203 VSS 4.73e-20 
C6041 VCC.n2204 VSS 6.59e-20 
C6042 VCC.n2205 VSS 5.15e-20 
C6043 VCC.n2206 VSS 2.47e-20 
C6044 VCC.n2207 VSS 7.41e-20 
C6045 VCC.n2208 VSS 9.47e-20 
C6046 VCC.n2209 VSS 1.32e-19 
C6047 VCC.n2210 VSS 7.71e-19 
C6048 VCC.n2211 VSS 9.83e-19 
C6049 VCC.n2212 VSS 2.36e-19 
C6050 VCC.n2213 VSS 3.21e-19 
C6051 VCC.n2214 VSS 2.61e-19 
C6052 VCC.n2215 VSS 0.00189f 
C6053 VCC.n2216 VSS 0.00276f 
C6054 VCC.n2217 VSS 5.76e-20 
C6055 VCC.n2218 VSS 2.88e-20 
C6056 VCC.n2219 VSS 3.5e-20 
C6057 VCC.n2220 VSS 9.83e-19 
C6058 VCC.n2221 VSS 9.47e-20 
C6059 VCC.n2222 VSS 1.17e-19 
C6060 VCC.n2223 VSS 2.06e-19 
C6061 VCC.n2224 VSS 1.36e-19 
C6062 VCC.n2225 VSS 1.01e-19 
C6063 VCC.n2226 VSS 3.5e-20 
C6064 VCC.n2227 VSS 3.09e-20 
C6065 VCC.n2228 VSS 3.29e-20 
C6066 VCC.n2229 VSS 3.29e-20 
C6067 VCC.n2230 VSS 4.73e-20 
C6068 VCC.n2231 VSS 1.44e-20 
C6069 VCC.n2232 VSS 3.5e-20 
C6070 VCC.n2233 VSS 7.41e-20 
C6071 VCC.n2234 VSS 2.47e-20 
C6072 VCC.t46 VSS 1.56e-19 
C6073 VCC.n2235 VSS 5.76e-20 
C6074 VCC.n2236 VSS 2.06e-20 
C6075 VCC.n2237 VSS 5.76e-20 
C6076 VCC.n2238 VSS 3.7e-20 
C6077 VCC.n2239 VSS 4.32e-20 
C6078 VCC.n2240 VSS 2.68e-20 
C6079 VCC.n2241 VSS 3.91e-20 
C6080 VCC.n2242 VSS 6.38e-20 
C6081 VCC.n2243 VSS 1.85e-20 
C6082 VCC.n2244 VSS 3.5e-20 
C6083 VCC.n2245 VSS 3.09e-20 
C6084 VCC.n2246 VSS 3.7e-20 
C6085 VCC.n2247 VSS 3.09e-20 
C6086 VCC.n2248 VSS 2.26e-20 
C6087 VCC.n2249 VSS 1.05e-19 
C6088 VCC.n2250 VSS 3.5e-20 
C6089 VCC.n2251 VSS 3.5e-20 
C6090 VCC.n2252 VSS 8.42e-19 
C6091 VCC.n2253 VSS 2.18e-19 
C6092 VCC.n2254 VSS 1.4e-19 
C6093 VCC.n2255 VSS 4.32e-20 
C6094 VCC.n2256 VSS 7.82e-20 
C6095 VCC.n2257 VSS 5.76e-20 
C6096 VCC.n2258 VSS 2.68e-20 
C6097 VCC.n2259 VSS 4.32e-20 
C6098 VCC.n2260 VSS 3.91e-20 
C6099 VCC.n2261 VSS 3.7e-20 
C6100 VCC.n2262 VSS 3.7e-20 
C6101 VCC.n2263 VSS 5.76e-20 
C6102 VCC.n2264 VSS 4.73e-20 
C6103 VCC.n2265 VSS 3.5e-20 
C6104 VCC.t188 VSS 1.56e-19 
C6105 VCC.n2266 VSS 7.97e-19 
C6106 VCC.n2267 VSS 3.09e-20 
C6107 VCC.n2268 VSS 1.01e-19 
C6108 VCC.n2269 VSS 3.5e-20 
C6109 VCC.n2270 VSS 1.36e-19 
C6110 VCC.n2271 VSS 3.5e-20 
C6111 VCC.n2272 VSS 3.33e-19 
C6112 VCC.n2273 VSS 1.17e-19 
C6113 VCC.n2274 VSS 1.09e-19 
C6114 VCC.n2275 VSS 3.5e-20 
C6115 VCC.n2276 VSS 4.73e-20 
C6116 VCC.n2277 VSS 5.56e-20 
C6117 VCC.n2278 VSS 2.88e-20 
C6118 VCC.n2279 VSS 2.26e-20 
C6119 VCC.n2280 VSS 5.76e-20 
C6120 VCC.n2281 VSS 2.68e-20 
C6121 VCC.n2282 VSS 2.68e-20 
C6122 VCC.n2283 VSS 1.9e-19 
C6123 VCC.n2284 VSS 5.76e-20 
C6124 VCC.n2285 VSS 2.68e-20 
C6125 VCC.n2286 VSS 2.68e-20 
C6126 VCC.n2287 VSS 2.68e-20 
C6127 VCC.n2288 VSS 5.76e-20 
C6128 VCC.n2289 VSS 2.26e-20 
C6129 VCC.n2290 VSS 3.09e-20 
C6130 VCC.n2291 VSS 2.26e-20 
C6131 VCC.n2292 VSS 5.15e-20 
C6132 VCC.n2293 VSS 4.73e-20 
C6133 VCC.n2294 VSS 3.7e-20 
C6134 VCC.n2295 VSS 3.5e-20 
C6135 VCC.n2296 VSS 7.41e-20 
C6136 VCC.n2297 VSS 1.91e-19 
C6137 VCC.n2298 VSS 9.88e-20 
C6138 VCC.n2299 VSS 3e-20 
C6139 VCC.n2300 VSS 5.12e-19 
C6140 VCC.n2301 VSS 1.18e-19 
C6141 VCC.n2302 VSS 3.5e-20 
C6142 VCC.n2303 VSS 3.5e-20 
C6143 VCC.n2304 VSS 5.15e-20 
C6144 VCC.n2305 VSS 4.32e-20 
C6145 VCC.n2306 VSS 2.68e-20 
C6146 VCC.n2307 VSS 3.91e-20 
C6147 VCC.n2308 VSS 1.44e-20 
C6148 VCC.n2309 VSS 3.5e-20 
C6149 VCC.n2310 VSS 3e-20 
C6150 VCC.n2311 VSS 7.95e-19 
C6151 VCC.n2312 VSS 1.83e-19 
C6152 VCC.n2313 VSS 2.88e-20 
C6153 VCC.n2314 VSS 2.68e-20 
C6154 VCC.n2315 VSS 2.68e-20 
C6155 VCC.n2316 VSS 2.68e-20 
C6156 VCC.n2317 VSS 4.53e-20 
C6157 VCC.n2318 VSS 3.7e-20 
C6158 VCC.n2319 VSS 7.82e-20 
C6159 VCC.n2320 VSS 1.17e-19 
C6160 VCC.n2321 VSS 3.91e-20 
C6161 VCC.n2322 VSS 1.65e-20 
C6162 VCC.n2323 VSS 2.68e-20 
C6163 VCC.n2324 VSS 3.5e-20 
C6164 VCC.n2325 VSS 3e-20 
C6165 VCC.n2326 VSS 5.12e-19 
C6166 VCC.n2327 VSS 1.18e-19 
C6167 VCC.n2328 VSS 3.5e-20 
C6168 VCC.n2329 VSS 3.5e-20 
C6169 VCC.t196 VSS 1.55e-19 
C6170 VCC.n2330 VSS 7.57e-19 
C6171 VCC.n2331 VSS 4.73e-20 
C6172 VCC.n2332 VSS 1.54e-19 
C6173 VCC.n2333 VSS 2.88e-20 
C6174 VCC.n2334 VSS 2.88e-20 
C6175 VCC.n2335 VSS 3.5e-20 
C6176 VCC.n2336 VSS 5.76e-20 
C6177 VCC.n2337 VSS 9.88e-20 
C6178 VCC.n2338 VSS 1.3e-19 
C6179 VCC.n2339 VSS 3e-20 
C6180 VCC.t194 VSS 0.005f 
C6181 VCC.t229 VSS 0.00453f 
C6182 VCC.n2340 VSS 0.00229f 
C6183 VCC.n2341 VSS 1.91e-19 
C6184 VCC.n2342 VSS 3.5e-20 
C6185 VCC.n2343 VSS 3.14e-19 
C6186 VCC.n2344 VSS 3.5e-20 
C6187 VCC.n2345 VSS 2.47e-20 
C6188 VCC.n2346 VSS 5.76e-20 
C6189 VCC.n2347 VSS 2.47e-20 
C6190 VCC.n2348 VSS 8.23e-21 
C6191 VCC.n2349 VSS 2.88e-20 
C6192 VCC.n2350 VSS 5.76e-20 
C6193 VCC.n2351 VSS 2.47e-20 
C6194 VCC.n2352 VSS 2.88e-20 
C6195 VCC.n2353 VSS 2.47e-20 
C6196 VCC.n2354 VSS 5.15e-20 
C6197 VCC.n2355 VSS 4.73e-20 
C6198 VCC.n2356 VSS 3.7e-20 
C6199 VCC.n2357 VSS 3.5e-20 
C6200 VCC.n2358 VSS 7.41e-20 
C6201 VCC.t32 VSS 6.42e-19 
C6202 VCC.n2359 VSS 3e-20 
C6203 VCC.n2360 VSS 5.97e-20 
C6204 VCC.n2361 VSS 4.13e-19 
C6205 VCC.n2362 VSS 9.53e-20 
C6206 VCC.n2363 VSS 3.5e-20 
C6207 VCC.n2364 VSS 3.5e-20 
C6208 VCC.n2365 VSS 5.35e-20 
C6209 VCC.n2366 VSS 4.32e-20 
C6210 VCC.n2367 VSS 2.68e-20 
C6211 VCC.n2368 VSS 3.7e-20 
C6212 VCC.n2369 VSS 1.65e-20 
C6213 VCC.n2370 VSS 4.53e-20 
C6214 VCC.n2371 VSS 1.2e-19 
C6215 VCC.n2372 VSS 5.2e-19 
C6216 VCC.n2373 VSS 1.2e-19 
C6217 VCC.n2374 VSS 6.38e-20 
C6218 VCC.n2375 VSS 2.47e-20 
C6219 VCC.n2376 VSS 4.53e-20 
C6220 VCC.n2377 VSS 3.5e-20 
C6221 VCC.n2378 VSS 3.5e-20 
C6222 VCC.n2379 VSS 2.68e-20 
C6223 VCC.n2380 VSS 2.68e-20 
C6224 VCC.n2381 VSS 2.47e-20 
C6225 VCC.n2382 VSS 4.53e-20 
C6226 VCC.n2383 VSS 2.68e-20 
C6227 VCC.n2384 VSS 4.32e-20 
C6228 VCC.n2385 VSS 2.68e-20 
C6229 VCC.n2386 VSS 3.91e-20 
C6230 VCC.n2387 VSS 2.88e-20 
C6231 VCC.n2388 VSS 4.73e-20 
C6232 VCC.n2389 VSS 3.7e-20 
C6233 VCC.n2390 VSS 3.7e-20 
C6234 VCC.n2391 VSS 3.5e-20 
C6235 VCC.n2392 VSS 5.76e-20 
C6236 VCC.n2393 VSS 4.73e-20 
C6237 VCC.n2394 VSS 3.09e-20 
C6238 VCC.n2395 VSS 3.5e-20 
C6239 VCC.n2396 VSS 3.5e-20 
C6240 VCC.n2397 VSS 3.5e-20 
C6241 VCC.n2398 VSS 1.18e-19 
C6242 VCC.n2399 VSS 3e-20 
C6243 VCC.n2400 VSS 1.15e-19 
C6244 VCC.n2401 VSS 9.88e-20 
C6245 VCC.n2402 VSS 5.76e-20 
C6246 VCC.n2403 VSS 3.5e-20 
C6247 VCC.n2404 VSS 3.09e-20 
C6248 VCC.n2405 VSS 3.09e-20 
C6249 VCC.n2406 VSS 2.26e-20 
C6250 VCC.n2407 VSS 5.76e-20 
C6251 VCC.n2408 VSS 2.68e-20 
C6252 VCC.n2409 VSS 2.68e-20 
C6253 VCC.n2410 VSS 0.00185f 
C6254 VCC.n2411 VSS 2.72e-19 
C6255 VCC.n2412 VSS 2.26e-20 
C6256 VCC.n2413 VSS 1.87e-19 
C6257 VCC.n2414 VSS 3.5e-20 
C6258 VCC.n2415 VSS 2.68e-20 
C6259 VCC.n2416 VSS 5.97e-20 
C6260 VCC.n2417 VSS 4.73e-20 
C6261 VCC.n2418 VSS 4.73e-20 
C6262 VCC.n2419 VSS 5.15e-20 
C6263 VCC.n2420 VSS 7.41e-20 
C6264 VCC.n2421 VSS 3.7e-20 
C6265 VCC.n2422 VSS 2.26e-20 
C6266 VCC.n2423 VSS 6.38e-20 
C6267 VCC.n2424 VSS 4.73e-20 
C6268 VCC.n2425 VSS 3.29e-20 
C6269 VCC.n2426 VSS 3.5e-20 
C6270 VCC.n2427 VSS 3e-20 
C6271 VCC.t228 VSS 0.005f 
C6272 VCC.t313 VSS 0.00453f 
C6273 VCC.n2428 VSS 0.00228f 
C6274 VCC.n2429 VSS 1.3e-19 
C6275 VCC.t226 VSS 4.05e-19 
C6276 VCC.n2430 VSS 4.05e-19 
C6277 VCC.n2431 VSS 1.15e-19 
C6278 VCC.n2432 VSS 3.36e-19 
C6279 VCC.n2433 VSS 6.17e-21 
C6280 VCC.n2434 VSS 3.12e-19 
C6281 VCC.n2435 VSS 1.65e-20 
C6282 VCC.n2436 VSS 1.54e-19 
C6283 VCC.n2437 VSS 1.54e-19 
C6284 VCC.n2438 VSS 1.65e-20 
C6285 VCC.n2439 VSS 1.03e-20 
C6286 VCC.n2440 VSS 3.5e-20 
C6287 VCC.n2441 VSS 2.26e-20 
C6288 VCC.n2442 VSS 4.73e-20 
C6289 VCC.n2443 VSS 3.5e-20 
C6290 VCC.n2444 VSS 3e-20 
C6291 VCC.n2445 VSS 1.3e-19 
C6292 VCC.n2446 VSS 5.12e-19 
C6293 VCC.n2447 VSS 1.3e-19 
C6294 VCC.n2448 VSS 4.13e-19 
C6295 VCC.n2449 VSS 9.53e-20 
C6296 VCC.n2450 VSS 5.76e-20 
C6297 VCC.n2451 VSS 7.41e-20 
C6298 VCC.n2452 VSS 5.56e-20 
C6299 VCC.t227 VSS 1.55e-19 
C6300 VCC.n2453 VSS 3.91e-20 
C6301 VCC.n2454 VSS 3.91e-20 
C6302 VCC.n2455 VSS 1.85e-20 
C6303 VCC.n2456 VSS 7.55e-19 
C6304 VCC.n2457 VSS 4.94e-20 
C6305 VCC.n2458 VSS 5.15e-20 
C6306 VCC.n2459 VSS 7.2e-20 
C6307 VCC.n2460 VSS 1.38e-19 
C6308 VCC.n2461 VSS 1.17e-19 
C6309 VCC.n2462 VSS 4.32e-20 
C6310 VCC.n2463 VSS 2.88e-20 
C6311 VCC.n2464 VSS 2.68e-20 
C6312 VCC.n2465 VSS 3.5e-20 
C6313 VCC.n2466 VSS 3.5e-20 
C6314 VCC.n2467 VSS 2.88e-20 
C6315 VCC.n2468 VSS 2.68e-20 
C6316 VCC.n2469 VSS 2.68e-20 
C6317 VCC.n2470 VSS 2.68e-20 
C6318 VCC.n2471 VSS 4.12e-20 
C6319 VCC.n2472 VSS 4.12e-20 
C6320 VCC.n2473 VSS 3.91e-20 
C6321 VCC.n2474 VSS 4.53e-20 
C6322 VCC.n2475 VSS 4.53e-20 
C6323 VCC.n2476 VSS 1.05e-19 
C6324 VCC.n2477 VSS 1.05e-19 
C6325 VCC.n2478 VSS 4.32e-20 
C6326 VCC.n2479 VSS 3.7e-20 
C6327 VCC.n2480 VSS 2.68e-20 
C6328 VCC.n2481 VSS 2.68e-20 
C6329 VCC.n2482 VSS 6.79e-20 
C6330 VCC.n2483 VSS 9.26e-20 
C6331 VCC.n2484 VSS 1.83e-19 
C6332 VCC.n2485 VSS 7.95e-19 
C6333 VCC.n2486 VSS 5.2e-19 
C6334 VCC.n2487 VSS 1.3e-19 
C6335 VCC.n2488 VSS 3e-20 
C6336 VCC.n2489 VSS 3.5e-20 
C6337 VCC.n2490 VSS 5.97e-20 
C6338 VCC.n2491 VSS 7.41e-20 
C6339 VCC.n2492 VSS 5.15e-20 
C6340 VCC.n2493 VSS 5.15e-20 
C6341 VCC.n2494 VSS 3.09e-20 
C6342 VCC.n2495 VSS 3.09e-20 
C6343 VCC.n2496 VSS 3.7e-20 
C6344 VCC.n2497 VSS 2.68e-20 
C6345 VCC.n2498 VSS 3.91e-20 
C6346 VCC.n2499 VSS 1.17e-19 
C6347 VCC.n2500 VSS 1.38e-19 
C6348 VCC.n2501 VSS 7e-20 
C6349 VCC.n2502 VSS 4.73e-20 
C6350 VCC.n2503 VSS 3.5e-20 
C6351 VCC.n2504 VSS 3.5e-20 
C6352 VCC.n2505 VSS 3.5e-20 
C6353 VCC.n2506 VSS 4.53e-20 
C6354 VCC.n2507 VSS 1.18e-19 
C6355 VCC.n2508 VSS 5.12e-19 
C6356 VCC.n2509 VSS 1.3e-19 
C6357 VCC.n2510 VSS 1.61e-19 
C6358 VCC.n2511 VSS 9.9e-20 
C6359 VCC.n2512 VSS 0.00243f 
C6360 VCC.n2513 VSS 2.26e-20 
C6361 VCC.n2514 VSS 4.13e-19 
C6362 VCC.n2515 VSS 3.5e-20 
C6363 VCC.n2516 VSS 3.5e-20 
C6364 VCC.n2517 VSS 2.47e-20 
C6365 VCC.n2518 VSS 2.06e-20 
C6366 VCC.n2519 VSS 6.17e-20 
C6367 VCC.n2520 VSS 6.17e-20 
C6368 VCC.n2521 VSS 4.73e-20 
C6369 VCC.n2522 VSS 4.73e-20 
C6370 VCC.n2523 VSS 2.88e-20 
C6371 VCC.n2524 VSS 1.44e-20 
C6372 VCC.n2525 VSS 1.65e-20 
C6373 VCC.n2526 VSS 1.54e-19 
C6374 VCC.n2527 VSS 1.54e-19 
C6375 VCC.n2528 VSS 1.65e-20 
C6376 VCC.n2529 VSS 3.09e-20 
C6377 VCC.t33 VSS 1.55e-19 
C6378 VCC.n2530 VSS 0.00102f 
C6379 VCC.n2531 VSS 2.73e-19 
C6380 VCC.n2532 VSS 0.00136f 
C6381 VCC.n2533 VSS 2.73e-19 
C6382 VCC.n2534 VSS 0.00181f 
C6383 VCC.n2535 VSS 5.76e-20 
C6384 VCC.n2536 VSS 1.54e-19 
C6385 VCC.n2537 VSS 1.65e-20 
C6386 VCC.n2538 VSS 6.17e-20 
C6387 VCC.n2539 VSS 2.47e-20 
C6388 VCC.n2540 VSS 4.73e-20 
C6389 VCC.n2541 VSS 4.73e-20 
C6390 VCC.n2542 VSS 5.15e-20 
C6391 VCC.n2543 VSS 3.5e-20 
C6392 VCC.n2544 VSS 7.41e-20 
C6393 VCC.n2545 VSS 3.7e-20 
C6394 VCC.n2546 VSS 2.26e-20 
C6395 VCC.n2547 VSS 6.17e-20 
C6396 VCC.n2548 VSS 4.73e-20 
C6397 VCC.n2549 VSS 2.88e-20 
C6398 VCC.n2550 VSS 2.88e-20 
C6399 VCC.n2551 VSS 3.4e-19 
C6400 VCC.n2552 VSS 1.15e-19 
C6401 VCC.n2553 VSS 3.98e-19 
C6402 VCC.t195 VSS 4.05e-19 
C6403 VCC.n2554 VSS 1.22e-19 
C6404 VCC.n2555 VSS 1.3e-19 
C6405 VCC.n2556 VSS 3e-20 
C6406 VCC.n2557 VSS 3.5e-20 
C6407 VCC.n2558 VSS 3.5e-20 
C6408 VCC.n2559 VSS 4.73e-20 
C6409 VCC.n2560 VSS 2.47e-20 
C6410 VCC.n2561 VSS 1.23e-20 
C6411 VCC.n2562 VSS 1.65e-20 
C6412 VCC.n2563 VSS 2.47e-20 
C6413 VCC.n2564 VSS 5.76e-20 
C6414 VCC.n2565 VSS 1.38e-19 
C6415 VCC.n2566 VSS 7e-20 
C6416 VCC.n2567 VSS 3.7e-20 
C6417 VCC.n2568 VSS 2.47e-20 
C6418 VCC.n2569 VSS 3.7e-20 
C6419 VCC.n2570 VSS 1.85e-20 
C6420 VCC.n2571 VSS 3.09e-20 
C6421 VCC.n2572 VSS 5.35e-20 
C6422 VCC.n2573 VSS 4.73e-20 
C6423 VCC.n2574 VSS 5.35e-20 
C6424 VCC.n2575 VSS 7.41e-20 
C6425 VCC.n2576 VSS 5.76e-20 
C6426 VCC.n2577 VSS 9.53e-20 
C6427 VCC.n2578 VSS 4.13e-19 
C6428 VCC.n2579 VSS 1.3e-19 
C6429 VCC.n2580 VSS 5.2e-19 
C6430 VCC.n2581 VSS 1.2e-19 
C6431 VCC.n2582 VSS 4.73e-20 
C6432 VCC.n2583 VSS 2.68e-20 
C6433 VCC.n2584 VSS 3.5e-20 
C6434 VCC.n2585 VSS 3.5e-20 
C6435 VCC.n2586 VSS 2.68e-20 
C6436 VCC.n2587 VSS 2.68e-20 
C6437 VCC.n2588 VSS 4.32e-20 
C6438 VCC.n2589 VSS 4.32e-20 
C6439 VCC.n2590 VSS 4.32e-20 
C6440 VCC.n2591 VSS 2.88e-20 
C6441 VCC.n2592 VSS 3.5e-20 
C6442 VCC.n2593 VSS 2.68e-20 
C6443 VCC.n2594 VSS 7.82e-20 
C6444 VCC.n2595 VSS 4.73e-20 
C6445 VCC.n2596 VSS 4.73e-20 
C6446 VCC.n2597 VSS 1.05e-19 
C6447 VCC.n2598 VSS 1.05e-19 
C6448 VCC.n2599 VSS 4.53e-20 
C6449 VCC.n2600 VSS 2.68e-20 
C6450 VCC.n2601 VSS 2.68e-20 
C6451 VCC.n2602 VSS 6.59e-20 
C6452 VCC.n2603 VSS 9.26e-20 
C6453 VCC.n2604 VSS 6.59e-20 
C6454 VCC.n2605 VSS 2.47e-20 
C6455 VCC.n2606 VSS 2.47e-20 
C6456 VCC.n2607 VSS 2.88e-20 
C6457 VCC.n2608 VSS 3.5e-20 
C6458 VCC.n2609 VSS 3.5e-20 
C6459 VCC.n2610 VSS 4.53e-20 
C6460 VCC.n2611 VSS 1.2e-19 
C6461 VCC.n2612 VSS 5.2e-19 
C6462 VCC.n2613 VSS 1.3e-19 
C6463 VCC.n2614 VSS 4.13e-19 
C6464 VCC.n2615 VSS 9.53e-20 
C6465 VCC.n2616 VSS 5.97e-20 
C6466 VCC.n2617 VSS 7.41e-20 
C6467 VCC.n2618 VSS 5.35e-20 
C6468 VCC.n2619 VSS 5.15e-20 
C6469 VCC.n2620 VSS 3.09e-20 
C6470 VCC.n2621 VSS 3.09e-20 
C6471 VCC.n2622 VSS 3.91e-20 
C6472 VCC.n2623 VSS 2.47e-20 
C6473 VCC.n2624 VSS 3.7e-20 
C6474 VCC.n2625 VSS 1.17e-19 
C6475 VCC.n2626 VSS 1.38e-19 
C6476 VCC.n2627 VSS 7.2e-20 
C6477 VCC.n2628 VSS 4.73e-20 
C6478 VCC.n2629 VSS 3.5e-20 
C6479 VCC.n2630 VSS 3.5e-20 
C6480 VCC.n2631 VSS 4.53e-20 
C6481 VCC.n2632 VSS 5.97e-20 
C6482 VCC.n2633 VSS 3.5e-20 
C6483 VCC.n2634 VSS 3e-20 
C6484 VCC.n2635 VSS 1.3e-19 
C6485 VCC.n2636 VSS 1.53e-19 
C6486 VCC.t143 VSS 4.05e-19 
C6487 VCC.n2637 VSS 1.35e-19 
C6488 VCC.t187 VSS 4.21e-19 
C6489 VCC.n2638 VSS 2.06e-19 
C6490 VCC.n2639 VSS 1.32e-19 
C6491 VCC.n2640 VSS 9.67e-20 
C6492 VCC.n2641 VSS 3.35e-20 
C6493 VCC.n2642 VSS 3.5e-20 
C6494 VCC.n2643 VSS 2.36e-19 
C6495 VCC.n2644 VSS 0.0023f 
C6496 VCC.t190 VSS 0.0031f 
C6497 VCC.t197 VSS 0.00366f 
C6498 VCC.t189 VSS 0.00365f 
C6499 VCC.t200 VSS 0.00386f 
C6500 VCC.n2645 VSS 0.00569f 
C6501 VCC.n2646 VSS 1.3e-19 
C6502 VCC.n2647 VSS 3.67e-19 
C6503 VCC.n2648 VSS 1.15e-19 
C6504 VCC.n2649 VSS 3.38e-19 
C6505 VCC.n2650 VSS 3.5e-20 
C6506 VCC.n2651 VSS 3.5e-20 
C6507 VCC.n2652 VSS 2.68e-20 
C6508 VCC.n2653 VSS 2.06e-20 
C6509 VCC.n2654 VSS 6.38e-20 
C6510 VCC.n2655 VSS 5.97e-20 
C6511 VCC.n2656 VSS 4.73e-20 
C6512 VCC.n2657 VSS 4.73e-20 
C6513 VCC.n2658 VSS 3.09e-20 
C6514 VCC.n2659 VSS 1.23e-20 
C6515 VCC.n2660 VSS 1.65e-20 
C6516 VCC.n2661 VSS 1.54e-19 
C6517 VCC.n2662 VSS 1.54e-19 
C6518 VCC.n2663 VSS 1.65e-20 
C6519 VCC.n2664 VSS 3.29e-20 
C6520 VCC.t144 VSS 1.67e-19 
C6521 VCC.n2665 VSS 0.00101f 
C6522 VCC.n2666 VSS 2.71e-19 
C6523 VCC.n2667 VSS 7.46e-19 
C6524 VCC.n2668 VSS 0.00333f 
C6525 VCC.n2669 VSS 2.46e-19 
C6526 VCC.n2670 VSS 3.02e-19 
C6527 VCC.n2671 VSS 3.7e-20 
C6528 VCC.n2672 VSS 5.15e-20 
C6529 VCC.n2673 VSS 5.97e-20 
C6530 VCC.n2674 VSS 6.38e-20 
C6531 VCC.n2675 VSS 4.73e-20 
C6532 VCC.n2676 VSS 4.73e-20 
C6533 VCC.n2677 VSS 2.68e-20 
C6534 VCC.n2678 VSS 3.29e-20 
C6535 VCC.n2679 VSS 1.65e-20 
C6536 VCC.n2680 VSS 1.54e-19 
C6537 VCC.n2681 VSS 1.54e-19 
C6538 VCC.n2682 VSS 1.65e-20 
C6539 VCC.n2683 VSS 3.09e-20 
C6540 VCC.n2684 VSS 3.09e-20 
C6541 VCC.n2685 VSS 4.73e-20 
C6542 VCC.n2686 VSS 4.32e-20 
C6543 VCC.n2687 VSS 3.5e-20 
C6544 VCC.n2688 VSS 3.5e-20 
C6545 VCC.n2689 VSS 1.35e-19 
C6546 VCC.n2690 VSS 5.24e-19 
C6547 VCC.n2691 VSS 1.4e-19 
C6548 VCC.n2692 VSS 5.4e-19 
C6549 VCC.n2693 VSS 1.35e-19 
C6550 VCC.n2694 VSS 4.37e-19 
C6551 VCC.n2695 VSS 1.13e-19 
C6552 VCC.n2696 VSS 8.23e-21 
C6553 VCC.n2697 VSS 1.65e-20 
C6554 VCC.n2698 VSS 3.5e-20 
C6555 VCC.n2699 VSS 3.91e-20 
C6556 VCC.n2700 VSS 3.09e-20 
C6557 VCC.n2701 VSS 1.85e-20 
C6558 VCC.n2702 VSS 3.5e-20 
C6559 VCC.n2703 VSS 1.05e-19 
C6560 VCC.n2704 VSS 2.06e-20 
C6561 VCC.n2705 VSS 2.26e-20 
C6562 VCC.n2706 VSS 3.7e-20 
C6563 VCC.n2707 VSS 5.15e-20 
C6564 VCC.n2708 VSS 1.38e-19 
C6565 VCC.n2709 VSS 1.17e-19 
C6566 VCC.n2710 VSS 4.32e-20 
C6567 VCC.n2711 VSS 2.88e-20 
C6568 VCC.n2712 VSS 2.68e-20 
C6569 VCC.n2713 VSS 6.59e-20 
C6570 VCC.n2714 VSS 5.56e-20 
C6571 VCC.n2715 VSS 2.68e-20 
C6572 VCC.n2716 VSS 4.32e-20 
C6573 VCC.n2717 VSS 1.05e-19 
C6574 VCC.n2718 VSS 3.09e-20 
C6575 VCC.n2719 VSS 3.7e-20 
C6576 VCC.n2720 VSS 4.32e-20 
C6577 VCC.n2721 VSS 1.05e-19 
C6578 VCC.n2722 VSS 4.53e-20 
C6579 VCC.n2723 VSS 4.53e-20 
C6580 VCC.n2724 VSS 7.82e-20 
C6581 VCC.n2725 VSS 2.18e-19 
C6582 VCC.n2726 VSS 1.4e-19 
C6583 VCC.n2727 VSS 1.4e-19 
C6584 VCC.n2728 VSS 5.4e-19 
C6585 VCC.n2729 VSS 1.35e-19 
C6586 VCC.t45 VSS 4.21e-19 
C6587 VCC.n2730 VSS 3.33e-19 
C6588 VCC.n2731 VSS 1.13e-19 
C6589 VCC.n2732 VSS 8.23e-21 
C6590 VCC.n2733 VSS 1.65e-20 
C6591 VCC.n2734 VSS 3.5e-20 
C6592 VCC.n2735 VSS 3.5e-20 
C6593 VCC.n2736 VSS 3.5e-20 
C6594 VCC.n2737 VSS 1.17e-19 
C6595 VCC.n2738 VSS 1.38e-19 
C6596 VCC.n2739 VSS 5.15e-20 
C6597 VCC.n2740 VSS 4.73e-20 
C6598 VCC.n2741 VSS 7.2e-20 
C6599 VCC.n2742 VSS 2.68e-20 
C6600 VCC.n2743 VSS 1.65e-20 
C6601 VCC.n2744 VSS 1.54e-19 
C6602 VCC.n2745 VSS 1.54e-19 
C6603 VCC.n2746 VSS 1.65e-20 
C6604 VCC.n2747 VSS 2.47e-20 
C6605 VCC.n2748 VSS 1.23e-20 
C6606 VCC.n2749 VSS 7.62e-19 
C6607 VCC.n2750 VSS 4.12e-20 
C6608 VCC.n2751 VSS 5.15e-20 
C6609 VCC.n2752 VSS 6.59e-20 
C6610 VCC.n2753 VSS 5.76e-20 
C6611 VCC.n2754 VSS 4.73e-20 
C6612 VCC.n2755 VSS 2.26e-20 
C6613 VCC.n2756 VSS 2.68e-20 
C6614 VCC.n2757 VSS 1.03e-20 
C6615 VCC.n2758 VSS 3.5e-20 
C6616 VCC.n2759 VSS 3.5e-20 
C6617 VCC.n2760 VSS 1.35e-19 
C6618 VCC.n2761 VSS 4.53e-19 
C6619 VCC.n2762 VSS 7.71e-19 
C6620 VCC.n2763 VSS 1.32e-19 
C6621 VCC.n2764 VSS 3.5e-20 
C6622 VCC.n2765 VSS 3.42e-20 
C6623 VCC.n2766 VSS 2.36e-19 
C6624 VCC.n2767 VSS 3.21e-19 
C6625 VCC.n2768 VSS 2.61e-19 
C6626 VCC.n2769 VSS 0.00189f 
C6627 VCC.n2770 VSS 2.68e-19 
C6628 VCC.n2771 VSS 3.52e-19 
C6629 VCC.n2772 VSS 5.76e-20 
C6630 VCC.n2773 VSS 2.88e-20 
C6631 VCC.n2774 VSS 3.5e-20 
C6632 VCC.n2775 VSS 3.42e-20 
C6633 VCC.n2776 VSS 3.5e-20 
C6634 VCC.n2777 VSS 4.53e-19 
C6635 VCC.n2778 VSS 1.17e-19 
C6636 VCC.n2779 VSS 3.5e-20 
C6637 VCC.n2780 VSS 1.44e-20 
C6638 VCC.n2781 VSS 4.12e-20 
C6639 VCC.n2782 VSS 5.76e-20 
C6640 VCC.n2783 VSS 5.76e-20 
C6641 VCC.n2784 VSS 2.06e-20 
C6642 VCC.n2785 VSS 3.29e-20 
C6643 VCC.n2786 VSS 7.2e-20 
C6644 VCC.n2787 VSS 3.29e-20 
C6645 VCC.n2788 VSS 4.73e-20 
C6646 VCC.n2789 VSS 2.26e-20 
C6647 VCC.n2790 VSS 1.01e-19 
C6648 VCC.n2791 VSS 1.36e-19 
C6649 VCC.n2792 VSS 1.35e-19 
C6650 VCC.n2793 VSS 3.5e-20 
C6651 VCC.n2794 VSS 3.5e-20 
C6652 VCC.n2795 VSS 3.5e-20 
C6653 VCC.n2796 VSS 3.5e-20 
C6654 VCC.n2797 VSS 3.09e-20 
C6655 VCC.n2798 VSS 3.91e-20 
C6656 VCC.n2799 VSS 4.73e-20 
C6657 VCC.n2800 VSS 4.32e-20 
C6658 VCC.n2801 VSS 2.68e-20 
C6659 VCC.n2802 VSS 4.53e-20 
C6660 VCC.n2803 VSS 4.53e-20 
C6661 VCC.n2804 VSS 3.09e-20 
C6662 VCC.n2805 VSS 4.32e-20 
C6663 VCC.n2806 VSS 2.68e-20 
C6664 VCC.n2807 VSS 7.82e-20 
C6665 VCC.n2808 VSS 5.56e-20 
C6666 VCC.n2809 VSS 1.4e-19 
C6667 VCC.n2810 VSS 2.18e-19 
C6668 VCC.n2811 VSS 1.35e-19 
C6669 VCC.n2812 VSS 1.13e-19 
C6670 VCC.n2813 VSS 3.5e-20 
C6671 VCC.n2814 VSS 1.85e-20 
C6672 VCC.n2815 VSS 3.7e-20 
C6673 VCC.n2816 VSS 3.09e-20 
C6674 VCC.n2817 VSS 6.59e-20 
C6675 VCC.n2818 VSS 2.68e-20 
C6676 VCC.n2819 VSS 5.76e-20 
C6677 VCC.n2820 VSS 4.73e-20 
C6678 VCC.n2821 VSS 3.5e-20 
C6679 VCC.t96 VSS 1.56e-19 
C6680 VCC.n2822 VSS 7.97e-19 
C6681 VCC.n2823 VSS 3.09e-20 
C6682 VCC.n2824 VSS 3.5e-20 
C6683 VCC.n2825 VSS 3.5e-20 
C6684 VCC.t95 VSS 4.21e-19 
C6685 VCC.n2826 VSS 1.32e-19 
C6686 VCC.n2827 VSS 1.09e-19 
C6687 VCC.n2828 VSS 3.5e-20 
C6688 VCC.n2829 VSS 3.09e-20 
C6689 VCC.n2830 VSS 5.97e-20 
C6690 VCC.n2831 VSS 2.26e-20 
C6691 VCC.n2832 VSS 5.76e-20 
C6692 VCC.n2833 VSS 2.68e-20 
C6693 VCC.n2834 VSS 2.68e-20 
C6694 VCC.n2835 VSS 1.9e-19 
C6695 VCC.n2836 VSS 5.76e-20 
C6696 VCC.n2837 VSS 2.68e-20 
C6697 VCC.n2838 VSS 2.68e-20 
C6698 VCC.n2839 VSS 2.68e-20 
C6699 VCC.n2840 VSS 5.76e-20 
C6700 VCC.n2841 VSS 2.26e-20 
C6701 VCC.n2842 VSS 3.09e-20 
C6702 VCC.n2843 VSS 2.26e-20 
C6703 VCC.n2844 VSS 5.15e-20 
C6704 VCC.n2845 VSS 4.73e-20 
C6705 VCC.n2846 VSS 3.7e-20 
C6706 VCC.n2847 VSS 3.5e-20 
C6707 VCC.n2848 VSS 7.41e-20 
C6708 VCC.n2849 VSS 1.91e-19 
C6709 VCC.n2850 VSS 9.88e-20 
C6710 VCC.n2851 VSS 3e-20 
C6711 VCC.n2852 VSS 5.12e-19 
C6712 VCC.n2853 VSS 1.18e-19 
C6713 VCC.n2854 VSS 3.5e-20 
C6714 VCC.n2855 VSS 3.5e-20 
C6715 VCC.n2856 VSS 5.15e-20 
C6716 VCC.n2857 VSS 4.32e-20 
C6717 VCC.n2858 VSS 2.68e-20 
C6718 VCC.n2859 VSS 3.91e-20 
C6719 VCC.n2860 VSS 1.44e-20 
C6720 VCC.n2861 VSS 3.5e-20 
C6721 VCC.n2862 VSS 3e-20 
C6722 VCC.n2863 VSS 7.95e-19 
C6723 VCC.n2864 VSS 1.83e-19 
C6724 VCC.n2865 VSS 2.88e-20 
C6725 VCC.n2866 VSS 2.68e-20 
C6726 VCC.n2867 VSS 2.68e-20 
C6727 VCC.n2868 VSS 2.68e-20 
C6728 VCC.n2869 VSS 4.53e-20 
C6729 VCC.n2870 VSS 3.7e-20 
C6730 VCC.n2871 VSS 7.82e-20 
C6731 VCC.n2872 VSS 1.17e-19 
C6732 VCC.n2873 VSS 3.91e-20 
C6733 VCC.n2874 VSS 1.65e-20 
C6734 VCC.n2875 VSS 2.68e-20 
C6735 VCC.n2876 VSS 3.5e-20 
C6736 VCC.n2877 VSS 3e-20 
C6737 VCC.n2878 VSS 5.12e-19 
C6738 VCC.n2879 VSS 1.18e-19 
C6739 VCC.n2880 VSS 3.5e-20 
C6740 VCC.n2881 VSS 3.5e-20 
C6741 VCC.t293 VSS 1.55e-19 
C6742 VCC.n2882 VSS 7.57e-19 
C6743 VCC.n2883 VSS 4.73e-20 
C6744 VCC.n2884 VSS 1.54e-19 
C6745 VCC.n2885 VSS 2.88e-20 
C6746 VCC.n2886 VSS 2.88e-20 
C6747 VCC.n2887 VSS 3.5e-20 
C6748 VCC.n2888 VSS 5.76e-20 
C6749 VCC.n2889 VSS 9.88e-20 
C6750 VCC.n2890 VSS 1.3e-19 
C6751 VCC.n2891 VSS 3e-20 
C6752 VCC.t291 VSS 0.005f 
C6753 VCC.t183 VSS 0.00453f 
C6754 VCC.n2892 VSS 0.00229f 
C6755 VCC.n2893 VSS 1.91e-19 
C6756 VCC.n2894 VSS 3.5e-20 
C6757 VCC.n2895 VSS 3.14e-19 
C6758 VCC.n2896 VSS 2.47e-20 
C6759 VCC.n2897 VSS 5.76e-20 
C6760 VCC.n2898 VSS 2.47e-20 
C6761 VCC.n2899 VSS 8.23e-21 
C6762 VCC.n2900 VSS 2.88e-20 
C6763 VCC.n2901 VSS 5.76e-20 
C6764 VCC.n2902 VSS 2.47e-20 
C6765 VCC.n2903 VSS 2.88e-20 
C6766 VCC.n2904 VSS 2.47e-20 
C6767 VCC.n2905 VSS 5.15e-20 
C6768 VCC.n2906 VSS 4.73e-20 
C6769 VCC.n2907 VSS 3.7e-20 
C6770 VCC.n2908 VSS 3.5e-20 
C6771 VCC.n2909 VSS 7.41e-20 
C6772 VCC.t147 VSS 6.42e-19 
C6773 VCC.n2910 VSS 3e-20 
C6774 VCC.n2911 VSS 5.97e-20 
C6775 VCC.n2912 VSS 4.13e-19 
C6776 VCC.n2913 VSS 9.53e-20 
C6777 VCC.n2914 VSS 3.5e-20 
C6778 VCC.n2915 VSS 3.5e-20 
C6779 VCC.n2916 VSS 5.35e-20 
C6780 VCC.n2917 VSS 4.32e-20 
C6781 VCC.n2918 VSS 2.68e-20 
C6782 VCC.n2919 VSS 3.7e-20 
C6783 VCC.n2920 VSS 1.65e-20 
C6784 VCC.n2921 VSS 4.53e-20 
C6785 VCC.n2922 VSS 1.2e-19 
C6786 VCC.n2923 VSS 5.2e-19 
C6787 VCC.n2924 VSS 1.2e-19 
C6788 VCC.n2925 VSS 6.38e-20 
C6789 VCC.n2926 VSS 2.47e-20 
C6790 VCC.n2927 VSS 4.53e-20 
C6791 VCC.n2928 VSS 3.5e-20 
C6792 VCC.n2929 VSS 3.5e-20 
C6793 VCC.n2930 VSS 2.68e-20 
C6794 VCC.n2931 VSS 2.68e-20 
C6795 VCC.n2932 VSS 2.47e-20 
C6796 VCC.n2933 VSS 4.53e-20 
C6797 VCC.n2934 VSS 2.68e-20 
C6798 VCC.n2935 VSS 4.32e-20 
C6799 VCC.n2936 VSS 2.68e-20 
C6800 VCC.n2937 VSS 3.91e-20 
C6801 VCC.n2938 VSS 2.88e-20 
C6802 VCC.n2939 VSS 4.73e-20 
C6803 VCC.n2940 VSS 3.7e-20 
C6804 VCC.n2941 VSS 3.7e-20 
C6805 VCC.n2942 VSS 3.5e-20 
C6806 VCC.n2943 VSS 5.76e-20 
C6807 VCC.n2944 VSS 4.73e-20 
C6808 VCC.n2945 VSS 3.09e-20 
C6809 VCC.n2946 VSS 3.5e-20 
C6810 VCC.n2947 VSS 3.5e-20 
C6811 VCC.n2948 VSS 3.5e-20 
C6812 VCC.n2949 VSS 1.18e-19 
C6813 VCC.n2950 VSS 3e-20 
C6814 VCC.n2951 VSS 1.15e-19 
C6815 VCC.n2952 VSS 9.88e-20 
C6816 VCC.n2953 VSS 5.76e-20 
C6817 VCC.n2954 VSS 3.5e-20 
C6818 VCC.n2955 VSS 3.09e-20 
C6819 VCC.n2956 VSS 3.09e-20 
C6820 VCC.n2957 VSS 2.26e-20 
C6821 VCC.n2958 VSS 5.76e-20 
C6822 VCC.n2959 VSS 2.68e-20 
C6823 VCC.n2960 VSS 2.68e-20 
C6824 VCC.n2961 VSS 0.00185f 
C6825 VCC.n2962 VSS 2.72e-19 
C6826 VCC.n2963 VSS 2.26e-20 
C6827 VCC.n2964 VSS 1.87e-19 
C6828 VCC.n2965 VSS 3.5e-20 
C6829 VCC.n2966 VSS 2.68e-20 
C6830 VCC.n2967 VSS 5.97e-20 
C6831 VCC.n2968 VSS 4.73e-20 
C6832 VCC.n2969 VSS 4.73e-20 
C6833 VCC.n2970 VSS 5.15e-20 
C6834 VCC.n2971 VSS 7.41e-20 
C6835 VCC.n2972 VSS 3.7e-20 
C6836 VCC.n2973 VSS 2.26e-20 
C6837 VCC.n2974 VSS 6.38e-20 
C6838 VCC.n2975 VSS 4.73e-20 
C6839 VCC.n2976 VSS 3.29e-20 
C6840 VCC.n2977 VSS 3.5e-20 
C6841 VCC.n2978 VSS 3e-20 
C6842 VCC.t184 VSS 0.005f 
C6843 VCC.t127 VSS 0.00453f 
C6844 VCC.n2979 VSS 0.00228f 
C6845 VCC.n2980 VSS 1.3e-19 
C6846 VCC.t185 VSS 4.05e-19 
C6847 VCC.n2981 VSS 4.05e-19 
C6848 VCC.n2982 VSS 1.15e-19 
C6849 VCC.n2983 VSS 3.36e-19 
C6850 VCC.n2984 VSS 6.17e-21 
C6851 VCC.n2985 VSS 3.12e-19 
C6852 VCC.n2986 VSS 1.65e-20 
C6853 VCC.n2987 VSS 1.54e-19 
C6854 VCC.n2988 VSS 1.54e-19 
C6855 VCC.n2989 VSS 1.65e-20 
C6856 VCC.n2990 VSS 1.03e-20 
C6857 VCC.n2991 VSS 3.5e-20 
C6858 VCC.n2992 VSS 2.26e-20 
C6859 VCC.n2993 VSS 4.73e-20 
C6860 VCC.n2994 VSS 3.5e-20 
C6861 VCC.n2995 VSS 3e-20 
C6862 VCC.n2996 VSS 1.3e-19 
C6863 VCC.n2997 VSS 5.12e-19 
C6864 VCC.n2998 VSS 1.3e-19 
C6865 VCC.n2999 VSS 4.13e-19 
C6866 VCC.n3000 VSS 9.53e-20 
C6867 VCC.n3001 VSS 5.76e-20 
C6868 VCC.n3002 VSS 7.41e-20 
C6869 VCC.n3003 VSS 5.56e-20 
C6870 VCC.t186 VSS 1.55e-19 
C6871 VCC.n3004 VSS 3.91e-20 
C6872 VCC.n3005 VSS 3.91e-20 
C6873 VCC.n3006 VSS 1.85e-20 
C6874 VCC.n3007 VSS 7.55e-19 
C6875 VCC.n3008 VSS 4.94e-20 
C6876 VCC.n3009 VSS 5.15e-20 
C6877 VCC.n3010 VSS 7.2e-20 
C6878 VCC.n3011 VSS 1.38e-19 
C6879 VCC.n3012 VSS 1.17e-19 
C6880 VCC.n3013 VSS 4.32e-20 
C6881 VCC.n3014 VSS 2.88e-20 
C6882 VCC.n3015 VSS 2.68e-20 
C6883 VCC.n3016 VSS 3.5e-20 
C6884 VCC.n3017 VSS 3.5e-20 
C6885 VCC.n3018 VSS 2.88e-20 
C6886 VCC.n3019 VSS 2.68e-20 
C6887 VCC.n3020 VSS 2.68e-20 
C6888 VCC.n3021 VSS 2.68e-20 
C6889 VCC.n3022 VSS 4.12e-20 
C6890 VCC.n3023 VSS 4.12e-20 
C6891 VCC.n3024 VSS 3.91e-20 
C6892 VCC.n3025 VSS 4.53e-20 
C6893 VCC.n3026 VSS 4.53e-20 
C6894 VCC.n3027 VSS 1.05e-19 
C6895 VCC.n3028 VSS 1.05e-19 
C6896 VCC.n3029 VSS 4.32e-20 
C6897 VCC.n3030 VSS 3.7e-20 
C6898 VCC.n3031 VSS 2.68e-20 
C6899 VCC.n3032 VSS 2.68e-20 
C6900 VCC.n3033 VSS 6.79e-20 
C6901 VCC.n3034 VSS 9.26e-20 
C6902 VCC.n3035 VSS 1.83e-19 
C6903 VCC.n3036 VSS 7.95e-19 
C6904 VCC.n3037 VSS 5.2e-19 
C6905 VCC.n3038 VSS 1.3e-19 
C6906 VCC.n3039 VSS 3e-20 
C6907 VCC.n3040 VSS 3.5e-20 
C6908 VCC.n3041 VSS 5.97e-20 
C6909 VCC.n3042 VSS 7.41e-20 
C6910 VCC.n3043 VSS 5.15e-20 
C6911 VCC.n3044 VSS 5.15e-20 
C6912 VCC.n3045 VSS 3.09e-20 
C6913 VCC.n3046 VSS 3.09e-20 
C6914 VCC.n3047 VSS 3.7e-20 
C6915 VCC.n3048 VSS 2.68e-20 
C6916 VCC.n3049 VSS 3.91e-20 
C6917 VCC.n3050 VSS 1.17e-19 
C6918 VCC.n3051 VSS 1.38e-19 
C6919 VCC.n3052 VSS 7e-20 
C6920 VCC.n3053 VSS 4.73e-20 
C6921 VCC.n3054 VSS 3.5e-20 
C6922 VCC.n3055 VSS 3.5e-20 
C6923 VCC.n3056 VSS 3.5e-20 
C6924 VCC.n3057 VSS 4.53e-20 
C6925 VCC.n3058 VSS 1.18e-19 
C6926 VCC.n3059 VSS 5.12e-19 
C6927 VCC.n3060 VSS 1.3e-19 
C6928 VCC.n3061 VSS 1.61e-19 
C6929 VCC.n3062 VSS 9.9e-20 
C6930 VCC.n3063 VSS 0.00243f 
C6931 VCC.n3064 VSS 2.26e-20 
C6932 VCC.n3065 VSS 4.13e-19 
C6933 VCC.n3066 VSS 3.5e-20 
C6934 VCC.n3067 VSS 3.5e-20 
C6935 VCC.n3068 VSS 2.47e-20 
C6936 VCC.n3069 VSS 2.06e-20 
C6937 VCC.n3070 VSS 6.17e-20 
C6938 VCC.n3071 VSS 6.17e-20 
C6939 VCC.n3072 VSS 4.73e-20 
C6940 VCC.n3073 VSS 4.73e-20 
C6941 VCC.n3074 VSS 2.88e-20 
C6942 VCC.n3075 VSS 1.44e-20 
C6943 VCC.n3076 VSS 1.65e-20 
C6944 VCC.n3077 VSS 1.54e-19 
C6945 VCC.n3078 VSS 1.54e-19 
C6946 VCC.n3079 VSS 1.65e-20 
C6947 VCC.n3080 VSS 3.09e-20 
C6948 VCC.t148 VSS 1.55e-19 
C6949 VCC.n3081 VSS 0.00102f 
C6950 VCC.n3082 VSS 2.73e-19 
C6951 VCC.n3083 VSS 0.00136f 
C6952 VCC.n3084 VSS 2.73e-19 
C6953 VCC.n3085 VSS 0.00181f 
C6954 VCC.n3086 VSS 5.76e-20 
C6955 VCC.n3087 VSS 1.54e-19 
C6956 VCC.n3088 VSS 1.65e-20 
C6957 VCC.n3089 VSS 2.88e-20 
C6958 VCC.n3090 VSS 2.47e-20 
C6959 VCC.n3091 VSS 6.17e-20 
C6960 VCC.n3092 VSS 4.73e-20 
C6961 VCC.n3093 VSS 4.73e-20 
C6962 VCC.n3094 VSS 5.15e-20 
C6963 VCC.n3095 VSS 3.5e-20 
C6964 VCC.n3096 VSS 7.41e-20 
C6965 VCC.n3097 VSS 3.7e-20 
C6966 VCC.n3098 VSS 2.26e-20 
C6967 VCC.n3099 VSS 6.17e-20 
C6968 VCC.n3100 VSS 4.73e-20 
C6969 VCC.n3101 VSS 3.5e-20 
C6970 VCC.n3102 VSS 2.88e-20 
C6971 VCC.n3103 VSS 3.4e-19 
C6972 VCC.n3104 VSS 1.15e-19 
C6973 VCC.n3105 VSS 3.98e-19 
C6974 VCC.t292 VSS 4.05e-19 
C6975 VCC.n3106 VSS 1.22e-19 
C6976 VCC.n3107 VSS 1.3e-19 
C6977 VCC.n3108 VSS 3e-20 
C6978 VCC.n3109 VSS 3.5e-20 
C6979 VCC.n3110 VSS 3.5e-20 
C6980 VCC.n3111 VSS 4.73e-20 
C6981 VCC.n3112 VSS 2.47e-20 
C6982 VCC.n3113 VSS 1.23e-20 
C6983 VCC.n3114 VSS 1.65e-20 
C6984 VCC.n3115 VSS 2.47e-20 
C6985 VCC.n3116 VSS 5.76e-20 
C6986 VCC.n3117 VSS 1.38e-19 
C6987 VCC.n3118 VSS 7e-20 
C6988 VCC.n3119 VSS 3.7e-20 
C6989 VCC.n3120 VSS 2.47e-20 
C6990 VCC.n3121 VSS 3.7e-20 
C6991 VCC.n3122 VSS 1.85e-20 
C6992 VCC.n3123 VSS 3.09e-20 
C6993 VCC.n3124 VSS 5.35e-20 
C6994 VCC.n3125 VSS 4.73e-20 
C6995 VCC.n3126 VSS 5.35e-20 
C6996 VCC.n3127 VSS 7.41e-20 
C6997 VCC.n3128 VSS 5.76e-20 
C6998 VCC.n3129 VSS 9.53e-20 
C6999 VCC.n3130 VSS 4.13e-19 
C7000 VCC.n3131 VSS 1.3e-19 
C7001 VCC.n3132 VSS 5.2e-19 
C7002 VCC.n3133 VSS 1.2e-19 
C7003 VCC.n3134 VSS 4.73e-20 
C7004 VCC.n3135 VSS 2.68e-20 
C7005 VCC.n3136 VSS 3.5e-20 
C7006 VCC.n3137 VSS 3.5e-20 
C7007 VCC.n3138 VSS 2.68e-20 
C7008 VCC.n3139 VSS 2.68e-20 
C7009 VCC.n3140 VSS 4.32e-20 
C7010 VCC.n3141 VSS 4.32e-20 
C7011 VCC.n3142 VSS 4.32e-20 
C7012 VCC.n3143 VSS 2.88e-20 
C7013 VCC.n3144 VSS 3.5e-20 
C7014 VCC.n3145 VSS 2.68e-20 
C7015 VCC.n3146 VSS 7.82e-20 
C7016 VCC.n3147 VSS 4.73e-20 
C7017 VCC.n3148 VSS 4.73e-20 
C7018 VCC.n3149 VSS 1.05e-19 
C7019 VCC.n3150 VSS 1.05e-19 
C7020 VCC.n3151 VSS 4.53e-20 
C7021 VCC.n3152 VSS 2.68e-20 
C7022 VCC.n3153 VSS 2.68e-20 
C7023 VCC.n3154 VSS 6.59e-20 
C7024 VCC.n3155 VSS 9.26e-20 
C7025 VCC.n3156 VSS 6.59e-20 
C7026 VCC.n3157 VSS 2.47e-20 
C7027 VCC.n3158 VSS 2.47e-20 
C7028 VCC.n3159 VSS 2.88e-20 
C7029 VCC.n3160 VSS 3.5e-20 
C7030 VCC.n3161 VSS 3.5e-20 
C7031 VCC.n3162 VSS 4.53e-20 
C7032 VCC.n3163 VSS 1.2e-19 
C7033 VCC.n3164 VSS 5.2e-19 
C7034 VCC.n3165 VSS 1.3e-19 
C7035 VCC.n3166 VSS 4.13e-19 
C7036 VCC.n3167 VSS 9.53e-20 
C7037 VCC.n3168 VSS 5.97e-20 
C7038 VCC.n3169 VSS 7.41e-20 
C7039 VCC.n3170 VSS 5.35e-20 
C7040 VCC.n3171 VSS 5.15e-20 
C7041 VCC.n3172 VSS 3.09e-20 
C7042 VCC.n3173 VSS 3.09e-20 
C7043 VCC.n3174 VSS 3.91e-20 
C7044 VCC.n3175 VSS 2.47e-20 
C7045 VCC.n3176 VSS 3.7e-20 
C7046 VCC.n3177 VSS 1.17e-19 
C7047 VCC.n3178 VSS 1.38e-19 
C7048 VCC.n3179 VSS 7.2e-20 
C7049 VCC.n3180 VSS 4.73e-20 
C7050 VCC.n3181 VSS 3.5e-20 
C7051 VCC.n3182 VSS 3.5e-20 
C7052 VCC.n3183 VSS 4.53e-20 
C7053 VCC.n3184 VSS 5.97e-20 
C7054 VCC.n3185 VSS 3.5e-20 
C7055 VCC.n3186 VSS 3e-20 
C7056 VCC.n3187 VSS 1.3e-19 
C7057 VCC.n3188 VSS 1.53e-19 
C7058 VCC.t230 VSS 4.05e-19 
C7059 VCC.n3189 VSS 2.06e-19 
C7060 VCC.n3190 VSS 1.35e-19 
C7061 VCC.n3191 VSS 9.67e-20 
C7062 VCC.n3192 VSS 3.35e-20 
C7063 VCC.n3193 VSS 3.5e-20 
C7064 VCC.n3194 VSS 2.36e-19 
C7065 VCC.n3195 VSS 0.0023f 
C7066 VCC.t94 VSS 0.0031f 
C7067 VCC.t272 VSS 0.00366f 
C7068 VCC.t97 VSS 0.00365f 
C7069 VCC.t273 VSS 0.00386f 
C7070 VCC.n3196 VSS 0.00569f 
C7071 VCC.n3197 VSS 1.3e-19 
C7072 VCC.n3198 VSS 3.67e-19 
C7073 VCC.n3199 VSS 1.15e-19 
C7074 VCC.n3200 VSS 3.38e-19 
C7075 VCC.n3201 VSS 3.5e-20 
C7076 VCC.n3202 VSS 3.5e-20 
C7077 VCC.n3203 VSS 2.68e-20 
C7078 VCC.n3204 VSS 2.06e-20 
C7079 VCC.n3205 VSS 6.38e-20 
C7080 VCC.n3206 VSS 5.97e-20 
C7081 VCC.n3207 VSS 4.73e-20 
C7082 VCC.n3208 VSS 4.73e-20 
C7083 VCC.n3209 VSS 3.09e-20 
C7084 VCC.n3210 VSS 1.23e-20 
C7085 VCC.n3211 VSS 1.65e-20 
C7086 VCC.n3212 VSS 1.54e-19 
C7087 VCC.n3213 VSS 1.54e-19 
C7088 VCC.n3214 VSS 1.65e-20 
C7089 VCC.n3215 VSS 3.29e-20 
C7090 VCC.t231 VSS 1.67e-19 
C7091 VCC.n3216 VSS 0.00101f 
C7092 VCC.n3217 VSS 2.71e-19 
C7093 VCC.n3218 VSS 7.46e-19 
C7094 VCC.n3219 VSS 0.00333f 
C7095 VCC.n3220 VSS 2.46e-19 
C7096 VCC.n3221 VSS 3.02e-19 
C7097 VCC.n3222 VSS 3.7e-20 
C7098 VCC.n3223 VSS 5.15e-20 
C7099 VCC.n3224 VSS 6.38e-20 
C7100 VCC.n3225 VSS 4.73e-20 
C7101 VCC.n3226 VSS 4.73e-20 
C7102 VCC.n3227 VSS 2.68e-20 
C7103 VCC.n3228 VSS 3.29e-20 
C7104 VCC.n3229 VSS 1.65e-20 
C7105 VCC.n3230 VSS 1.54e-19 
C7106 VCC.n3231 VSS 1.54e-19 
C7107 VCC.n3232 VSS 5.56e-20 
C7108 VCC.n3233 VSS 2.88e-20 
C7109 VCC.n3234 VSS 1.65e-20 
C7110 VCC.n3235 VSS 3.09e-20 
C7111 VCC.n3236 VSS 4.73e-20 
C7112 VCC.n3237 VSS 4.73e-20 
C7113 VCC.n3238 VSS 4.32e-20 
C7114 VCC.n3239 VSS 1.17e-19 
C7115 VCC.n3240 VSS 3.33e-19 
C7116 VCC.n3241 VSS 1.35e-19 
C7117 VCC.n3242 VSS 4.37e-19 
C7118 VCC.n3243 VSS 5.24e-19 
C7119 VCC.n3244 VSS 1.36e-19 
C7120 VCC.n3245 VSS 1.01e-19 
C7121 VCC.n3246 VSS 1.05e-19 
C7122 VCC.n3247 VSS 2.06e-20 
C7123 VCC.n3248 VSS 2.26e-20 
C7124 VCC.n3249 VSS 3.7e-20 
C7125 VCC.n3250 VSS 5.15e-20 
C7126 VCC.n3251 VSS 1.38e-19 
C7127 VCC.n3252 VSS 3.91e-20 
C7128 VCC.n3253 VSS 2.88e-20 
C7129 VCC.n3254 VSS 4.32e-20 
C7130 VCC.n3255 VSS 1.17e-19 
C7131 VCC.n3256 VSS 3.7e-20 
C7132 VCC.n3257 VSS 3.91e-20 
C7133 VCC.n3258 VSS 3.5e-20 
C7134 VCC.n3259 VSS 1.65e-20 
C7135 VCC.n3260 VSS 8.23e-21 
C7136 VCC.n3261 VSS 3.5e-20 
C7137 VCC.n3262 VSS 3.5e-20 
C7138 VCC.n3263 VSS 1.4e-19 
C7139 VCC.n3264 VSS 5.4e-19 
C7140 VCC.n3265 VSS 8.42e-19 
C7141 VCC.n3266 VSS 5.4e-19 
C7142 VCC.n3267 VSS 1.4e-19 
C7143 VCC.n3268 VSS 1.4e-19 
C7144 VCC.n3269 VSS 2.18e-19 
C7145 VCC.n3270 VSS 7.82e-20 
C7146 VCC.n3271 VSS 4.32e-20 
C7147 VCC.n3272 VSS 4.32e-20 
C7148 VCC.n3273 VSS 1.05e-19 
C7149 VCC.n3274 VSS 1.05e-19 
C7150 VCC.n3275 VSS 4.32e-20 
C7151 VCC.n3276 VSS 3.7e-20 
C7152 VCC.n3277 VSS 2.68e-20 
C7153 VCC.n3278 VSS 5.76e-20 
C7154 VCC.n3279 VSS 6.38e-20 
C7155 VCC.n3280 VSS 3.5e-20 
C7156 VCC.n3281 VSS 3.5e-20 
C7157 VCC.n3282 VSS 1.17e-19 
C7158 VCC.n3283 VSS 1.38e-19 
C7159 VCC.n3284 VSS 5.15e-20 
C7160 VCC.n3285 VSS 1.05e-19 
C7161 VCC.n3286 VSS 2.26e-20 
C7162 VCC.n3287 VSS 5.76e-20 
C7163 VCC.n3288 VSS 3.7e-20 
C7164 VCC.n3289 VSS 3.7e-20 
C7165 VCC.n3290 VSS 3.09e-20 
C7166 VCC.n3291 VSS 1.85e-20 
C7167 VCC.n3292 VSS 1.65e-20 
C7168 VCC.n3293 VSS 8.23e-21 
C7169 VCC.n3294 VSS 1.13e-19 
C7170 VCC.n3295 VSS 3.33e-19 
C7171 VCC.t198 VSS 4.21e-19 
C7172 VCC.n3296 VSS 2.06e-19 
C7173 VCC.n3297 VSS 1.35e-19 
C7174 VCC.n3298 VSS 3.5e-20 
C7175 VCC.n3299 VSS 3.5e-20 
C7176 VCC.n3300 VSS 3.5e-20 
C7177 VCC.n3301 VSS 1.03e-20 
C7178 VCC.n3302 VSS 2.68e-20 
C7179 VCC.n3303 VSS 3.09e-20 
C7180 VCC.n3304 VSS 2.68e-20 
C7181 VCC.n3305 VSS 1.65e-20 
C7182 VCC.n3306 VSS 1.54e-19 
C7183 VCC.n3307 VSS 1.54e-19 
C7184 VCC.n3308 VSS 1.65e-20 
C7185 VCC.t199 VSS 1.56e-19 
C7186 VCC.n3309 VSS 7.62e-19 
C7187 VCC.n3310 VSS 1.23e-20 
C7188 VCC.n3311 VSS 2.47e-20 
C7189 VCC.n3312 VSS 4.73e-20 
C7190 VCC.n3313 VSS 6.59e-20 
C7191 VCC.n3314 VSS 5.15e-20 
C7192 VCC.n3315 VSS 2.47e-20 
C7193 VCC.n3316 VSS 7.41e-20 
C7194 VCC.n3317 VSS 9.47e-20 
C7195 VCC.n3318 VSS 1.32e-19 
C7196 VCC.n3319 VSS 7.71e-19 
C7197 VCC.n3320 VSS 9.83e-19 
C7198 VCC.n3321 VSS 2.36e-19 
C7199 VCC.n3322 VSS 3.21e-19 
C7200 VCC.n3323 VSS 2.61e-19 
C7201 VCC.n3324 VSS 0.00189f 
C7202 VCC.n3325 VSS 0.00274f 
C7203 VCC.n3326 VSS 5.76e-20 
C7204 VCC.n3327 VSS 2.88e-20 
C7205 VCC.n3328 VSS 3.5e-20 
C7206 VCC.n3329 VSS 9.83e-19 
C7207 VCC.n3330 VSS 9.47e-20 
C7208 VCC.n3331 VSS 1.17e-19 
C7209 VCC.n3332 VSS 2.06e-19 
C7210 VCC.n3333 VSS 1.36e-19 
C7211 VCC.n3334 VSS 1.01e-19 
C7212 VCC.n3335 VSS 3.5e-20 
C7213 VCC.n3336 VSS 3.09e-20 
C7214 VCC.n3337 VSS 3.29e-20 
C7215 VCC.n3338 VSS 3.29e-20 
C7216 VCC.n3339 VSS 4.73e-20 
C7217 VCC.n3340 VSS 1.44e-20 
C7218 VCC.n3341 VSS 3.5e-20 
C7219 VCC.n3342 VSS 7.41e-20 
C7220 VCC.n3343 VSS 2.47e-20 
C7221 VCC.t275 VSS 1.56e-19 
C7222 VCC.n3344 VSS 5.76e-20 
C7223 VCC.n3345 VSS 2.06e-20 
C7224 VCC.n3346 VSS 5.76e-20 
C7225 VCC.n3347 VSS 3.7e-20 
C7226 VCC.n3348 VSS 4.32e-20 
C7227 VCC.n3349 VSS 2.68e-20 
C7228 VCC.n3350 VSS 3.91e-20 
C7229 VCC.n3351 VSS 6.38e-20 
C7230 VCC.n3352 VSS 1.85e-20 
C7231 VCC.n3353 VSS 3.5e-20 
C7232 VCC.n3354 VSS 3.09e-20 
C7233 VCC.n3355 VSS 3.7e-20 
C7234 VCC.n3356 VSS 3.09e-20 
C7235 VCC.n3357 VSS 2.26e-20 
C7236 VCC.n3358 VSS 1.05e-19 
C7237 VCC.n3359 VSS 3.5e-20 
C7238 VCC.n3360 VSS 3.5e-20 
C7239 VCC.n3361 VSS 8.42e-19 
C7240 VCC.n3362 VSS 2.18e-19 
C7241 VCC.n3363 VSS 1.4e-19 
C7242 VCC.n3364 VSS 4.32e-20 
C7243 VCC.n3365 VSS 7.82e-20 
C7244 VCC.n3366 VSS 5.76e-20 
C7245 VCC.n3367 VSS 2.68e-20 
C7246 VCC.n3368 VSS 4.32e-20 
C7247 VCC.n3369 VSS 3.91e-20 
C7248 VCC.n3370 VSS 3.7e-20 
C7249 VCC.n3371 VSS 3.7e-20 
C7250 VCC.n3372 VSS 5.76e-20 
C7251 VCC.n3373 VSS 4.73e-20 
C7252 VCC.n3374 VSS 3.5e-20 
C7253 VCC.t270 VSS 1.56e-19 
C7254 VCC.n3375 VSS 7.97e-19 
C7255 VCC.n3376 VSS 3.09e-20 
C7256 VCC.n3377 VSS 1.01e-19 
C7257 VCC.n3378 VSS 3.5e-20 
C7258 VCC.n3379 VSS 1.36e-19 
C7259 VCC.n3380 VSS 3.5e-20 
C7260 VCC.n3381 VSS 3.33e-19 
C7261 VCC.n3382 VSS 1.17e-19 
C7262 VCC.n3383 VSS 1.09e-19 
C7263 VCC.n3384 VSS 3.5e-20 
C7264 VCC.n3385 VSS 4.73e-20 
C7265 VCC.n3386 VSS 5.56e-20 
C7266 VCC.n3387 VSS 2.88e-20 
C7267 VCC.n3388 VSS 2.26e-20 
C7268 VCC.n3389 VSS 5.76e-20 
C7269 VCC.n3390 VSS 2.68e-20 
C7270 VCC.n3391 VSS 2.68e-20 
C7271 VCC.n3392 VSS 1.9e-19 
C7272 VCC.n3393 VSS 5.76e-20 
C7273 VCC.n3394 VSS 2.68e-20 
C7274 VCC.n3395 VSS 2.68e-20 
C7275 VCC.n3396 VSS 2.68e-20 
C7276 VCC.n3397 VSS 5.76e-20 
C7277 VCC.n3398 VSS 2.26e-20 
C7278 VCC.n3399 VSS 3.09e-20 
C7279 VCC.n3400 VSS 2.26e-20 
C7280 VCC.n3401 VSS 5.15e-20 
C7281 VCC.n3402 VSS 4.73e-20 
C7282 VCC.n3403 VSS 3.7e-20 
C7283 VCC.n3404 VSS 3.5e-20 
C7284 VCC.n3405 VSS 7.41e-20 
C7285 VCC.n3406 VSS 1.91e-19 
C7286 VCC.n3407 VSS 9.88e-20 
C7287 VCC.n3408 VSS 3e-20 
C7288 VCC.n3409 VSS 5.12e-19 
C7289 VCC.n3410 VSS 1.18e-19 
C7290 VCC.n3411 VSS 3.5e-20 
C7291 VCC.n3412 VSS 3.5e-20 
C7292 VCC.n3413 VSS 5.15e-20 
C7293 VCC.n3414 VSS 4.32e-20 
C7294 VCC.n3415 VSS 2.68e-20 
C7295 VCC.n3416 VSS 3.91e-20 
C7296 VCC.n3417 VSS 1.44e-20 
C7297 VCC.n3418 VSS 3.5e-20 
C7298 VCC.n3419 VSS 3e-20 
C7299 VCC.n3420 VSS 7.95e-19 
C7300 VCC.n3421 VSS 1.83e-19 
C7301 VCC.n3422 VSS 2.88e-20 
C7302 VCC.n3423 VSS 2.68e-20 
C7303 VCC.n3424 VSS 2.68e-20 
C7304 VCC.n3425 VSS 2.68e-20 
C7305 VCC.n3426 VSS 4.53e-20 
C7306 VCC.n3427 VSS 3.7e-20 
C7307 VCC.n3428 VSS 7.82e-20 
C7308 VCC.n3429 VSS 1.17e-19 
C7309 VCC.n3430 VSS 3.91e-20 
C7310 VCC.n3431 VSS 1.65e-20 
C7311 VCC.n3432 VSS 2.68e-20 
C7312 VCC.n3433 VSS 3.5e-20 
C7313 VCC.n3434 VSS 3e-20 
C7314 VCC.n3435 VSS 5.12e-19 
C7315 VCC.n3436 VSS 1.18e-19 
C7316 VCC.n3437 VSS 3.5e-20 
C7317 VCC.n3438 VSS 3.5e-20 
C7318 VCC.t179 VSS 1.55e-19 
C7319 VCC.n3439 VSS 7.57e-19 
C7320 VCC.n3440 VSS 4.73e-20 
C7321 VCC.n3441 VSS 1.54e-19 
C7322 VCC.n3442 VSS 2.88e-20 
C7323 VCC.n3443 VSS 2.88e-20 
C7324 VCC.n3444 VSS 3.5e-20 
C7325 VCC.n3445 VSS 5.76e-20 
C7326 VCC.n3446 VSS 9.88e-20 
C7327 VCC.n3447 VSS 1.3e-19 
C7328 VCC.n3448 VSS 3e-20 
C7329 VCC.t180 VSS 0.005f 
C7330 VCC.t93 VSS 0.00453f 
C7331 VCC.n3449 VSS 0.00229f 
C7332 VCC.n3450 VSS 1.91e-19 
C7333 VCC.n3451 VSS 3.5e-20 
C7334 VCC.n3452 VSS 3.14e-19 
C7335 VCC.n3453 VSS 3.5e-20 
C7336 VCC.n3454 VSS 2.47e-20 
C7337 VCC.n3455 VSS 5.76e-20 
C7338 VCC.n3456 VSS 2.47e-20 
C7339 VCC.n3457 VSS 8.23e-21 
C7340 VCC.n3458 VSS 2.88e-20 
C7341 VCC.n3459 VSS 5.76e-20 
C7342 VCC.n3460 VSS 2.47e-20 
C7343 VCC.n3461 VSS 2.88e-20 
C7344 VCC.n3462 VSS 2.47e-20 
C7345 VCC.n3463 VSS 5.15e-20 
C7346 VCC.n3464 VSS 4.73e-20 
C7347 VCC.n3465 VSS 3.7e-20 
C7348 VCC.n3466 VSS 3.5e-20 
C7349 VCC.n3467 VSS 7.41e-20 
C7350 VCC.t311 VSS 6.42e-19 
C7351 VCC.n3468 VSS 3e-20 
C7352 VCC.n3469 VSS 5.97e-20 
C7353 VCC.n3470 VSS 4.13e-19 
C7354 VCC.n3471 VSS 9.53e-20 
C7355 VCC.n3472 VSS 3.5e-20 
C7356 VCC.n3473 VSS 3.5e-20 
C7357 VCC.n3474 VSS 5.35e-20 
C7358 VCC.n3475 VSS 4.32e-20 
C7359 VCC.n3476 VSS 2.68e-20 
C7360 VCC.n3477 VSS 3.7e-20 
C7361 VCC.n3478 VSS 1.65e-20 
C7362 VCC.n3479 VSS 4.53e-20 
C7363 VCC.n3480 VSS 1.2e-19 
C7364 VCC.n3481 VSS 5.2e-19 
C7365 VCC.n3482 VSS 1.2e-19 
C7366 VCC.n3483 VSS 6.38e-20 
C7367 VCC.n3484 VSS 2.47e-20 
C7368 VCC.n3485 VSS 4.53e-20 
C7369 VCC.n3486 VSS 3.5e-20 
C7370 VCC.n3487 VSS 3.5e-20 
C7371 VCC.n3488 VSS 2.68e-20 
C7372 VCC.n3489 VSS 2.68e-20 
C7373 VCC.n3490 VSS 2.47e-20 
C7374 VCC.n3491 VSS 4.53e-20 
C7375 VCC.n3492 VSS 2.68e-20 
C7376 VCC.n3493 VSS 4.32e-20 
C7377 VCC.n3494 VSS 2.68e-20 
C7378 VCC.n3495 VSS 3.91e-20 
C7379 VCC.n3496 VSS 2.88e-20 
C7380 VCC.n3497 VSS 4.73e-20 
C7381 VCC.n3498 VSS 3.7e-20 
C7382 VCC.n3499 VSS 3.7e-20 
C7383 VCC.n3500 VSS 3.5e-20 
C7384 VCC.n3501 VSS 5.76e-20 
C7385 VCC.n3502 VSS 4.73e-20 
C7386 VCC.n3503 VSS 3.09e-20 
C7387 VCC.n3504 VSS 3.5e-20 
C7388 VCC.n3505 VSS 3.5e-20 
C7389 VCC.n3506 VSS 3.5e-20 
C7390 VCC.n3507 VSS 1.18e-19 
C7391 VCC.n3508 VSS 3e-20 
C7392 VCC.n3509 VSS 1.15e-19 
C7393 VCC.n3510 VSS 9.88e-20 
C7394 VCC.n3511 VSS 5.76e-20 
C7395 VCC.n3512 VSS 3.5e-20 
C7396 VCC.n3513 VSS 3.09e-20 
C7397 VCC.n3514 VSS 3.09e-20 
C7398 VCC.n3515 VSS 2.26e-20 
C7399 VCC.n3516 VSS 5.76e-20 
C7400 VCC.n3517 VSS 2.68e-20 
C7401 VCC.n3518 VSS 2.68e-20 
C7402 VCC.n3519 VSS 0.00185f 
C7403 VCC.n3520 VSS 2.72e-19 
C7404 VCC.n3521 VSS 2.26e-20 
C7405 VCC.n3522 VSS 1.87e-19 
C7406 VCC.n3523 VSS 3.5e-20 
C7407 VCC.n3524 VSS 2.68e-20 
C7408 VCC.n3525 VSS 5.97e-20 
C7409 VCC.n3526 VSS 4.73e-20 
C7410 VCC.n3527 VSS 4.73e-20 
C7411 VCC.n3528 VSS 5.15e-20 
C7412 VCC.n3529 VSS 7.41e-20 
C7413 VCC.n3530 VSS 3.7e-20 
C7414 VCC.n3531 VSS 2.26e-20 
C7415 VCC.n3532 VSS 6.38e-20 
C7416 VCC.n3533 VSS 4.73e-20 
C7417 VCC.n3534 VSS 3.29e-20 
C7418 VCC.n3535 VSS 3.5e-20 
C7419 VCC.n3536 VSS 3e-20 
C7420 VCC.t286 VSS 0.005f 
C7421 VCC.t177 VSS 0.00453f 
C7422 VCC.n3537 VSS 0.00228f 
C7423 VCC.n3538 VSS 1.3e-19 
C7424 VCC.t287 VSS 4.05e-19 
C7425 VCC.n3539 VSS 4.05e-19 
C7426 VCC.n3540 VSS 1.15e-19 
C7427 VCC.n3541 VSS 3.36e-19 
C7428 VCC.n3542 VSS 6.17e-21 
C7429 VCC.n3543 VSS 3.12e-19 
C7430 VCC.n3544 VSS 1.65e-20 
C7431 VCC.n3545 VSS 1.54e-19 
C7432 VCC.n3546 VSS 1.54e-19 
C7433 VCC.n3547 VSS 1.65e-20 
C7434 VCC.n3548 VSS 1.03e-20 
C7435 VCC.n3549 VSS 3.5e-20 
C7436 VCC.n3550 VSS 2.26e-20 
C7437 VCC.n3551 VSS 4.73e-20 
C7438 VCC.n3552 VSS 3.5e-20 
C7439 VCC.n3553 VSS 3e-20 
C7440 VCC.n3554 VSS 1.3e-19 
C7441 VCC.n3555 VSS 5.12e-19 
C7442 VCC.n3556 VSS 1.3e-19 
C7443 VCC.n3557 VSS 4.13e-19 
C7444 VCC.n3558 VSS 9.53e-20 
C7445 VCC.n3559 VSS 5.76e-20 
C7446 VCC.n3560 VSS 7.41e-20 
C7447 VCC.n3561 VSS 5.56e-20 
C7448 VCC.t288 VSS 1.55e-19 
C7449 VCC.n3562 VSS 3.91e-20 
C7450 VCC.n3563 VSS 3.91e-20 
C7451 VCC.n3564 VSS 1.85e-20 
C7452 VCC.n3565 VSS 7.55e-19 
C7453 VCC.n3566 VSS 4.94e-20 
C7454 VCC.n3567 VSS 5.15e-20 
C7455 VCC.n3568 VSS 7.2e-20 
C7456 VCC.n3569 VSS 1.38e-19 
C7457 VCC.n3570 VSS 1.17e-19 
C7458 VCC.n3571 VSS 4.32e-20 
C7459 VCC.n3572 VSS 2.88e-20 
C7460 VCC.n3573 VSS 2.68e-20 
C7461 VCC.n3574 VSS 3.5e-20 
C7462 VCC.n3575 VSS 3.5e-20 
C7463 VCC.n3576 VSS 2.88e-20 
C7464 VCC.n3577 VSS 2.68e-20 
C7465 VCC.n3578 VSS 2.68e-20 
C7466 VCC.n3579 VSS 2.68e-20 
C7467 VCC.n3580 VSS 4.12e-20 
C7468 VCC.n3581 VSS 4.12e-20 
C7469 VCC.n3582 VSS 3.91e-20 
C7470 VCC.n3583 VSS 4.53e-20 
C7471 VCC.n3584 VSS 4.53e-20 
C7472 VCC.n3585 VSS 1.05e-19 
C7473 VCC.n3586 VSS 1.05e-19 
C7474 VCC.n3587 VSS 4.32e-20 
C7475 VCC.n3588 VSS 3.7e-20 
C7476 VCC.n3589 VSS 2.68e-20 
C7477 VCC.n3590 VSS 2.68e-20 
C7478 VCC.n3591 VSS 6.79e-20 
C7479 VCC.n3592 VSS 9.26e-20 
C7480 VCC.n3593 VSS 1.83e-19 
C7481 VCC.n3594 VSS 7.95e-19 
C7482 VCC.n3595 VSS 5.2e-19 
C7483 VCC.n3596 VSS 1.3e-19 
C7484 VCC.n3597 VSS 3e-20 
C7485 VCC.n3598 VSS 3.5e-20 
C7486 VCC.n3599 VSS 5.97e-20 
C7487 VCC.n3600 VSS 7.41e-20 
C7488 VCC.n3601 VSS 5.15e-20 
C7489 VCC.n3602 VSS 5.15e-20 
C7490 VCC.n3603 VSS 3.09e-20 
C7491 VCC.n3604 VSS 3.09e-20 
C7492 VCC.n3605 VSS 3.7e-20 
C7493 VCC.n3606 VSS 2.68e-20 
C7494 VCC.n3607 VSS 3.91e-20 
C7495 VCC.n3608 VSS 1.17e-19 
C7496 VCC.n3609 VSS 1.38e-19 
C7497 VCC.n3610 VSS 7e-20 
C7498 VCC.n3611 VSS 4.73e-20 
C7499 VCC.n3612 VSS 3.5e-20 
C7500 VCC.n3613 VSS 3.5e-20 
C7501 VCC.n3614 VSS 3.5e-20 
C7502 VCC.n3615 VSS 4.53e-20 
C7503 VCC.n3616 VSS 1.18e-19 
C7504 VCC.n3617 VSS 5.12e-19 
C7505 VCC.n3618 VSS 1.3e-19 
C7506 VCC.n3619 VSS 1.61e-19 
C7507 VCC.n3620 VSS 9.9e-20 
C7508 VCC.n3621 VSS 0.00243f 
C7509 VCC.n3622 VSS 2.26e-20 
C7510 VCC.n3623 VSS 4.13e-19 
C7511 VCC.n3624 VSS 3.5e-20 
C7512 VCC.n3625 VSS 3.5e-20 
C7513 VCC.n3626 VSS 2.47e-20 
C7514 VCC.n3627 VSS 2.06e-20 
C7515 VCC.n3628 VSS 6.17e-20 
C7516 VCC.n3629 VSS 6.17e-20 
C7517 VCC.n3630 VSS 4.73e-20 
C7518 VCC.n3631 VSS 4.73e-20 
C7519 VCC.n3632 VSS 2.88e-20 
C7520 VCC.n3633 VSS 1.44e-20 
C7521 VCC.n3634 VSS 1.65e-20 
C7522 VCC.n3635 VSS 1.54e-19 
C7523 VCC.n3636 VSS 1.54e-19 
C7524 VCC.n3637 VSS 1.65e-20 
C7525 VCC.n3638 VSS 3.09e-20 
C7526 VCC.t312 VSS 1.55e-19 
C7527 VCC.n3639 VSS 0.00102f 
C7528 VCC.n3640 VSS 2.73e-19 
C7529 VCC.n3641 VSS 0.00136f 
C7530 VCC.n3642 VSS 2.73e-19 
C7531 VCC.n3643 VSS 0.00181f 
C7532 VCC.n3644 VSS 5.76e-20 
C7533 VCC.n3645 VSS 1.54e-19 
C7534 VCC.n3646 VSS 1.65e-20 
C7535 VCC.n3647 VSS 6.17e-20 
C7536 VCC.n3648 VSS 2.47e-20 
C7537 VCC.n3649 VSS 4.73e-20 
C7538 VCC.n3650 VSS 4.73e-20 
C7539 VCC.n3651 VSS 5.15e-20 
C7540 VCC.n3652 VSS 3.5e-20 
C7541 VCC.n3653 VSS 7.41e-20 
C7542 VCC.n3654 VSS 3.7e-20 
C7543 VCC.n3655 VSS 2.26e-20 
C7544 VCC.n3656 VSS 6.17e-20 
C7545 VCC.n3657 VSS 4.73e-20 
C7546 VCC.n3658 VSS 2.88e-20 
C7547 VCC.n3659 VSS 2.88e-20 
C7548 VCC.n3660 VSS 3.4e-19 
C7549 VCC.n3661 VSS 1.15e-19 
C7550 VCC.n3662 VSS 3.98e-19 
C7551 VCC.t178 VSS 4.05e-19 
C7552 VCC.n3663 VSS 1.22e-19 
C7553 VCC.n3664 VSS 1.3e-19 
C7554 VCC.n3665 VSS 3e-20 
C7555 VCC.n3666 VSS 3.5e-20 
C7556 VCC.n3667 VSS 3.5e-20 
C7557 VCC.n3668 VSS 4.73e-20 
C7558 VCC.n3669 VSS 2.47e-20 
C7559 VCC.n3670 VSS 1.23e-20 
C7560 VCC.n3671 VSS 1.65e-20 
C7561 VCC.n3672 VSS 2.47e-20 
C7562 VCC.n3673 VSS 5.76e-20 
C7563 VCC.n3674 VSS 1.38e-19 
C7564 VCC.n3675 VSS 7e-20 
C7565 VCC.n3676 VSS 3.7e-20 
C7566 VCC.n3677 VSS 2.47e-20 
C7567 VCC.n3678 VSS 3.7e-20 
C7568 VCC.n3679 VSS 1.85e-20 
C7569 VCC.n3680 VSS 3.09e-20 
C7570 VCC.n3681 VSS 5.35e-20 
C7571 VCC.n3682 VSS 4.73e-20 
C7572 VCC.n3683 VSS 5.35e-20 
C7573 VCC.n3684 VSS 7.41e-20 
C7574 VCC.n3685 VSS 5.76e-20 
C7575 VCC.n3686 VSS 9.53e-20 
C7576 VCC.n3687 VSS 4.13e-19 
C7577 VCC.n3688 VSS 1.3e-19 
C7578 VCC.n3689 VSS 5.2e-19 
C7579 VCC.n3690 VSS 1.2e-19 
C7580 VCC.n3691 VSS 4.73e-20 
C7581 VCC.n3692 VSS 2.68e-20 
C7582 VCC.n3693 VSS 3.5e-20 
C7583 VCC.n3694 VSS 3.5e-20 
C7584 VCC.n3695 VSS 2.68e-20 
C7585 VCC.n3696 VSS 2.68e-20 
C7586 VCC.n3697 VSS 4.32e-20 
C7587 VCC.n3698 VSS 4.32e-20 
C7588 VCC.n3699 VSS 4.32e-20 
C7589 VCC.n3700 VSS 2.88e-20 
C7590 VCC.n3701 VSS 3.5e-20 
C7591 VCC.n3702 VSS 2.68e-20 
C7592 VCC.n3703 VSS 7.82e-20 
C7593 VCC.n3704 VSS 4.73e-20 
C7594 VCC.n3705 VSS 4.73e-20 
C7595 VCC.n3706 VSS 1.05e-19 
C7596 VCC.n3707 VSS 1.05e-19 
C7597 VCC.n3708 VSS 4.53e-20 
C7598 VCC.n3709 VSS 2.68e-20 
C7599 VCC.n3710 VSS 2.68e-20 
C7600 VCC.n3711 VSS 6.59e-20 
C7601 VCC.n3712 VSS 9.26e-20 
C7602 VCC.n3713 VSS 6.59e-20 
C7603 VCC.n3714 VSS 2.47e-20 
C7604 VCC.n3715 VSS 2.47e-20 
C7605 VCC.n3716 VSS 2.88e-20 
C7606 VCC.n3717 VSS 3.5e-20 
C7607 VCC.n3718 VSS 3.5e-20 
C7608 VCC.n3719 VSS 4.53e-20 
C7609 VCC.n3720 VSS 1.2e-19 
C7610 VCC.n3721 VSS 5.2e-19 
C7611 VCC.n3722 VSS 1.3e-19 
C7612 VCC.n3723 VSS 4.13e-19 
C7613 VCC.n3724 VSS 9.53e-20 
C7614 VCC.n3725 VSS 5.97e-20 
C7615 VCC.n3726 VSS 7.41e-20 
C7616 VCC.n3727 VSS 5.35e-20 
C7617 VCC.n3728 VSS 5.15e-20 
C7618 VCC.n3729 VSS 3.09e-20 
C7619 VCC.n3730 VSS 3.09e-20 
C7620 VCC.n3731 VSS 3.91e-20 
C7621 VCC.n3732 VSS 2.47e-20 
C7622 VCC.n3733 VSS 3.7e-20 
C7623 VCC.n3734 VSS 1.17e-19 
C7624 VCC.n3735 VSS 1.38e-19 
C7625 VCC.n3736 VSS 7.2e-20 
C7626 VCC.n3737 VSS 4.73e-20 
C7627 VCC.n3738 VSS 3.5e-20 
C7628 VCC.n3739 VSS 3.5e-20 
C7629 VCC.n3740 VSS 4.53e-20 
C7630 VCC.n3741 VSS 5.97e-20 
C7631 VCC.n3742 VSS 3.5e-20 
C7632 VCC.n3743 VSS 3e-20 
C7633 VCC.n3744 VSS 1.3e-19 
C7634 VCC.n3745 VSS 1.53e-19 
C7635 VCC.t181 VSS 4.05e-19 
C7636 VCC.n3746 VSS 1.35e-19 
C7637 VCC.t269 VSS 4.21e-19 
C7638 VCC.n3747 VSS 2.06e-19 
C7639 VCC.n3748 VSS 1.32e-19 
C7640 VCC.n3749 VSS 9.67e-20 
C7641 VCC.n3750 VSS 3.35e-20 
C7642 VCC.n3751 VSS 3.5e-20 
C7643 VCC.n3752 VSS 2.36e-19 
C7644 VCC.n3753 VSS 0.0023f 
C7645 VCC.t268 VSS 0.0031f 
C7646 VCC.t98 VSS 0.00366f 
C7647 VCC.t271 VSS 0.00365f 
C7648 VCC.t101 VSS 0.00386f 
C7649 VCC.n3754 VSS 0.00569f 
C7650 VCC.n3755 VSS 1.3e-19 
C7651 VCC.n3756 VSS 3.67e-19 
C7652 VCC.n3757 VSS 1.15e-19 
C7653 VCC.n3758 VSS 3.38e-19 
C7654 VCC.n3759 VSS 3.5e-20 
C7655 VCC.n3760 VSS 3.5e-20 
C7656 VCC.n3761 VSS 2.68e-20 
C7657 VCC.n3762 VSS 2.06e-20 
C7658 VCC.n3763 VSS 6.38e-20 
C7659 VCC.n3764 VSS 5.97e-20 
C7660 VCC.n3765 VSS 4.73e-20 
C7661 VCC.n3766 VSS 4.73e-20 
C7662 VCC.n3767 VSS 3.09e-20 
C7663 VCC.n3768 VSS 1.23e-20 
C7664 VCC.n3769 VSS 1.65e-20 
C7665 VCC.n3770 VSS 1.54e-19 
C7666 VCC.n3771 VSS 1.54e-19 
C7667 VCC.n3772 VSS 1.65e-20 
C7668 VCC.n3773 VSS 3.29e-20 
C7669 VCC.t182 VSS 1.67e-19 
C7670 VCC.n3774 VSS 0.00101f 
C7671 VCC.n3775 VSS 2.71e-19 
C7672 VCC.n3776 VSS 7.46e-19 
C7673 VCC.n3777 VSS 0.00333f 
C7674 VCC.n3778 VSS 2.46e-19 
C7675 VCC.n3779 VSS 3.02e-19 
C7676 VCC.n3780 VSS 3.7e-20 
C7677 VCC.n3781 VSS 5.15e-20 
C7678 VCC.n3782 VSS 5.97e-20 
C7679 VCC.n3783 VSS 6.38e-20 
C7680 VCC.n3784 VSS 4.73e-20 
C7681 VCC.n3785 VSS 4.73e-20 
C7682 VCC.n3786 VSS 2.68e-20 
C7683 VCC.n3787 VSS 3.29e-20 
C7684 VCC.n3788 VSS 1.65e-20 
C7685 VCC.n3789 VSS 1.54e-19 
C7686 VCC.n3790 VSS 1.54e-19 
C7687 VCC.n3791 VSS 1.65e-20 
C7688 VCC.n3792 VSS 3.09e-20 
C7689 VCC.n3793 VSS 3.09e-20 
C7690 VCC.n3794 VSS 4.73e-20 
C7691 VCC.n3795 VSS 4.32e-20 
C7692 VCC.n3796 VSS 3.5e-20 
C7693 VCC.n3797 VSS 3.5e-20 
C7694 VCC.n3798 VSS 1.35e-19 
C7695 VCC.n3799 VSS 5.24e-19 
C7696 VCC.n3800 VSS 1.4e-19 
C7697 VCC.n3801 VSS 5.4e-19 
C7698 VCC.n3802 VSS 1.35e-19 
C7699 VCC.n3803 VSS 4.37e-19 
C7700 VCC.n3804 VSS 1.13e-19 
C7701 VCC.n3805 VSS 8.23e-21 
C7702 VCC.n3806 VSS 1.65e-20 
C7703 VCC.n3807 VSS 3.5e-20 
C7704 VCC.n3808 VSS 3.91e-20 
C7705 VCC.n3809 VSS 3.09e-20 
C7706 VCC.n3810 VSS 1.85e-20 
C7707 VCC.n3811 VSS 3.5e-20 
C7708 VCC.n3812 VSS 1.05e-19 
C7709 VCC.n3813 VSS 2.06e-20 
C7710 VCC.n3814 VSS 2.26e-20 
C7711 VCC.n3815 VSS 3.7e-20 
C7712 VCC.n3816 VSS 5.15e-20 
C7713 VCC.n3817 VSS 1.38e-19 
C7714 VCC.n3818 VSS 1.17e-19 
C7715 VCC.n3819 VSS 4.32e-20 
C7716 VCC.n3820 VSS 2.88e-20 
C7717 VCC.n3821 VSS 2.68e-20 
C7718 VCC.n3822 VSS 6.59e-20 
C7719 VCC.n3823 VSS 5.56e-20 
C7720 VCC.n3824 VSS 2.68e-20 
C7721 VCC.n3825 VSS 4.32e-20 
C7722 VCC.n3826 VSS 1.05e-19 
C7723 VCC.n3827 VSS 3.09e-20 
C7724 VCC.n3828 VSS 3.7e-20 
C7725 VCC.n3829 VSS 4.32e-20 
C7726 VCC.n3830 VSS 1.05e-19 
C7727 VCC.n3831 VSS 4.53e-20 
C7728 VCC.n3832 VSS 4.53e-20 
C7729 VCC.n3833 VSS 7.82e-20 
C7730 VCC.n3834 VSS 2.18e-19 
C7731 VCC.n3835 VSS 1.4e-19 
C7732 VCC.n3836 VSS 1.4e-19 
C7733 VCC.n3837 VSS 5.4e-19 
C7734 VCC.n3838 VSS 1.35e-19 
C7735 VCC.t274 VSS 4.21e-19 
C7736 VCC.n3839 VSS 3.33e-19 
C7737 VCC.n3840 VSS 1.13e-19 
C7738 VCC.n3841 VSS 8.23e-21 
C7739 VCC.n3842 VSS 1.65e-20 
C7740 VCC.n3843 VSS 3.5e-20 
C7741 VCC.n3844 VSS 3.5e-20 
C7742 VCC.n3845 VSS 3.5e-20 
C7743 VCC.n3846 VSS 1.17e-19 
C7744 VCC.n3847 VSS 1.38e-19 
C7745 VCC.n3848 VSS 5.15e-20 
C7746 VCC.n3849 VSS 4.73e-20 
C7747 VCC.n3850 VSS 7.2e-20 
C7748 VCC.n3851 VSS 2.68e-20 
C7749 VCC.n3852 VSS 1.65e-20 
C7750 VCC.n3853 VSS 1.54e-19 
C7751 VCC.n3854 VSS 1.54e-19 
C7752 VCC.n3855 VSS 1.65e-20 
C7753 VCC.n3856 VSS 2.47e-20 
C7754 VCC.n3857 VSS 1.23e-20 
C7755 VCC.n3858 VSS 7.62e-19 
C7756 VCC.n3859 VSS 4.12e-20 
C7757 VCC.n3860 VSS 5.15e-20 
C7758 VCC.n3861 VSS 6.59e-20 
C7759 VCC.n3862 VSS 5.76e-20 
C7760 VCC.n3863 VSS 4.73e-20 
C7761 VCC.n3864 VSS 2.26e-20 
C7762 VCC.n3865 VSS 2.68e-20 
C7763 VCC.n3866 VSS 1.03e-20 
C7764 VCC.n3867 VSS 3.5e-20 
C7765 VCC.n3868 VSS 3.5e-20 
C7766 VCC.n3869 VSS 1.35e-19 
C7767 VCC.n3870 VSS 4.53e-19 
C7768 VCC.n3871 VSS 7.71e-19 
C7769 VCC.n3872 VSS 1.32e-19 
C7770 VCC.n3873 VSS 3.5e-20 
C7771 VCC.n3874 VSS 3.42e-20 
C7772 VCC.n3875 VSS 2.36e-19 
C7773 VCC.n3876 VSS 3.21e-19 
C7774 VCC.n3877 VSS 2.61e-19 
C7775 VCC.n3878 VSS 0.00189f 
C7776 VCC.n3879 VSS 2.68e-19 
C7777 VCC.n3880 VSS 0.00246f 
C7778 VCC.n3881 VSS 5.76e-20 
C7779 VCC.n3882 VSS 2.88e-20 
C7780 VCC.n3883 VSS 3.5e-20 
C7781 VCC.n3884 VSS 3.42e-20 
C7782 VCC.n3885 VSS 3.5e-20 
C7783 VCC.n3886 VSS 4.53e-19 
C7784 VCC.n3887 VSS 1.17e-19 
C7785 VCC.n3888 VSS 3.5e-20 
C7786 VCC.n3889 VSS 1.44e-20 
C7787 VCC.n3890 VSS 4.12e-20 
C7788 VCC.n3891 VSS 5.76e-20 
C7789 VCC.n3892 VSS 5.76e-20 
C7790 VCC.n3893 VSS 2.06e-20 
C7791 VCC.n3894 VSS 3.29e-20 
C7792 VCC.n3895 VSS 7.2e-20 
C7793 VCC.n3896 VSS 3.29e-20 
C7794 VCC.n3897 VSS 4.73e-20 
C7795 VCC.n3898 VSS 2.26e-20 
C7796 VCC.n3899 VSS 1.01e-19 
C7797 VCC.n3900 VSS 1.36e-19 
C7798 VCC.n3901 VSS 1.35e-19 
C7799 VCC.n3902 VSS 3.5e-20 
C7800 VCC.n3903 VSS 3.5e-20 
C7801 VCC.n3904 VSS 3.5e-20 
C7802 VCC.n3905 VSS 3.5e-20 
C7803 VCC.n3906 VSS 3.09e-20 
C7804 VCC.n3907 VSS 3.91e-20 
C7805 VCC.n3908 VSS 4.73e-20 
C7806 VCC.n3909 VSS 4.32e-20 
C7807 VCC.n3910 VSS 2.68e-20 
C7808 VCC.n3911 VSS 4.53e-20 
C7809 VCC.n3912 VSS 4.53e-20 
C7810 VCC.n3913 VSS 3.09e-20 
C7811 VCC.n3914 VSS 4.32e-20 
C7812 VCC.n3915 VSS 2.68e-20 
C7813 VCC.n3916 VSS 7.82e-20 
C7814 VCC.n3917 VSS 5.56e-20 
C7815 VCC.n3918 VSS 1.4e-19 
C7816 VCC.n3919 VSS 2.18e-19 
C7817 VCC.n3920 VSS 1.35e-19 
C7818 VCC.n3921 VSS 1.13e-19 
C7819 VCC.n3922 VSS 3.5e-20 
C7820 VCC.n3923 VSS 1.85e-20 
C7821 VCC.n3924 VSS 3.7e-20 
C7822 VCC.n3925 VSS 3.09e-20 
C7823 VCC.n3926 VSS 6.59e-20 
C7824 VCC.n3927 VSS 2.68e-20 
C7825 VCC.n3928 VSS 5.76e-20 
C7826 VCC.n3929 VSS 4.73e-20 
C7827 VCC.n3930 VSS 3.5e-20 
C7828 VCC.t301 VSS 1.56e-19 
C7829 VCC.n3931 VSS 7.97e-19 
C7830 VCC.n3932 VSS 3.09e-20 
C7831 VCC.n3933 VSS 3.5e-20 
C7832 VCC.n3934 VSS 3.5e-20 
C7833 VCC.t300 VSS 4.21e-19 
C7834 VCC.n3935 VSS 1.32e-19 
C7835 VCC.n3936 VSS 1.09e-19 
C7836 VCC.n3937 VSS 3.5e-20 
C7837 VCC.n3938 VSS 3.09e-20 
C7838 VCC.n3939 VSS 5.97e-20 
C7839 VCC.n3940 VSS 2.26e-20 
C7840 VCC.n3941 VSS 5.76e-20 
C7841 VCC.n3942 VSS 2.68e-20 
C7842 VCC.n3943 VSS 2.68e-20 
C7843 VCC.n3944 VSS 1.9e-19 
C7844 VCC.n3945 VSS 5.76e-20 
C7845 VCC.n3946 VSS 2.68e-20 
C7846 VCC.n3947 VSS 2.68e-20 
C7847 VCC.n3948 VSS 2.68e-20 
C7848 VCC.n3949 VSS 5.76e-20 
C7849 VCC.n3950 VSS 2.26e-20 
C7850 VCC.n3951 VSS 3.09e-20 
C7851 VCC.n3952 VSS 2.26e-20 
C7852 VCC.n3953 VSS 5.15e-20 
C7853 VCC.n3954 VSS 4.73e-20 
C7854 VCC.n3955 VSS 3.7e-20 
C7855 VCC.n3956 VSS 3.5e-20 
C7856 VCC.n3957 VSS 7.41e-20 
C7857 VCC.n3958 VSS 1.91e-19 
C7858 VCC.n3959 VSS 9.88e-20 
C7859 VCC.n3960 VSS 3e-20 
C7860 VCC.n3961 VSS 5.12e-19 
C7861 VCC.n3962 VSS 1.18e-19 
C7862 VCC.n3963 VSS 3.5e-20 
C7863 VCC.n3964 VSS 3.5e-20 
C7864 VCC.n3965 VSS 5.15e-20 
C7865 VCC.n3966 VSS 4.32e-20 
C7866 VCC.n3967 VSS 2.68e-20 
C7867 VCC.n3968 VSS 3.91e-20 
C7868 VCC.n3969 VSS 1.44e-20 
C7869 VCC.n3970 VSS 3.5e-20 
C7870 VCC.n3971 VSS 3e-20 
C7871 VCC.n3972 VSS 7.95e-19 
C7872 VCC.n3973 VSS 1.83e-19 
C7873 VCC.n3974 VSS 2.88e-20 
C7874 VCC.n3975 VSS 2.68e-20 
C7875 VCC.n3976 VSS 2.68e-20 
C7876 VCC.n3977 VSS 2.68e-20 
C7877 VCC.n3978 VSS 4.53e-20 
C7878 VCC.n3979 VSS 3.7e-20 
C7879 VCC.n3980 VSS 7.82e-20 
C7880 VCC.n3981 VSS 1.17e-19 
C7881 VCC.n3982 VSS 3.91e-20 
C7882 VCC.n3983 VSS 1.65e-20 
C7883 VCC.n3984 VSS 2.68e-20 
C7884 VCC.n3985 VSS 3.5e-20 
C7885 VCC.n3986 VSS 3e-20 
C7886 VCC.n3987 VSS 5.12e-19 
C7887 VCC.n3988 VSS 1.18e-19 
C7888 VCC.n3989 VSS 3.5e-20 
C7889 VCC.n3990 VSS 3.5e-20 
C7890 VCC.t203 VSS 1.55e-19 
C7891 VCC.n3991 VSS 7.57e-19 
C7892 VCC.n3992 VSS 4.73e-20 
C7893 VCC.n3993 VSS 1.54e-19 
C7894 VCC.n3994 VSS 2.88e-20 
C7895 VCC.n3995 VSS 2.88e-20 
C7896 VCC.n3996 VSS 3.5e-20 
C7897 VCC.n3997 VSS 5.76e-20 
C7898 VCC.n3998 VSS 9.88e-20 
C7899 VCC.n3999 VSS 1.3e-19 
C7900 VCC.n4000 VSS 3e-20 
C7901 VCC.t201 VSS 0.005f 
C7902 VCC.t122 VSS 0.00453f 
C7903 VCC.n4001 VSS 0.00229f 
C7904 VCC.n4002 VSS 1.91e-19 
C7905 VCC.n4003 VSS 3.5e-20 
C7906 VCC.n4004 VSS 3.14e-19 
C7907 VCC.n4005 VSS 2.47e-20 
C7908 VCC.n4006 VSS 5.76e-20 
C7909 VCC.n4007 VSS 2.47e-20 
C7910 VCC.n4008 VSS 8.23e-21 
C7911 VCC.n4009 VSS 2.88e-20 
C7912 VCC.n4010 VSS 5.76e-20 
C7913 VCC.n4011 VSS 2.47e-20 
C7914 VCC.n4012 VSS 2.88e-20 
C7915 VCC.n4013 VSS 2.47e-20 
C7916 VCC.n4014 VSS 5.15e-20 
C7917 VCC.n4015 VSS 4.73e-20 
C7918 VCC.n4016 VSS 3.7e-20 
C7919 VCC.n4017 VSS 3.5e-20 
C7920 VCC.n4018 VSS 7.41e-20 
C7921 VCC.t298 VSS 6.42e-19 
C7922 VCC.n4019 VSS 3e-20 
C7923 VCC.n4020 VSS 5.97e-20 
C7924 VCC.n4021 VSS 4.13e-19 
C7925 VCC.n4022 VSS 9.53e-20 
C7926 VCC.n4023 VSS 3.5e-20 
C7927 VCC.n4024 VSS 3.5e-20 
C7928 VCC.n4025 VSS 5.35e-20 
C7929 VCC.n4026 VSS 4.32e-20 
C7930 VCC.n4027 VSS 2.68e-20 
C7931 VCC.n4028 VSS 3.7e-20 
C7932 VCC.n4029 VSS 1.65e-20 
C7933 VCC.n4030 VSS 4.53e-20 
C7934 VCC.n4031 VSS 1.2e-19 
C7935 VCC.n4032 VSS 5.2e-19 
C7936 VCC.n4033 VSS 1.2e-19 
C7937 VCC.n4034 VSS 6.38e-20 
C7938 VCC.n4035 VSS 2.47e-20 
C7939 VCC.n4036 VSS 4.53e-20 
C7940 VCC.n4037 VSS 3.5e-20 
C7941 VCC.n4038 VSS 3.5e-20 
C7942 VCC.n4039 VSS 2.68e-20 
C7943 VCC.n4040 VSS 2.68e-20 
C7944 VCC.n4041 VSS 2.47e-20 
C7945 VCC.n4042 VSS 4.53e-20 
C7946 VCC.n4043 VSS 2.68e-20 
C7947 VCC.n4044 VSS 4.32e-20 
C7948 VCC.n4045 VSS 2.68e-20 
C7949 VCC.n4046 VSS 3.91e-20 
C7950 VCC.n4047 VSS 2.88e-20 
C7951 VCC.n4048 VSS 4.73e-20 
C7952 VCC.n4049 VSS 3.7e-20 
C7953 VCC.n4050 VSS 3.7e-20 
C7954 VCC.n4051 VSS 3.5e-20 
C7955 VCC.n4052 VSS 5.76e-20 
C7956 VCC.n4053 VSS 4.73e-20 
C7957 VCC.n4054 VSS 3.09e-20 
C7958 VCC.n4055 VSS 3.5e-20 
C7959 VCC.n4056 VSS 3.5e-20 
C7960 VCC.n4057 VSS 3.5e-20 
C7961 VCC.n4058 VSS 1.18e-19 
C7962 VCC.n4059 VSS 3e-20 
C7963 VCC.n4060 VSS 1.15e-19 
C7964 VCC.n4061 VSS 9.88e-20 
C7965 VCC.n4062 VSS 5.76e-20 
C7966 VCC.n4063 VSS 3.5e-20 
C7967 VCC.n4064 VSS 3.09e-20 
C7968 VCC.n4065 VSS 3.09e-20 
C7969 VCC.n4066 VSS 2.26e-20 
C7970 VCC.n4067 VSS 5.76e-20 
C7971 VCC.n4068 VSS 2.68e-20 
C7972 VCC.n4069 VSS 2.68e-20 
C7973 VCC.n4070 VSS 0.00185f 
C7974 VCC.n4071 VSS 2.72e-19 
C7975 VCC.n4072 VSS 2.26e-20 
C7976 VCC.n4073 VSS 1.87e-19 
C7977 VCC.n4074 VSS 3.5e-20 
C7978 VCC.n4075 VSS 2.68e-20 
C7979 VCC.n4076 VSS 5.97e-20 
C7980 VCC.n4077 VSS 4.73e-20 
C7981 VCC.n4078 VSS 4.73e-20 
C7982 VCC.n4079 VSS 5.15e-20 
C7983 VCC.n4080 VSS 7.41e-20 
C7984 VCC.n4081 VSS 3.7e-20 
C7985 VCC.n4082 VSS 2.26e-20 
C7986 VCC.n4083 VSS 6.38e-20 
C7987 VCC.n4084 VSS 4.73e-20 
C7988 VCC.n4085 VSS 3.29e-20 
C7989 VCC.n4086 VSS 3.5e-20 
C7990 VCC.n4087 VSS 3e-20 
C7991 VCC.t75 VSS 0.005f 
C7992 VCC.t204 VSS 0.00453f 
C7993 VCC.n4088 VSS 0.00228f 
C7994 VCC.n4089 VSS 1.3e-19 
C7995 VCC.t73 VSS 4.05e-19 
C7996 VCC.n4090 VSS 4.05e-19 
C7997 VCC.n4091 VSS 1.15e-19 
C7998 VCC.n4092 VSS 3.36e-19 
C7999 VCC.n4093 VSS 6.17e-21 
C8000 VCC.n4094 VSS 3.12e-19 
C8001 VCC.n4095 VSS 1.65e-20 
C8002 VCC.n4096 VSS 1.54e-19 
C8003 VCC.n4097 VSS 1.54e-19 
C8004 VCC.n4098 VSS 1.65e-20 
C8005 VCC.n4099 VSS 1.03e-20 
C8006 VCC.n4100 VSS 3.5e-20 
C8007 VCC.n4101 VSS 2.26e-20 
C8008 VCC.n4102 VSS 4.73e-20 
C8009 VCC.n4103 VSS 3.5e-20 
C8010 VCC.n4104 VSS 3e-20 
C8011 VCC.n4105 VSS 1.3e-19 
C8012 VCC.n4106 VSS 5.12e-19 
C8013 VCC.n4107 VSS 1.3e-19 
C8014 VCC.n4108 VSS 4.13e-19 
C8015 VCC.n4109 VSS 9.53e-20 
C8016 VCC.n4110 VSS 5.76e-20 
C8017 VCC.n4111 VSS 7.41e-20 
C8018 VCC.n4112 VSS 5.56e-20 
C8019 VCC.t74 VSS 1.55e-19 
C8020 VCC.n4113 VSS 3.91e-20 
C8021 VCC.n4114 VSS 3.91e-20 
C8022 VCC.n4115 VSS 1.85e-20 
C8023 VCC.n4116 VSS 7.55e-19 
C8024 VCC.n4117 VSS 4.94e-20 
C8025 VCC.n4118 VSS 5.15e-20 
C8026 VCC.n4119 VSS 7.2e-20 
C8027 VCC.n4120 VSS 1.38e-19 
C8028 VCC.n4121 VSS 1.17e-19 
C8029 VCC.n4122 VSS 4.32e-20 
C8030 VCC.n4123 VSS 2.88e-20 
C8031 VCC.n4124 VSS 2.68e-20 
C8032 VCC.n4125 VSS 3.5e-20 
C8033 VCC.n4126 VSS 3.5e-20 
C8034 VCC.n4127 VSS 2.88e-20 
C8035 VCC.n4128 VSS 2.68e-20 
C8036 VCC.n4129 VSS 2.68e-20 
C8037 VCC.n4130 VSS 2.68e-20 
C8038 VCC.n4131 VSS 4.12e-20 
C8039 VCC.n4132 VSS 4.12e-20 
C8040 VCC.n4133 VSS 3.91e-20 
C8041 VCC.n4134 VSS 4.53e-20 
C8042 VCC.n4135 VSS 4.53e-20 
C8043 VCC.n4136 VSS 1.05e-19 
C8044 VCC.n4137 VSS 1.05e-19 
C8045 VCC.n4138 VSS 4.32e-20 
C8046 VCC.n4139 VSS 3.7e-20 
C8047 VCC.n4140 VSS 2.68e-20 
C8048 VCC.n4141 VSS 2.68e-20 
C8049 VCC.n4142 VSS 6.79e-20 
C8050 VCC.n4143 VSS 9.26e-20 
C8051 VCC.n4144 VSS 1.83e-19 
C8052 VCC.n4145 VSS 7.95e-19 
C8053 VCC.n4146 VSS 5.2e-19 
C8054 VCC.n4147 VSS 1.3e-19 
C8055 VCC.n4148 VSS 3e-20 
C8056 VCC.n4149 VSS 3.5e-20 
C8057 VCC.n4150 VSS 5.97e-20 
C8058 VCC.n4151 VSS 7.41e-20 
C8059 VCC.n4152 VSS 5.15e-20 
C8060 VCC.n4153 VSS 5.15e-20 
C8061 VCC.n4154 VSS 3.09e-20 
C8062 VCC.n4155 VSS 3.09e-20 
C8063 VCC.n4156 VSS 3.7e-20 
C8064 VCC.n4157 VSS 2.68e-20 
C8065 VCC.n4158 VSS 3.91e-20 
C8066 VCC.n4159 VSS 1.17e-19 
C8067 VCC.n4160 VSS 1.38e-19 
C8068 VCC.n4161 VSS 7e-20 
C8069 VCC.n4162 VSS 4.73e-20 
C8070 VCC.n4163 VSS 3.5e-20 
C8071 VCC.n4164 VSS 3.5e-20 
C8072 VCC.n4165 VSS 3.5e-20 
C8073 VCC.n4166 VSS 4.53e-20 
C8074 VCC.n4167 VSS 1.18e-19 
C8075 VCC.n4168 VSS 5.12e-19 
C8076 VCC.n4169 VSS 1.3e-19 
C8077 VCC.n4170 VSS 1.61e-19 
C8078 VCC.n4171 VSS 9.9e-20 
C8079 VCC.n4172 VSS 0.00243f 
C8080 VCC.n4173 VSS 2.26e-20 
C8081 VCC.n4174 VSS 4.13e-19 
C8082 VCC.n4175 VSS 3.5e-20 
C8083 VCC.n4176 VSS 3.5e-20 
C8084 VCC.n4177 VSS 2.47e-20 
C8085 VCC.n4178 VSS 2.06e-20 
C8086 VCC.n4179 VSS 6.17e-20 
C8087 VCC.n4180 VSS 6.17e-20 
C8088 VCC.n4181 VSS 4.73e-20 
C8089 VCC.n4182 VSS 4.73e-20 
C8090 VCC.n4183 VSS 2.88e-20 
C8091 VCC.n4184 VSS 1.44e-20 
C8092 VCC.n4185 VSS 1.65e-20 
C8093 VCC.n4186 VSS 1.54e-19 
C8094 VCC.n4187 VSS 1.54e-19 
C8095 VCC.n4188 VSS 1.65e-20 
C8096 VCC.n4189 VSS 3.09e-20 
C8097 VCC.t299 VSS 1.55e-19 
C8098 VCC.n4190 VSS 0.00102f 
C8099 VCC.n4191 VSS 2.73e-19 
C8100 VCC.n4192 VSS 0.00136f 
C8101 VCC.n4193 VSS 2.73e-19 
C8102 VCC.n4194 VSS 0.00181f 
C8103 VCC.n4195 VSS 5.76e-20 
C8104 VCC.n4196 VSS 1.54e-19 
C8105 VCC.n4197 VSS 1.65e-20 
C8106 VCC.n4198 VSS 2.88e-20 
C8107 VCC.n4199 VSS 2.47e-20 
C8108 VCC.n4200 VSS 6.17e-20 
C8109 VCC.n4201 VSS 4.73e-20 
C8110 VCC.n4202 VSS 4.73e-20 
C8111 VCC.n4203 VSS 5.15e-20 
C8112 VCC.n4204 VSS 3.5e-20 
C8113 VCC.n4205 VSS 7.41e-20 
C8114 VCC.n4206 VSS 3.7e-20 
C8115 VCC.n4207 VSS 2.26e-20 
C8116 VCC.n4208 VSS 6.17e-20 
C8117 VCC.n4209 VSS 4.73e-20 
C8118 VCC.n4210 VSS 3.5e-20 
C8119 VCC.n4211 VSS 2.88e-20 
C8120 VCC.n4212 VSS 3.4e-19 
C8121 VCC.n4213 VSS 1.15e-19 
C8122 VCC.n4214 VSS 3.98e-19 
C8123 VCC.t202 VSS 4.05e-19 
C8124 VCC.n4215 VSS 1.22e-19 
C8125 VCC.n4216 VSS 1.3e-19 
C8126 VCC.n4217 VSS 3e-20 
C8127 VCC.n4218 VSS 3.5e-20 
C8128 VCC.n4219 VSS 3.5e-20 
C8129 VCC.n4220 VSS 4.73e-20 
C8130 VCC.n4221 VSS 2.47e-20 
C8131 VCC.n4222 VSS 1.23e-20 
C8132 VCC.n4223 VSS 1.65e-20 
C8133 VCC.n4224 VSS 2.47e-20 
C8134 VCC.n4225 VSS 5.76e-20 
C8135 VCC.n4226 VSS 1.38e-19 
C8136 VCC.n4227 VSS 7e-20 
C8137 VCC.n4228 VSS 3.7e-20 
C8138 VCC.n4229 VSS 2.47e-20 
C8139 VCC.n4230 VSS 3.7e-20 
C8140 VCC.n4231 VSS 1.85e-20 
C8141 VCC.n4232 VSS 3.09e-20 
C8142 VCC.n4233 VSS 5.35e-20 
C8143 VCC.n4234 VSS 4.73e-20 
C8144 VCC.n4235 VSS 5.35e-20 
C8145 VCC.n4236 VSS 7.41e-20 
C8146 VCC.n4237 VSS 5.76e-20 
C8147 VCC.n4238 VSS 9.53e-20 
C8148 VCC.n4239 VSS 4.13e-19 
C8149 VCC.n4240 VSS 1.3e-19 
C8150 VCC.n4241 VSS 5.2e-19 
C8151 VCC.n4242 VSS 1.2e-19 
C8152 VCC.n4243 VSS 4.73e-20 
C8153 VCC.n4244 VSS 2.68e-20 
C8154 VCC.n4245 VSS 3.5e-20 
C8155 VCC.n4246 VSS 3.5e-20 
C8156 VCC.n4247 VSS 2.68e-20 
C8157 VCC.n4248 VSS 2.68e-20 
C8158 VCC.n4249 VSS 4.32e-20 
C8159 VCC.n4250 VSS 4.32e-20 
C8160 VCC.n4251 VSS 4.32e-20 
C8161 VCC.n4252 VSS 2.88e-20 
C8162 VCC.n4253 VSS 3.5e-20 
C8163 VCC.n4254 VSS 2.68e-20 
C8164 VCC.n4255 VSS 7.82e-20 
C8165 VCC.n4256 VSS 4.73e-20 
C8166 VCC.n4257 VSS 4.73e-20 
C8167 VCC.n4258 VSS 1.05e-19 
C8168 VCC.n4259 VSS 1.05e-19 
C8169 VCC.n4260 VSS 4.53e-20 
C8170 VCC.n4261 VSS 2.68e-20 
C8171 VCC.n4262 VSS 2.68e-20 
C8172 VCC.n4263 VSS 6.59e-20 
C8173 VCC.n4264 VSS 9.26e-20 
C8174 VCC.n4265 VSS 6.59e-20 
C8175 VCC.n4266 VSS 2.47e-20 
C8176 VCC.n4267 VSS 2.47e-20 
C8177 VCC.n4268 VSS 2.88e-20 
C8178 VCC.n4269 VSS 3.5e-20 
C8179 VCC.n4270 VSS 3.5e-20 
C8180 VCC.n4271 VSS 4.53e-20 
C8181 VCC.n4272 VSS 1.2e-19 
C8182 VCC.n4273 VSS 5.2e-19 
C8183 VCC.n4274 VSS 1.3e-19 
C8184 VCC.n4275 VSS 4.13e-19 
C8185 VCC.n4276 VSS 9.53e-20 
C8186 VCC.n4277 VSS 5.97e-20 
C8187 VCC.n4278 VSS 7.41e-20 
C8188 VCC.n4279 VSS 5.35e-20 
C8189 VCC.n4280 VSS 5.15e-20 
C8190 VCC.n4281 VSS 3.09e-20 
C8191 VCC.n4282 VSS 3.09e-20 
C8192 VCC.n4283 VSS 3.91e-20 
C8193 VCC.n4284 VSS 2.47e-20 
C8194 VCC.n4285 VSS 3.7e-20 
C8195 VCC.n4286 VSS 1.17e-19 
C8196 VCC.n4287 VSS 1.38e-19 
C8197 VCC.n4288 VSS 7.2e-20 
C8198 VCC.n4289 VSS 4.73e-20 
C8199 VCC.n4290 VSS 3.5e-20 
C8200 VCC.n4291 VSS 3.5e-20 
C8201 VCC.n4292 VSS 4.53e-20 
C8202 VCC.n4293 VSS 5.97e-20 
C8203 VCC.n4294 VSS 3.5e-20 
C8204 VCC.n4295 VSS 3e-20 
C8205 VCC.n4296 VSS 1.3e-19 
C8206 VCC.n4297 VSS 1.53e-19 
C8207 VCC.t91 VSS 4.05e-19 
C8208 VCC.n4298 VSS 2.06e-19 
C8209 VCC.n4299 VSS 1.35e-19 
C8210 VCC.n4300 VSS 9.67e-20 
C8211 VCC.n4301 VSS 3.35e-20 
C8212 VCC.n4302 VSS 3.5e-20 
C8213 VCC.n4303 VSS 2.36e-19 
C8214 VCC.n4304 VSS 0.0023f 
C8215 VCC.t303 VSS 0.0031f 
C8216 VCC.t266 VSS 0.00366f 
C8217 VCC.t302 VSS 0.00365f 
C8218 VCC.t267 VSS 0.00386f 
C8219 VCC.n4305 VSS 0.00569f 
C8220 VCC.n4306 VSS 1.3e-19 
C8221 VCC.n4307 VSS 3.67e-19 
C8222 VCC.n4308 VSS 1.15e-19 
C8223 VCC.n4309 VSS 3.38e-19 
C8224 VCC.n4310 VSS 3.5e-20 
C8225 VCC.n4311 VSS 3.5e-20 
C8226 VCC.n4312 VSS 2.68e-20 
C8227 VCC.n4313 VSS 2.06e-20 
C8228 VCC.n4314 VSS 6.38e-20 
C8229 VCC.n4315 VSS 5.97e-20 
C8230 VCC.n4316 VSS 4.73e-20 
C8231 VCC.n4317 VSS 4.73e-20 
C8232 VCC.n4318 VSS 3.09e-20 
C8233 VCC.n4319 VSS 1.23e-20 
C8234 VCC.n4320 VSS 1.65e-20 
C8235 VCC.n4321 VSS 1.54e-19 
C8236 VCC.n4322 VSS 1.54e-19 
C8237 VCC.n4323 VSS 1.65e-20 
C8238 VCC.n4324 VSS 3.29e-20 
C8239 VCC.t92 VSS 1.67e-19 
C8240 VCC.n4325 VSS 0.00101f 
C8241 VCC.n4326 VSS 2.71e-19 
C8242 VCC.n4327 VSS 7.46e-19 
C8243 VCC.n4328 VSS 0.00333f 
C8244 VCC.n4329 VSS 2.46e-19 
C8245 VCC.n4330 VSS 3.02e-19 
C8246 VCC.n4331 VSS 3.7e-20 
C8247 VCC.n4332 VSS 5.15e-20 
C8248 VCC.n4333 VSS 6.38e-20 
C8249 VCC.n4334 VSS 4.73e-20 
C8250 VCC.n4335 VSS 4.73e-20 
C8251 VCC.n4336 VSS 2.68e-20 
C8252 VCC.n4337 VSS 3.29e-20 
C8253 VCC.n4338 VSS 1.65e-20 
C8254 VCC.n4339 VSS 1.54e-19 
C8255 VCC.n4340 VSS 1.54e-19 
C8256 VCC.n4341 VSS 5.56e-20 
C8257 VCC.n4342 VSS 2.88e-20 
C8258 VCC.n4343 VSS 1.65e-20 
C8259 VCC.n4344 VSS 3.09e-20 
C8260 VCC.n4345 VSS 4.73e-20 
C8261 VCC.n4346 VSS 4.73e-20 
C8262 VCC.n4347 VSS 4.32e-20 
C8263 VCC.n4348 VSS 1.17e-19 
C8264 VCC.n4349 VSS 3.33e-19 
C8265 VCC.n4350 VSS 1.35e-19 
C8266 VCC.n4351 VSS 4.37e-19 
C8267 VCC.n4352 VSS 5.24e-19 
C8268 VCC.n4353 VSS 1.36e-19 
C8269 VCC.n4354 VSS 1.01e-19 
C8270 VCC.n4355 VSS 1.05e-19 
C8271 VCC.n4356 VSS 2.06e-20 
C8272 VCC.n4357 VSS 2.26e-20 
C8273 VCC.n4358 VSS 3.7e-20 
C8274 VCC.n4359 VSS 5.15e-20 
C8275 VCC.n4360 VSS 1.38e-19 
C8276 VCC.n4361 VSS 3.91e-20 
C8277 VCC.n4362 VSS 2.88e-20 
C8278 VCC.n4363 VSS 4.32e-20 
C8279 VCC.n4364 VSS 1.17e-19 
C8280 VCC.n4365 VSS 3.7e-20 
C8281 VCC.n4366 VSS 3.91e-20 
C8282 VCC.n4367 VSS 3.5e-20 
C8283 VCC.n4368 VSS 1.65e-20 
C8284 VCC.n4369 VSS 8.23e-21 
C8285 VCC.n4370 VSS 3.5e-20 
C8286 VCC.n4371 VSS 3.5e-20 
C8287 VCC.n4372 VSS 1.4e-19 
C8288 VCC.n4373 VSS 5.4e-19 
C8289 VCC.n4374 VSS 8.42e-19 
C8290 VCC.n4375 VSS 5.4e-19 
C8291 VCC.n4376 VSS 1.4e-19 
C8292 VCC.n4377 VSS 1.4e-19 
C8293 VCC.n4378 VSS 2.18e-19 
C8294 VCC.n4379 VSS 7.82e-20 
C8295 VCC.n4380 VSS 4.32e-20 
C8296 VCC.n4381 VSS 4.32e-20 
C8297 VCC.n4382 VSS 1.05e-19 
C8298 VCC.n4383 VSS 1.05e-19 
C8299 VCC.n4384 VSS 4.32e-20 
C8300 VCC.n4385 VSS 3.7e-20 
C8301 VCC.n4386 VSS 2.68e-20 
C8302 VCC.n4387 VSS 5.76e-20 
C8303 VCC.n4388 VSS 6.38e-20 
C8304 VCC.n4389 VSS 3.5e-20 
C8305 VCC.n4390 VSS 3.5e-20 
C8306 VCC.n4391 VSS 1.17e-19 
C8307 VCC.n4392 VSS 1.38e-19 
C8308 VCC.n4393 VSS 5.15e-20 
C8309 VCC.n4394 VSS 1.05e-19 
C8310 VCC.n4395 VSS 2.26e-20 
C8311 VCC.n4396 VSS 5.76e-20 
C8312 VCC.n4397 VSS 3.7e-20 
C8313 VCC.n4398 VSS 3.7e-20 
C8314 VCC.n4399 VSS 3.09e-20 
C8315 VCC.n4400 VSS 1.85e-20 
C8316 VCC.n4401 VSS 1.65e-20 
C8317 VCC.n4402 VSS 8.23e-21 
C8318 VCC.n4403 VSS 1.13e-19 
C8319 VCC.n4404 VSS 3.33e-19 
C8320 VCC.t99 VSS 4.21e-19 
C8321 VCC.n4405 VSS 2.06e-19 
C8322 VCC.n4406 VSS 1.35e-19 
C8323 VCC.n4407 VSS 3.5e-20 
C8324 VCC.n4408 VSS 3.5e-20 
C8325 VCC.n4409 VSS 3.5e-20 
C8326 VCC.n4410 VSS 1.03e-20 
C8327 VCC.n4411 VSS 2.68e-20 
C8328 VCC.n4412 VSS 3.09e-20 
C8329 VCC.n4413 VSS 2.68e-20 
C8330 VCC.n4414 VSS 1.65e-20 
C8331 VCC.n4415 VSS 1.54e-19 
C8332 VCC.n4416 VSS 1.54e-19 
C8333 VCC.n4417 VSS 1.65e-20 
C8334 VCC.t100 VSS 1.56e-19 
C8335 VCC.n4418 VSS 7.62e-19 
C8336 VCC.n4419 VSS 1.23e-20 
C8337 VCC.n4420 VSS 2.47e-20 
C8338 VCC.n4421 VSS 4.73e-20 
C8339 VCC.n4422 VSS 6.59e-20 
C8340 VCC.n4423 VSS 5.15e-20 
C8341 VCC.n4424 VSS 2.47e-20 
C8342 VCC.n4425 VSS 7.41e-20 
C8343 VCC.n4426 VSS 9.47e-20 
C8344 VCC.n4427 VSS 1.32e-19 
C8345 VCC.n4428 VSS 7.71e-19 
C8346 VCC.n4429 VSS 9.83e-19 
C8347 VCC.n4430 VSS 2.36e-19 
C8348 VCC.n4431 VSS 3.21e-19 
C8349 VCC.n4432 VSS 2.61e-19 
C8350 VCC.n4433 VSS 0.00189f 
C8351 VCC.n4434 VSS 0.00259f 
C8352 VCC.n4435 VSS 5.76e-20 
C8353 VCC.n4436 VSS 2.88e-20 
C8354 VCC.n4437 VSS 3.5e-20 
C8355 VCC.n4438 VSS 9.83e-19 
C8356 VCC.n4439 VSS 9.47e-20 
C8357 VCC.n4440 VSS 1.17e-19 
C8358 VCC.n4441 VSS 2.06e-19 
C8359 VCC.n4442 VSS 1.36e-19 
C8360 VCC.n4443 VSS 1.01e-19 
C8361 VCC.n4444 VSS 3.5e-20 
C8362 VCC.n4445 VSS 3.09e-20 
C8363 VCC.n4446 VSS 3.29e-20 
C8364 VCC.n4447 VSS 3.29e-20 
C8365 VCC.n4448 VSS 4.73e-20 
C8366 VCC.n4449 VSS 1.44e-20 
C8367 VCC.n4450 VSS 3.5e-20 
C8368 VCC.n4451 VSS 7.41e-20 
C8369 VCC.n4452 VSS 2.47e-20 
C8370 VCC.t265 VSS 1.56e-19 
C8371 VCC.n4453 VSS 5.76e-20 
C8372 VCC.n4454 VSS 2.06e-20 
C8373 VCC.n4455 VSS 5.76e-20 
C8374 VCC.n4456 VSS 3.7e-20 
C8375 VCC.n4457 VSS 4.32e-20 
C8376 VCC.n4458 VSS 2.68e-20 
C8377 VCC.n4459 VSS 3.91e-20 
C8378 VCC.n4460 VSS 6.38e-20 
C8379 VCC.n4461 VSS 1.85e-20 
C8380 VCC.n4462 VSS 3.5e-20 
C8381 VCC.n4463 VSS 3.09e-20 
C8382 VCC.n4464 VSS 3.7e-20 
C8383 VCC.n4465 VSS 3.09e-20 
C8384 VCC.n4466 VSS 2.26e-20 
C8385 VCC.n4467 VSS 1.05e-19 
C8386 VCC.n4468 VSS 3.5e-20 
C8387 VCC.n4469 VSS 3.5e-20 
C8388 VCC.n4470 VSS 8.42e-19 
C8389 VCC.n4471 VSS 2.18e-19 
C8390 VCC.n4472 VSS 1.4e-19 
C8391 VCC.n4473 VSS 4.32e-20 
C8392 VCC.n4474 VSS 7.82e-20 
C8393 VCC.n4475 VSS 5.76e-20 
C8394 VCC.n4476 VSS 2.68e-20 
C8395 VCC.n4477 VSS 4.32e-20 
C8396 VCC.n4478 VSS 3.91e-20 
C8397 VCC.n4479 VSS 3.7e-20 
C8398 VCC.n4480 VSS 3.7e-20 
C8399 VCC.n4481 VSS 5.76e-20 
C8400 VCC.n4482 VSS 4.73e-20 
C8401 VCC.n4483 VSS 3.5e-20 
C8402 VCC.t114 VSS 1.56e-19 
C8403 VCC.n4484 VSS 7.97e-19 
C8404 VCC.n4485 VSS 3.09e-20 
C8405 VCC.n4486 VSS 1.01e-19 
C8406 VCC.n4487 VSS 3.5e-20 
C8407 VCC.n4488 VSS 1.36e-19 
C8408 VCC.n4489 VSS 3.5e-20 
C8409 VCC.n4490 VSS 3.33e-19 
C8410 VCC.n4491 VSS 1.17e-19 
C8411 VCC.n4492 VSS 1.09e-19 
C8412 VCC.n4493 VSS 3.5e-20 
C8413 VCC.n4494 VSS 4.73e-20 
C8414 VCC.n4495 VSS 5.56e-20 
C8415 VCC.n4496 VSS 2.88e-20 
C8416 VCC.n4497 VSS 2.26e-20 
C8417 VCC.n4498 VSS 5.76e-20 
C8418 VCC.n4499 VSS 2.68e-20 
C8419 VCC.n4500 VSS 2.68e-20 
C8420 VCC.n4501 VSS 1.9e-19 
C8421 VCC.n4502 VSS 5.76e-20 
C8422 VCC.n4503 VSS 2.68e-20 
C8423 VCC.n4504 VSS 2.68e-20 
C8424 VCC.n4505 VSS 2.68e-20 
C8425 VCC.n4506 VSS 5.76e-20 
C8426 VCC.n4507 VSS 2.26e-20 
C8427 VCC.n4508 VSS 3.09e-20 
C8428 VCC.n4509 VSS 2.26e-20 
C8429 VCC.n4510 VSS 5.15e-20 
C8430 VCC.n4511 VSS 4.73e-20 
C8431 VCC.n4512 VSS 3.7e-20 
C8432 VCC.n4513 VSS 3.5e-20 
C8433 VCC.n4514 VSS 7.41e-20 
C8434 VCC.n4515 VSS 1.91e-19 
C8435 VCC.n4516 VSS 9.88e-20 
C8436 VCC.n4517 VSS 3e-20 
C8437 VCC.n4518 VSS 5.12e-19 
C8438 VCC.n4519 VSS 1.18e-19 
C8439 VCC.n4520 VSS 3.5e-20 
C8440 VCC.n4521 VSS 3.5e-20 
C8441 VCC.n4522 VSS 5.15e-20 
C8442 VCC.n4523 VSS 4.32e-20 
C8443 VCC.n4524 VSS 2.68e-20 
C8444 VCC.n4525 VSS 3.91e-20 
C8445 VCC.n4526 VSS 1.44e-20 
C8446 VCC.n4527 VSS 3.5e-20 
C8447 VCC.n4528 VSS 3e-20 
C8448 VCC.n4529 VSS 7.95e-19 
C8449 VCC.n4530 VSS 1.83e-19 
C8450 VCC.n4531 VSS 2.88e-20 
C8451 VCC.n4532 VSS 2.68e-20 
C8452 VCC.n4533 VSS 2.68e-20 
C8453 VCC.n4534 VSS 2.68e-20 
C8454 VCC.n4535 VSS 4.53e-20 
C8455 VCC.n4536 VSS 3.7e-20 
C8456 VCC.n4537 VSS 7.82e-20 
C8457 VCC.n4538 VSS 1.17e-19 
C8458 VCC.n4539 VSS 3.91e-20 
C8459 VCC.n4540 VSS 1.65e-20 
C8460 VCC.n4541 VSS 2.68e-20 
C8461 VCC.n4542 VSS 3.5e-20 
C8462 VCC.n4543 VSS 3e-20 
C8463 VCC.n4544 VSS 5.12e-19 
C8464 VCC.n4545 VSS 1.18e-19 
C8465 VCC.n4546 VSS 3.5e-20 
C8466 VCC.n4547 VSS 3.5e-20 
C8467 VCC.t160 VSS 1.55e-19 
C8468 VCC.n4548 VSS 7.57e-19 
C8469 VCC.n4549 VSS 4.73e-20 
C8470 VCC.n4550 VSS 1.54e-19 
C8471 VCC.n4551 VSS 2.88e-20 
C8472 VCC.n4552 VSS 2.88e-20 
C8473 VCC.n4553 VSS 3.5e-20 
C8474 VCC.n4554 VSS 5.76e-20 
C8475 VCC.n4555 VSS 9.88e-20 
C8476 VCC.n4556 VSS 1.3e-19 
C8477 VCC.n4557 VSS 3e-20 
C8478 VCC.t158 VSS 0.005f 
C8479 VCC.t163 VSS 0.00453f 
C8480 VCC.n4558 VSS 0.00229f 
C8481 VCC.n4559 VSS 1.91e-19 
C8482 VCC.n4560 VSS 3.5e-20 
C8483 VCC.n4561 VSS 3.14e-19 
C8484 VCC.n4562 VSS 3.5e-20 
C8485 VCC.n4563 VSS 2.47e-20 
C8486 VCC.n4564 VSS 5.76e-20 
C8487 VCC.n4565 VSS 2.47e-20 
C8488 VCC.n4566 VSS 8.23e-21 
C8489 VCC.n4567 VSS 2.88e-20 
C8490 VCC.n4568 VSS 5.76e-20 
C8491 VCC.n4569 VSS 2.47e-20 
C8492 VCC.n4570 VSS 2.88e-20 
C8493 VCC.n4571 VSS 2.47e-20 
C8494 VCC.n4572 VSS 5.15e-20 
C8495 VCC.n4573 VSS 4.73e-20 
C8496 VCC.n4574 VSS 3.7e-20 
C8497 VCC.n4575 VSS 3.5e-20 
C8498 VCC.n4576 VSS 7.41e-20 
C8499 VCC.t175 VSS 6.42e-19 
C8500 VCC.n4577 VSS 3e-20 
C8501 VCC.n4578 VSS 5.97e-20 
C8502 VCC.n4579 VSS 4.13e-19 
C8503 VCC.n4580 VSS 9.53e-20 
C8504 VCC.n4581 VSS 3.5e-20 
C8505 VCC.n4582 VSS 3.5e-20 
C8506 VCC.n4583 VSS 5.35e-20 
C8507 VCC.n4584 VSS 4.32e-20 
C8508 VCC.n4585 VSS 2.68e-20 
C8509 VCC.n4586 VSS 3.7e-20 
C8510 VCC.n4587 VSS 1.65e-20 
C8511 VCC.n4588 VSS 4.53e-20 
C8512 VCC.n4589 VSS 1.2e-19 
C8513 VCC.n4590 VSS 5.2e-19 
C8514 VCC.n4591 VSS 1.2e-19 
C8515 VCC.n4592 VSS 6.38e-20 
C8516 VCC.n4593 VSS 2.47e-20 
C8517 VCC.n4594 VSS 4.53e-20 
C8518 VCC.n4595 VSS 3.5e-20 
C8519 VCC.n4596 VSS 3.5e-20 
C8520 VCC.n4597 VSS 2.68e-20 
C8521 VCC.n4598 VSS 2.68e-20 
C8522 VCC.n4599 VSS 2.47e-20 
C8523 VCC.n4600 VSS 4.53e-20 
C8524 VCC.n4601 VSS 2.68e-20 
C8525 VCC.n4602 VSS 4.32e-20 
C8526 VCC.n4603 VSS 2.68e-20 
C8527 VCC.n4604 VSS 3.91e-20 
C8528 VCC.n4605 VSS 2.88e-20 
C8529 VCC.n4606 VSS 4.73e-20 
C8530 VCC.n4607 VSS 3.7e-20 
C8531 VCC.n4608 VSS 3.7e-20 
C8532 VCC.n4609 VSS 3.5e-20 
C8533 VCC.n4610 VSS 5.76e-20 
C8534 VCC.n4611 VSS 4.73e-20 
C8535 VCC.n4612 VSS 3.09e-20 
C8536 VCC.n4613 VSS 3.5e-20 
C8537 VCC.n4614 VSS 3.5e-20 
C8538 VCC.n4615 VSS 3.5e-20 
C8539 VCC.n4616 VSS 1.18e-19 
C8540 VCC.n4617 VSS 3e-20 
C8541 VCC.n4618 VSS 1.15e-19 
C8542 VCC.n4619 VSS 9.88e-20 
C8543 VCC.n4620 VSS 5.76e-20 
C8544 VCC.n4621 VSS 3.5e-20 
C8545 VCC.n4622 VSS 3.09e-20 
C8546 VCC.n4623 VSS 3.09e-20 
C8547 VCC.n4624 VSS 2.26e-20 
C8548 VCC.n4625 VSS 5.76e-20 
C8549 VCC.n4626 VSS 2.68e-20 
C8550 VCC.n4627 VSS 2.68e-20 
C8551 VCC.n4628 VSS 0.00185f 
C8552 VCC.n4629 VSS 2.72e-19 
C8553 VCC.n4630 VSS 2.26e-20 
C8554 VCC.n4631 VSS 1.87e-19 
C8555 VCC.n4632 VSS 3.5e-20 
C8556 VCC.n4633 VSS 2.68e-20 
C8557 VCC.n4634 VSS 5.97e-20 
C8558 VCC.n4635 VSS 4.73e-20 
C8559 VCC.n4636 VSS 4.73e-20 
C8560 VCC.n4637 VSS 5.15e-20 
C8561 VCC.n4638 VSS 7.41e-20 
C8562 VCC.n4639 VSS 3.7e-20 
C8563 VCC.n4640 VSS 2.26e-20 
C8564 VCC.n4641 VSS 6.38e-20 
C8565 VCC.n4642 VSS 4.73e-20 
C8566 VCC.n4643 VSS 3.29e-20 
C8567 VCC.n4644 VSS 3.5e-20 
C8568 VCC.n4645 VSS 3e-20 
C8569 VCC.t58 VSS 0.005f 
C8570 VCC.t258 VSS 0.00453f 
C8571 VCC.n4646 VSS 0.00228f 
C8572 VCC.n4647 VSS 1.3e-19 
C8573 VCC.t56 VSS 4.05e-19 
C8574 VCC.n4648 VSS 4.05e-19 
C8575 VCC.n4649 VSS 1.15e-19 
C8576 VCC.n4650 VSS 3.36e-19 
C8577 VCC.n4651 VSS 6.17e-21 
C8578 VCC.n4652 VSS 3.12e-19 
C8579 VCC.n4653 VSS 1.65e-20 
C8580 VCC.n4654 VSS 1.54e-19 
C8581 VCC.n4655 VSS 1.54e-19 
C8582 VCC.n4656 VSS 1.65e-20 
C8583 VCC.n4657 VSS 1.03e-20 
C8584 VCC.n4658 VSS 3.5e-20 
C8585 VCC.n4659 VSS 2.26e-20 
C8586 VCC.n4660 VSS 4.73e-20 
C8587 VCC.n4661 VSS 3.5e-20 
C8588 VCC.n4662 VSS 3e-20 
C8589 VCC.n4663 VSS 1.3e-19 
C8590 VCC.n4664 VSS 5.12e-19 
C8591 VCC.n4665 VSS 1.3e-19 
C8592 VCC.n4666 VSS 4.13e-19 
C8593 VCC.n4667 VSS 9.53e-20 
C8594 VCC.n4668 VSS 5.76e-20 
C8595 VCC.n4669 VSS 7.41e-20 
C8596 VCC.n4670 VSS 5.56e-20 
C8597 VCC.t57 VSS 1.55e-19 
C8598 VCC.n4671 VSS 3.91e-20 
C8599 VCC.n4672 VSS 3.91e-20 
C8600 VCC.n4673 VSS 1.85e-20 
C8601 VCC.n4674 VSS 7.55e-19 
C8602 VCC.n4675 VSS 4.94e-20 
C8603 VCC.n4676 VSS 5.15e-20 
C8604 VCC.n4677 VSS 7.2e-20 
C8605 VCC.n4678 VSS 1.38e-19 
C8606 VCC.n4679 VSS 1.17e-19 
C8607 VCC.n4680 VSS 4.32e-20 
C8608 VCC.n4681 VSS 2.88e-20 
C8609 VCC.n4682 VSS 2.68e-20 
C8610 VCC.n4683 VSS 3.5e-20 
C8611 VCC.n4684 VSS 3.5e-20 
C8612 VCC.n4685 VSS 2.88e-20 
C8613 VCC.n4686 VSS 2.68e-20 
C8614 VCC.n4687 VSS 2.68e-20 
C8615 VCC.n4688 VSS 2.68e-20 
C8616 VCC.n4689 VSS 4.12e-20 
C8617 VCC.n4690 VSS 4.12e-20 
C8618 VCC.n4691 VSS 3.91e-20 
C8619 VCC.n4692 VSS 4.53e-20 
C8620 VCC.n4693 VSS 4.53e-20 
C8621 VCC.n4694 VSS 1.05e-19 
C8622 VCC.n4695 VSS 1.05e-19 
C8623 VCC.n4696 VSS 4.32e-20 
C8624 VCC.n4697 VSS 3.7e-20 
C8625 VCC.n4698 VSS 2.68e-20 
C8626 VCC.n4699 VSS 2.68e-20 
C8627 VCC.n4700 VSS 6.79e-20 
C8628 VCC.n4701 VSS 9.26e-20 
C8629 VCC.n4702 VSS 1.83e-19 
C8630 VCC.n4703 VSS 7.95e-19 
C8631 VCC.n4704 VSS 5.2e-19 
C8632 VCC.n4705 VSS 1.3e-19 
C8633 VCC.n4706 VSS 3e-20 
C8634 VCC.n4707 VSS 3.5e-20 
C8635 VCC.n4708 VSS 5.97e-20 
C8636 VCC.n4709 VSS 7.41e-20 
C8637 VCC.n4710 VSS 5.15e-20 
C8638 VCC.n4711 VSS 5.15e-20 
C8639 VCC.n4712 VSS 3.09e-20 
C8640 VCC.n4713 VSS 3.09e-20 
C8641 VCC.n4714 VSS 3.7e-20 
C8642 VCC.n4715 VSS 2.68e-20 
C8643 VCC.n4716 VSS 3.91e-20 
C8644 VCC.n4717 VSS 1.17e-19 
C8645 VCC.n4718 VSS 1.38e-19 
C8646 VCC.n4719 VSS 7e-20 
C8647 VCC.n4720 VSS 4.73e-20 
C8648 VCC.n4721 VSS 3.5e-20 
C8649 VCC.n4722 VSS 3.5e-20 
C8650 VCC.n4723 VSS 3.5e-20 
C8651 VCC.n4724 VSS 4.53e-20 
C8652 VCC.n4725 VSS 1.18e-19 
C8653 VCC.n4726 VSS 5.12e-19 
C8654 VCC.n4727 VSS 1.3e-19 
C8655 VCC.n4728 VSS 1.61e-19 
C8656 VCC.n4729 VSS 9.9e-20 
C8657 VCC.n4730 VSS 0.00243f 
C8658 VCC.n4731 VSS 2.26e-20 
C8659 VCC.n4732 VSS 4.13e-19 
C8660 VCC.n4733 VSS 3.5e-20 
C8661 VCC.n4734 VSS 3.5e-20 
C8662 VCC.n4735 VSS 2.47e-20 
C8663 VCC.n4736 VSS 2.06e-20 
C8664 VCC.n4737 VSS 6.17e-20 
C8665 VCC.n4738 VSS 6.17e-20 
C8666 VCC.n4739 VSS 4.73e-20 
C8667 VCC.n4740 VSS 4.73e-20 
C8668 VCC.n4741 VSS 2.88e-20 
C8669 VCC.n4742 VSS 1.44e-20 
C8670 VCC.n4743 VSS 1.65e-20 
C8671 VCC.n4744 VSS 1.54e-19 
C8672 VCC.n4745 VSS 1.54e-19 
C8673 VCC.n4746 VSS 1.65e-20 
C8674 VCC.n4747 VSS 3.09e-20 
C8675 VCC.t176 VSS 1.55e-19 
C8676 VCC.n4748 VSS 0.00102f 
C8677 VCC.n4749 VSS 2.73e-19 
C8678 VCC.n4750 VSS 0.00136f 
C8679 VCC.n4751 VSS 2.73e-19 
C8680 VCC.n4752 VSS 0.00181f 
C8681 VCC.n4753 VSS 5.76e-20 
C8682 VCC.n4754 VSS 1.54e-19 
C8683 VCC.n4755 VSS 1.65e-20 
C8684 VCC.n4756 VSS 6.17e-20 
C8685 VCC.n4757 VSS 2.47e-20 
C8686 VCC.n4758 VSS 4.73e-20 
C8687 VCC.n4759 VSS 4.73e-20 
C8688 VCC.n4760 VSS 5.15e-20 
C8689 VCC.n4761 VSS 3.5e-20 
C8690 VCC.n4762 VSS 7.41e-20 
C8691 VCC.n4763 VSS 3.7e-20 
C8692 VCC.n4764 VSS 2.26e-20 
C8693 VCC.n4765 VSS 6.17e-20 
C8694 VCC.n4766 VSS 4.73e-20 
C8695 VCC.n4767 VSS 2.88e-20 
C8696 VCC.n4768 VSS 2.88e-20 
C8697 VCC.n4769 VSS 3.4e-19 
C8698 VCC.n4770 VSS 1.15e-19 
C8699 VCC.n4771 VSS 3.98e-19 
C8700 VCC.t159 VSS 4.05e-19 
C8701 VCC.n4772 VSS 1.22e-19 
C8702 VCC.n4773 VSS 1.3e-19 
C8703 VCC.n4774 VSS 3e-20 
C8704 VCC.n4775 VSS 3.5e-20 
C8705 VCC.n4776 VSS 3.5e-20 
C8706 VCC.n4777 VSS 4.73e-20 
C8707 VCC.n4778 VSS 2.47e-20 
C8708 VCC.n4779 VSS 1.23e-20 
C8709 VCC.n4780 VSS 1.65e-20 
C8710 VCC.n4781 VSS 2.47e-20 
C8711 VCC.n4782 VSS 5.76e-20 
C8712 VCC.n4783 VSS 1.38e-19 
C8713 VCC.n4784 VSS 7e-20 
C8714 VCC.n4785 VSS 3.7e-20 
C8715 VCC.n4786 VSS 2.47e-20 
C8716 VCC.n4787 VSS 3.7e-20 
C8717 VCC.n4788 VSS 1.85e-20 
C8718 VCC.n4789 VSS 3.09e-20 
C8719 VCC.n4790 VSS 5.35e-20 
C8720 VCC.n4791 VSS 4.73e-20 
C8721 VCC.n4792 VSS 5.35e-20 
C8722 VCC.n4793 VSS 7.41e-20 
C8723 VCC.n4794 VSS 5.76e-20 
C8724 VCC.n4795 VSS 9.53e-20 
C8725 VCC.n4796 VSS 4.13e-19 
C8726 VCC.n4797 VSS 1.3e-19 
C8727 VCC.n4798 VSS 5.2e-19 
C8728 VCC.n4799 VSS 1.2e-19 
C8729 VCC.n4800 VSS 4.73e-20 
C8730 VCC.n4801 VSS 2.68e-20 
C8731 VCC.n4802 VSS 3.5e-20 
C8732 VCC.n4803 VSS 3.5e-20 
C8733 VCC.n4804 VSS 2.68e-20 
C8734 VCC.n4805 VSS 2.68e-20 
C8735 VCC.n4806 VSS 4.32e-20 
C8736 VCC.n4807 VSS 4.32e-20 
C8737 VCC.n4808 VSS 4.32e-20 
C8738 VCC.n4809 VSS 2.88e-20 
C8739 VCC.n4810 VSS 3.5e-20 
C8740 VCC.n4811 VSS 2.68e-20 
C8741 VCC.n4812 VSS 7.82e-20 
C8742 VCC.n4813 VSS 4.73e-20 
C8743 VCC.n4814 VSS 4.73e-20 
C8744 VCC.n4815 VSS 1.05e-19 
C8745 VCC.n4816 VSS 1.05e-19 
C8746 VCC.n4817 VSS 4.53e-20 
C8747 VCC.n4818 VSS 2.68e-20 
C8748 VCC.n4819 VSS 2.68e-20 
C8749 VCC.n4820 VSS 6.59e-20 
C8750 VCC.n4821 VSS 9.26e-20 
C8751 VCC.n4822 VSS 6.59e-20 
C8752 VCC.n4823 VSS 2.47e-20 
C8753 VCC.n4824 VSS 2.47e-20 
C8754 VCC.n4825 VSS 2.88e-20 
C8755 VCC.n4826 VSS 3.5e-20 
C8756 VCC.n4827 VSS 3.5e-20 
C8757 VCC.n4828 VSS 4.53e-20 
C8758 VCC.n4829 VSS 1.2e-19 
C8759 VCC.n4830 VSS 5.2e-19 
C8760 VCC.n4831 VSS 1.3e-19 
C8761 VCC.n4832 VSS 4.13e-19 
C8762 VCC.n4833 VSS 9.53e-20 
C8763 VCC.n4834 VSS 5.97e-20 
C8764 VCC.n4835 VSS 7.41e-20 
C8765 VCC.n4836 VSS 5.35e-20 
C8766 VCC.n4837 VSS 5.15e-20 
C8767 VCC.n4838 VSS 3.09e-20 
C8768 VCC.n4839 VSS 3.09e-20 
C8769 VCC.n4840 VSS 3.91e-20 
C8770 VCC.n4841 VSS 2.47e-20 
C8771 VCC.n4842 VSS 3.7e-20 
C8772 VCC.n4843 VSS 1.17e-19 
C8773 VCC.n4844 VSS 1.38e-19 
C8774 VCC.n4845 VSS 7.2e-20 
C8775 VCC.n4846 VSS 4.73e-20 
C8776 VCC.n4847 VSS 3.5e-20 
C8777 VCC.n4848 VSS 3.5e-20 
C8778 VCC.n4849 VSS 4.53e-20 
C8779 VCC.n4850 VSS 5.97e-20 
C8780 VCC.n4851 VSS 3.5e-20 
C8781 VCC.n4852 VSS 3e-20 
C8782 VCC.n4853 VSS 1.3e-19 
C8783 VCC.n4854 VSS 1.53e-19 
C8784 VCC.t123 VSS 4.05e-19 
C8785 VCC.n4855 VSS 1.35e-19 
C8786 VCC.t113 VSS 4.21e-19 
C8787 VCC.n4856 VSS 2.06e-19 
C8788 VCC.n4857 VSS 1.32e-19 
C8789 VCC.n4858 VSS 9.67e-20 
C8790 VCC.n4859 VSS 3.35e-20 
C8791 VCC.n4860 VSS 3.5e-20 
C8792 VCC.n4861 VSS 2.36e-19 
C8793 VCC.n4862 VSS 0.0023f 
C8794 VCC.t112 VSS 0.0031f 
C8795 VCC.t115 VSS 0.00366f 
C8796 VCC.t111 VSS 0.00365f 
C8797 VCC.t118 VSS 0.00386f 
C8798 VCC.n4863 VSS 0.00569f 
C8799 VCC.n4864 VSS 1.3e-19 
C8800 VCC.n4865 VSS 3.67e-19 
C8801 VCC.n4866 VSS 1.15e-19 
C8802 VCC.n4867 VSS 3.38e-19 
C8803 VCC.n4868 VSS 3.5e-20 
C8804 VCC.n4869 VSS 3.5e-20 
C8805 VCC.n4870 VSS 2.68e-20 
C8806 VCC.n4871 VSS 2.06e-20 
C8807 VCC.n4872 VSS 6.38e-20 
C8808 VCC.n4873 VSS 5.97e-20 
C8809 VCC.n4874 VSS 4.73e-20 
C8810 VCC.n4875 VSS 4.73e-20 
C8811 VCC.n4876 VSS 3.09e-20 
C8812 VCC.n4877 VSS 1.23e-20 
C8813 VCC.n4878 VSS 1.65e-20 
C8814 VCC.n4879 VSS 1.54e-19 
C8815 VCC.n4880 VSS 1.54e-19 
C8816 VCC.n4881 VSS 1.65e-20 
C8817 VCC.n4882 VSS 3.29e-20 
C8818 VCC.t124 VSS 1.67e-19 
C8819 VCC.n4883 VSS 0.00101f 
C8820 VCC.n4884 VSS 2.71e-19 
C8821 VCC.n4885 VSS 7.46e-19 
C8822 VCC.n4886 VSS 0.00333f 
C8823 VCC.n4887 VSS 2.46e-19 
C8824 VCC.n4888 VSS 3.02e-19 
C8825 VCC.n4889 VSS 3.7e-20 
C8826 VCC.n4890 VSS 5.15e-20 
C8827 VCC.n4891 VSS 5.97e-20 
C8828 VCC.n4892 VSS 6.38e-20 
C8829 VCC.n4893 VSS 4.73e-20 
C8830 VCC.n4894 VSS 4.73e-20 
C8831 VCC.n4895 VSS 2.68e-20 
C8832 VCC.n4896 VSS 3.29e-20 
C8833 VCC.n4897 VSS 1.65e-20 
C8834 VCC.n4898 VSS 1.54e-19 
C8835 VCC.n4899 VSS 1.54e-19 
C8836 VCC.n4900 VSS 1.65e-20 
C8837 VCC.n4901 VSS 3.09e-20 
C8838 VCC.n4902 VSS 3.09e-20 
C8839 VCC.n4903 VSS 4.73e-20 
C8840 VCC.n4904 VSS 4.32e-20 
C8841 VCC.n4905 VSS 3.5e-20 
C8842 VCC.n4906 VSS 3.5e-20 
C8843 VCC.n4907 VSS 1.35e-19 
C8844 VCC.n4908 VSS 5.24e-19 
C8845 VCC.n4909 VSS 1.4e-19 
C8846 VCC.n4910 VSS 5.4e-19 
C8847 VCC.n4911 VSS 1.35e-19 
C8848 VCC.n4912 VSS 4.37e-19 
C8849 VCC.n4913 VSS 1.13e-19 
C8850 VCC.n4914 VSS 8.23e-21 
C8851 VCC.n4915 VSS 1.65e-20 
C8852 VCC.n4916 VSS 3.5e-20 
C8853 VCC.n4917 VSS 3.91e-20 
C8854 VCC.n4918 VSS 3.09e-20 
C8855 VCC.n4919 VSS 1.85e-20 
C8856 VCC.n4920 VSS 3.5e-20 
C8857 VCC.n4921 VSS 1.05e-19 
C8858 VCC.n4922 VSS 2.06e-20 
C8859 VCC.n4923 VSS 2.26e-20 
C8860 VCC.n4924 VSS 3.7e-20 
C8861 VCC.n4925 VSS 5.15e-20 
C8862 VCC.n4926 VSS 1.38e-19 
C8863 VCC.n4927 VSS 1.17e-19 
C8864 VCC.n4928 VSS 4.32e-20 
C8865 VCC.n4929 VSS 2.88e-20 
C8866 VCC.n4930 VSS 2.68e-20 
C8867 VCC.n4931 VSS 6.59e-20 
C8868 VCC.n4932 VSS 5.56e-20 
C8869 VCC.n4933 VSS 2.68e-20 
C8870 VCC.n4934 VSS 4.32e-20 
C8871 VCC.n4935 VSS 1.05e-19 
C8872 VCC.n4936 VSS 3.09e-20 
C8873 VCC.n4937 VSS 3.7e-20 
C8874 VCC.n4938 VSS 4.32e-20 
C8875 VCC.n4939 VSS 1.05e-19 
C8876 VCC.n4940 VSS 4.53e-20 
C8877 VCC.n4941 VSS 4.53e-20 
C8878 VCC.n4942 VSS 7.82e-20 
C8879 VCC.n4943 VSS 2.18e-19 
C8880 VCC.n4944 VSS 1.4e-19 
C8881 VCC.n4945 VSS 1.4e-19 
C8882 VCC.n4946 VSS 5.4e-19 
C8883 VCC.n4947 VSS 1.35e-19 
C8884 VCC.t264 VSS 4.21e-19 
C8885 VCC.n4948 VSS 3.33e-19 
C8886 VCC.n4949 VSS 1.13e-19 
C8887 VCC.n4950 VSS 8.23e-21 
C8888 VCC.n4951 VSS 1.65e-20 
C8889 VCC.n4952 VSS 3.5e-20 
C8890 VCC.n4953 VSS 3.5e-20 
C8891 VCC.n4954 VSS 3.5e-20 
C8892 VCC.n4955 VSS 1.17e-19 
C8893 VCC.n4956 VSS 1.38e-19 
C8894 VCC.n4957 VSS 5.15e-20 
C8895 VCC.n4958 VSS 4.73e-20 
C8896 VCC.n4959 VSS 7.2e-20 
C8897 VCC.n4960 VSS 2.68e-20 
C8898 VCC.n4961 VSS 1.65e-20 
C8899 VCC.n4962 VSS 1.54e-19 
C8900 VCC.n4963 VSS 1.54e-19 
C8901 VCC.n4964 VSS 1.65e-20 
C8902 VCC.n4965 VSS 2.47e-20 
C8903 VCC.n4966 VSS 1.23e-20 
C8904 VCC.n4967 VSS 7.62e-19 
C8905 VCC.n4968 VSS 4.12e-20 
C8906 VCC.n4969 VSS 5.15e-20 
C8907 VCC.n4970 VSS 6.59e-20 
C8908 VCC.n4971 VSS 5.76e-20 
C8909 VCC.n4972 VSS 4.73e-20 
C8910 VCC.n4973 VSS 2.26e-20 
C8911 VCC.n4974 VSS 2.68e-20 
C8912 VCC.n4975 VSS 1.03e-20 
C8913 VCC.n4976 VSS 3.5e-20 
C8914 VCC.n4977 VSS 3.5e-20 
C8915 VCC.n4978 VSS 1.35e-19 
C8916 VCC.n4979 VSS 4.53e-19 
C8917 VCC.n4980 VSS 7.71e-19 
C8918 VCC.n4981 VSS 1.32e-19 
C8919 VCC.n4982 VSS 3.5e-20 
C8920 VCC.n4983 VSS 3.42e-20 
C8921 VCC.n4984 VSS 2.36e-19 
C8922 VCC.n4985 VSS 3.21e-19 
C8923 VCC.n4986 VSS 2.61e-19 
C8924 VCC.n4987 VSS 0.00189f 
C8925 VCC.n4988 VSS 2.68e-19 
C8926 VCC.n4989 VSS 5.22e-19 
C8927 VCC.n4990 VSS 5.76e-20 
C8928 VCC.n4991 VSS 2.88e-20 
C8929 VCC.n4992 VSS 3.5e-20 
C8930 VCC.n4993 VSS 3.42e-20 
C8931 VCC.n4994 VSS 3.5e-20 
C8932 VCC.n4995 VSS 4.53e-19 
C8933 VCC.n4996 VSS 1.17e-19 
C8934 VCC.n4997 VSS 3.5e-20 
C8935 VCC.n4998 VSS 1.44e-20 
C8936 VCC.n4999 VSS 4.12e-20 
C8937 VCC.n5000 VSS 5.76e-20 
C8938 VCC.n5001 VSS 5.76e-20 
C8939 VCC.n5002 VSS 2.06e-20 
C8940 VCC.n5003 VSS 3.29e-20 
C8941 VCC.n5004 VSS 7.2e-20 
C8942 VCC.n5005 VSS 3.29e-20 
C8943 VCC.n5006 VSS 4.73e-20 
C8944 VCC.n5007 VSS 2.26e-20 
C8945 VCC.n5008 VSS 1.01e-19 
C8946 VCC.n5009 VSS 1.36e-19 
C8947 VCC.n5010 VSS 1.35e-19 
C8948 VCC.n5011 VSS 3.5e-20 
C8949 VCC.n5012 VSS 3.5e-20 
C8950 VCC.n5013 VSS 3.5e-20 
C8951 VCC.n5014 VSS 3.5e-20 
C8952 VCC.n5015 VSS 3.09e-20 
C8953 VCC.n5016 VSS 3.91e-20 
C8954 VCC.n5017 VSS 4.73e-20 
C8955 VCC.n5018 VSS 4.32e-20 
C8956 VCC.n5019 VSS 2.68e-20 
C8957 VCC.n5020 VSS 4.53e-20 
C8958 VCC.n5021 VSS 4.53e-20 
C8959 VCC.n5022 VSS 3.09e-20 
C8960 VCC.n5023 VSS 4.32e-20 
C8961 VCC.n5024 VSS 2.68e-20 
C8962 VCC.n5025 VSS 7.82e-20 
C8963 VCC.n5026 VSS 5.56e-20 
C8964 VCC.n5027 VSS 1.4e-19 
C8965 VCC.n5028 VSS 2.18e-19 
C8966 VCC.n5029 VSS 1.35e-19 
C8967 VCC.n5030 VSS 1.13e-19 
C8968 VCC.n5031 VSS 3.5e-20 
C8969 VCC.n5032 VSS 1.85e-20 
C8970 VCC.n5033 VSS 3.7e-20 
C8971 VCC.n5034 VSS 3.09e-20 
C8972 VCC.n5035 VSS 6.59e-20 
C8973 VCC.n5036 VSS 2.68e-20 
C8974 VCC.n5037 VSS 5.76e-20 
C8975 VCC.n5038 VSS 4.73e-20 
C8976 VCC.n5039 VSS 3.5e-20 
C8977 VCC.t224 VSS 1.56e-19 
C8978 VCC.n5040 VSS 7.97e-19 
C8979 VCC.n5041 VSS 3.09e-20 
C8980 VCC.n5042 VSS 3.5e-20 
C8981 VCC.n5043 VSS 3.5e-20 
C8982 VCC.t223 VSS 4.21e-19 
C8983 VCC.n5044 VSS 1.32e-19 
C8984 VCC.n5045 VSS 1.09e-19 
C8985 VCC.n5046 VSS 3.5e-20 
C8986 VCC.n5047 VSS 3.09e-20 
C8987 VCC.n5048 VSS 5.97e-20 
C8988 VCC.n5049 VSS 2.26e-20 
C8989 VCC.n5050 VSS 5.76e-20 
C8990 VCC.n5051 VSS 2.68e-20 
C8991 VCC.n5052 VSS 2.68e-20 
C8992 VCC.n5053 VSS 1.9e-19 
C8993 VCC.n5054 VSS 5.76e-20 
C8994 VCC.n5055 VSS 2.68e-20 
C8995 VCC.n5056 VSS 2.68e-20 
C8996 VCC.n5057 VSS 2.68e-20 
C8997 VCC.n5058 VSS 5.76e-20 
C8998 VCC.n5059 VSS 2.26e-20 
C8999 VCC.n5060 VSS 3.09e-20 
C9000 VCC.n5061 VSS 2.26e-20 
C9001 VCC.n5062 VSS 5.15e-20 
C9002 VCC.n5063 VSS 4.73e-20 
C9003 VCC.n5064 VSS 3.7e-20 
C9004 VCC.n5065 VSS 3.5e-20 
C9005 VCC.n5066 VSS 7.41e-20 
C9006 VCC.n5067 VSS 1.91e-19 
C9007 VCC.n5068 VSS 9.88e-20 
C9008 VCC.n5069 VSS 3e-20 
C9009 VCC.n5070 VSS 5.12e-19 
C9010 VCC.n5071 VSS 1.18e-19 
C9011 VCC.n5072 VSS 3.5e-20 
C9012 VCC.n5073 VSS 3.5e-20 
C9013 VCC.n5074 VSS 5.15e-20 
C9014 VCC.n5075 VSS 4.32e-20 
C9015 VCC.n5076 VSS 2.68e-20 
C9016 VCC.n5077 VSS 3.91e-20 
C9017 VCC.n5078 VSS 1.44e-20 
C9018 VCC.n5079 VSS 3.5e-20 
C9019 VCC.n5080 VSS 3e-20 
C9020 VCC.n5081 VSS 7.95e-19 
C9021 VCC.n5082 VSS 1.83e-19 
C9022 VCC.n5083 VSS 2.88e-20 
C9023 VCC.n5084 VSS 2.68e-20 
C9024 VCC.n5085 VSS 2.68e-20 
C9025 VCC.n5086 VSS 2.68e-20 
C9026 VCC.n5087 VSS 4.53e-20 
C9027 VCC.n5088 VSS 3.7e-20 
C9028 VCC.n5089 VSS 7.82e-20 
C9029 VCC.n5090 VSS 1.17e-19 
C9030 VCC.n5091 VSS 3.91e-20 
C9031 VCC.n5092 VSS 1.65e-20 
C9032 VCC.n5093 VSS 2.68e-20 
C9033 VCC.n5094 VSS 3.5e-20 
C9034 VCC.n5095 VSS 3e-20 
C9035 VCC.n5096 VSS 5.12e-19 
C9036 VCC.n5097 VSS 1.18e-19 
C9037 VCC.n5098 VSS 3.5e-20 
C9038 VCC.n5099 VSS 3.5e-20 
C9039 VCC.t234 VSS 1.55e-19 
C9040 VCC.n5100 VSS 7.57e-19 
C9041 VCC.n5101 VSS 4.73e-20 
C9042 VCC.n5102 VSS 1.54e-19 
C9043 VCC.n5103 VSS 2.88e-20 
C9044 VCC.n5104 VSS 2.88e-20 
C9045 VCC.n5105 VSS 3.5e-20 
C9046 VCC.n5106 VSS 5.76e-20 
C9047 VCC.n5107 VSS 9.88e-20 
C9048 VCC.n5108 VSS 1.3e-19 
C9049 VCC.n5109 VSS 3e-20 
C9050 VCC.t232 VSS 0.005f 
C9051 VCC.t241 VSS 0.00453f 
C9052 VCC.n5110 VSS 0.00229f 
C9053 VCC.n5111 VSS 1.91e-19 
C9054 VCC.n5112 VSS 3.5e-20 
C9055 VCC.n5113 VSS 3.14e-19 
C9056 VCC.n5114 VSS 2.47e-20 
C9057 VCC.n5115 VSS 5.76e-20 
C9058 VCC.n5116 VSS 2.47e-20 
C9059 VCC.n5117 VSS 8.23e-21 
C9060 VCC.n5118 VSS 2.88e-20 
C9061 VCC.n5119 VSS 5.76e-20 
C9062 VCC.n5120 VSS 2.47e-20 
C9063 VCC.n5121 VSS 2.88e-20 
C9064 VCC.n5122 VSS 2.47e-20 
C9065 VCC.n5123 VSS 5.15e-20 
C9066 VCC.n5124 VSS 4.73e-20 
C9067 VCC.n5125 VSS 3.7e-20 
C9068 VCC.n5126 VSS 3.5e-20 
C9069 VCC.n5127 VSS 7.41e-20 
C9070 VCC.t125 VSS 6.42e-19 
C9071 VCC.n5128 VSS 3e-20 
C9072 VCC.n5129 VSS 5.97e-20 
C9073 VCC.n5130 VSS 4.13e-19 
C9074 VCC.n5131 VSS 9.53e-20 
C9075 VCC.n5132 VSS 3.5e-20 
C9076 VCC.n5133 VSS 3.5e-20 
C9077 VCC.n5134 VSS 5.35e-20 
C9078 VCC.n5135 VSS 4.32e-20 
C9079 VCC.n5136 VSS 2.68e-20 
C9080 VCC.n5137 VSS 3.7e-20 
C9081 VCC.n5138 VSS 1.65e-20 
C9082 VCC.n5139 VSS 4.53e-20 
C9083 VCC.n5140 VSS 1.2e-19 
C9084 VCC.n5141 VSS 5.2e-19 
C9085 VCC.n5142 VSS 1.2e-19 
C9086 VCC.n5143 VSS 6.38e-20 
C9087 VCC.n5144 VSS 2.47e-20 
C9088 VCC.n5145 VSS 4.53e-20 
C9089 VCC.n5146 VSS 3.5e-20 
C9090 VCC.n5147 VSS 3.5e-20 
C9091 VCC.n5148 VSS 2.68e-20 
C9092 VCC.n5149 VSS 2.68e-20 
C9093 VCC.n5150 VSS 2.47e-20 
C9094 VCC.n5151 VSS 4.53e-20 
C9095 VCC.n5152 VSS 2.68e-20 
C9096 VCC.n5153 VSS 4.32e-20 
C9097 VCC.n5154 VSS 2.68e-20 
C9098 VCC.n5155 VSS 3.91e-20 
C9099 VCC.n5156 VSS 2.88e-20 
C9100 VCC.n5157 VSS 4.73e-20 
C9101 VCC.n5158 VSS 3.7e-20 
C9102 VCC.n5159 VSS 3.7e-20 
C9103 VCC.n5160 VSS 3.5e-20 
C9104 VCC.n5161 VSS 5.76e-20 
C9105 VCC.n5162 VSS 4.73e-20 
C9106 VCC.n5163 VSS 3.09e-20 
C9107 VCC.n5164 VSS 3.5e-20 
C9108 VCC.n5165 VSS 3.5e-20 
C9109 VCC.n5166 VSS 3.5e-20 
C9110 VCC.n5167 VSS 1.18e-19 
C9111 VCC.n5168 VSS 3e-20 
C9112 VCC.n5169 VSS 1.15e-19 
C9113 VCC.n5170 VSS 9.88e-20 
C9114 VCC.n5171 VSS 5.76e-20 
C9115 VCC.n5172 VSS 3.5e-20 
C9116 VCC.n5173 VSS 3.09e-20 
C9117 VCC.n5174 VSS 3.09e-20 
C9118 VCC.n5175 VSS 2.26e-20 
C9119 VCC.n5176 VSS 5.76e-20 
C9120 VCC.n5177 VSS 2.68e-20 
C9121 VCC.n5178 VSS 2.68e-20 
C9122 VCC.n5179 VSS 0.00185f 
C9123 VCC.n5180 VSS 2.72e-19 
C9124 VCC.n5181 VSS 2.26e-20 
C9125 VCC.n5182 VSS 1.87e-19 
C9126 VCC.n5183 VSS 3.5e-20 
C9127 VCC.n5184 VSS 2.68e-20 
C9128 VCC.n5185 VSS 5.97e-20 
C9129 VCC.n5186 VSS 4.73e-20 
C9130 VCC.n5187 VSS 4.73e-20 
C9131 VCC.n5188 VSS 5.15e-20 
C9132 VCC.n5189 VSS 7.41e-20 
C9133 VCC.n5190 VSS 3.7e-20 
C9134 VCC.n5191 VSS 2.26e-20 
C9135 VCC.n5192 VSS 6.38e-20 
C9136 VCC.n5193 VSS 4.73e-20 
C9137 VCC.n5194 VSS 3.29e-20 
C9138 VCC.n5195 VSS 3.5e-20 
C9139 VCC.n5196 VSS 3e-20 
C9140 VCC.t142 VSS 0.005f 
C9141 VCC.t171 VSS 0.00453f 
C9142 VCC.n5197 VSS 0.00228f 
C9143 VCC.n5198 VSS 1.3e-19 
C9144 VCC.t140 VSS 4.05e-19 
C9145 VCC.n5199 VSS 4.05e-19 
C9146 VCC.n5200 VSS 1.15e-19 
C9147 VCC.n5201 VSS 3.36e-19 
C9148 VCC.n5202 VSS 6.17e-21 
C9149 VCC.n5203 VSS 3.12e-19 
C9150 VCC.n5204 VSS 1.65e-20 
C9151 VCC.n5205 VSS 1.54e-19 
C9152 VCC.n5206 VSS 1.54e-19 
C9153 VCC.n5207 VSS 1.65e-20 
C9154 VCC.n5208 VSS 1.03e-20 
C9155 VCC.n5209 VSS 3.5e-20 
C9156 VCC.n5210 VSS 2.26e-20 
C9157 VCC.n5211 VSS 4.73e-20 
C9158 VCC.n5212 VSS 3.5e-20 
C9159 VCC.n5213 VSS 3e-20 
C9160 VCC.n5214 VSS 1.3e-19 
C9161 VCC.n5215 VSS 5.12e-19 
C9162 VCC.n5216 VSS 1.3e-19 
C9163 VCC.n5217 VSS 4.13e-19 
C9164 VCC.n5218 VSS 9.53e-20 
C9165 VCC.n5219 VSS 5.76e-20 
C9166 VCC.n5220 VSS 7.41e-20 
C9167 VCC.n5221 VSS 5.56e-20 
C9168 VCC.t141 VSS 1.55e-19 
C9169 VCC.n5222 VSS 3.91e-20 
C9170 VCC.n5223 VSS 3.91e-20 
C9171 VCC.n5224 VSS 1.85e-20 
C9172 VCC.n5225 VSS 7.55e-19 
C9173 VCC.n5226 VSS 4.94e-20 
C9174 VCC.n5227 VSS 5.15e-20 
C9175 VCC.n5228 VSS 7.2e-20 
C9176 VCC.n5229 VSS 1.38e-19 
C9177 VCC.n5230 VSS 1.17e-19 
C9178 VCC.n5231 VSS 4.32e-20 
C9179 VCC.n5232 VSS 2.88e-20 
C9180 VCC.n5233 VSS 2.68e-20 
C9181 VCC.n5234 VSS 3.5e-20 
C9182 VCC.n5235 VSS 3.5e-20 
C9183 VCC.n5236 VSS 2.88e-20 
C9184 VCC.n5237 VSS 2.68e-20 
C9185 VCC.n5238 VSS 2.68e-20 
C9186 VCC.n5239 VSS 2.68e-20 
C9187 VCC.n5240 VSS 4.12e-20 
C9188 VCC.n5241 VSS 4.12e-20 
C9189 VCC.n5242 VSS 3.91e-20 
C9190 VCC.n5243 VSS 4.53e-20 
C9191 VCC.n5244 VSS 4.53e-20 
C9192 VCC.n5245 VSS 1.05e-19 
C9193 VCC.n5246 VSS 1.05e-19 
C9194 VCC.n5247 VSS 4.32e-20 
C9195 VCC.n5248 VSS 3.7e-20 
C9196 VCC.n5249 VSS 2.68e-20 
C9197 VCC.n5250 VSS 2.68e-20 
C9198 VCC.n5251 VSS 6.79e-20 
C9199 VCC.n5252 VSS 9.26e-20 
C9200 VCC.n5253 VSS 1.83e-19 
C9201 VCC.n5254 VSS 7.95e-19 
C9202 VCC.n5255 VSS 5.2e-19 
C9203 VCC.n5256 VSS 1.3e-19 
C9204 VCC.n5257 VSS 3e-20 
C9205 VCC.n5258 VSS 3.5e-20 
C9206 VCC.n5259 VSS 5.97e-20 
C9207 VCC.n5260 VSS 7.41e-20 
C9208 VCC.n5261 VSS 5.15e-20 
C9209 VCC.n5262 VSS 5.15e-20 
C9210 VCC.n5263 VSS 3.09e-20 
C9211 VCC.n5264 VSS 3.09e-20 
C9212 VCC.n5265 VSS 3.7e-20 
C9213 VCC.n5266 VSS 2.68e-20 
C9214 VCC.n5267 VSS 3.91e-20 
C9215 VCC.n5268 VSS 1.17e-19 
C9216 VCC.n5269 VSS 1.38e-19 
C9217 VCC.n5270 VSS 7e-20 
C9218 VCC.n5271 VSS 4.73e-20 
C9219 VCC.n5272 VSS 3.5e-20 
C9220 VCC.n5273 VSS 3.5e-20 
C9221 VCC.n5274 VSS 3.5e-20 
C9222 VCC.n5275 VSS 4.53e-20 
C9223 VCC.n5276 VSS 1.18e-19 
C9224 VCC.n5277 VSS 5.12e-19 
C9225 VCC.n5278 VSS 1.3e-19 
C9226 VCC.n5279 VSS 1.61e-19 
C9227 VCC.n5280 VSS 9.9e-20 
C9228 VCC.n5281 VSS 0.00243f 
C9229 VCC.n5282 VSS 2.26e-20 
C9230 VCC.n5283 VSS 4.13e-19 
C9231 VCC.n5284 VSS 3.5e-20 
C9232 VCC.n5285 VSS 3.5e-20 
C9233 VCC.n5286 VSS 2.47e-20 
C9234 VCC.n5287 VSS 2.06e-20 
C9235 VCC.n5288 VSS 6.17e-20 
C9236 VCC.n5289 VSS 6.17e-20 
C9237 VCC.n5290 VSS 4.73e-20 
C9238 VCC.n5291 VSS 4.73e-20 
C9239 VCC.n5292 VSS 2.88e-20 
C9240 VCC.n5293 VSS 1.44e-20 
C9241 VCC.n5294 VSS 1.65e-20 
C9242 VCC.n5295 VSS 1.54e-19 
C9243 VCC.n5296 VSS 1.54e-19 
C9244 VCC.n5297 VSS 1.65e-20 
C9245 VCC.n5298 VSS 3.09e-20 
C9246 VCC.t126 VSS 1.55e-19 
C9247 VCC.n5299 VSS 0.00102f 
C9248 VCC.n5300 VSS 2.73e-19 
C9249 VCC.n5301 VSS 0.00136f 
C9250 VCC.n5302 VSS 2.73e-19 
C9251 VCC.n5303 VSS 0.00181f 
C9252 VCC.n5304 VSS 5.76e-20 
C9253 VCC.n5305 VSS 1.54e-19 
C9254 VCC.n5306 VSS 1.65e-20 
C9255 VCC.n5307 VSS 2.88e-20 
C9256 VCC.n5308 VSS 2.47e-20 
C9257 VCC.n5309 VSS 6.17e-20 
C9258 VCC.n5310 VSS 4.73e-20 
C9259 VCC.n5311 VSS 4.73e-20 
C9260 VCC.n5312 VSS 5.15e-20 
C9261 VCC.n5313 VSS 3.5e-20 
C9262 VCC.n5314 VSS 7.41e-20 
C9263 VCC.n5315 VSS 3.7e-20 
C9264 VCC.n5316 VSS 2.26e-20 
C9265 VCC.n5317 VSS 6.17e-20 
C9266 VCC.n5318 VSS 4.73e-20 
C9267 VCC.n5319 VSS 3.5e-20 
C9268 VCC.n5320 VSS 2.88e-20 
C9269 VCC.n5321 VSS 3.4e-19 
C9270 VCC.n5322 VSS 1.15e-19 
C9271 VCC.n5323 VSS 3.98e-19 
C9272 VCC.t233 VSS 4.05e-19 
C9273 VCC.n5324 VSS 1.22e-19 
C9274 VCC.n5325 VSS 1.3e-19 
C9275 VCC.n5326 VSS 3e-20 
C9276 VCC.n5327 VSS 3.5e-20 
C9277 VCC.n5328 VSS 3.5e-20 
C9278 VCC.n5329 VSS 4.73e-20 
C9279 VCC.n5330 VSS 2.47e-20 
C9280 VCC.n5331 VSS 1.23e-20 
C9281 VCC.n5332 VSS 1.65e-20 
C9282 VCC.n5333 VSS 2.47e-20 
C9283 VCC.n5334 VSS 5.76e-20 
C9284 VCC.n5335 VSS 1.38e-19 
C9285 VCC.n5336 VSS 7e-20 
C9286 VCC.n5337 VSS 3.7e-20 
C9287 VCC.n5338 VSS 2.47e-20 
C9288 VCC.n5339 VSS 3.7e-20 
C9289 VCC.n5340 VSS 1.85e-20 
C9290 VCC.n5341 VSS 3.09e-20 
C9291 VCC.n5342 VSS 5.35e-20 
C9292 VCC.n5343 VSS 4.73e-20 
C9293 VCC.n5344 VSS 5.35e-20 
C9294 VCC.n5345 VSS 7.41e-20 
C9295 VCC.n5346 VSS 5.76e-20 
C9296 VCC.n5347 VSS 9.53e-20 
C9297 VCC.n5348 VSS 4.13e-19 
C9298 VCC.n5349 VSS 1.3e-19 
C9299 VCC.n5350 VSS 5.2e-19 
C9300 VCC.n5351 VSS 1.2e-19 
C9301 VCC.n5352 VSS 4.73e-20 
C9302 VCC.n5353 VSS 2.68e-20 
C9303 VCC.n5354 VSS 3.5e-20 
C9304 VCC.n5355 VSS 3.5e-20 
C9305 VCC.n5356 VSS 2.68e-20 
C9306 VCC.n5357 VSS 2.68e-20 
C9307 VCC.n5358 VSS 4.32e-20 
C9308 VCC.n5359 VSS 4.32e-20 
C9309 VCC.n5360 VSS 4.32e-20 
C9310 VCC.n5361 VSS 2.88e-20 
C9311 VCC.n5362 VSS 3.5e-20 
C9312 VCC.n5363 VSS 2.68e-20 
C9313 VCC.n5364 VSS 7.82e-20 
C9314 VCC.n5365 VSS 4.73e-20 
C9315 VCC.n5366 VSS 4.73e-20 
C9316 VCC.n5367 VSS 1.05e-19 
C9317 VCC.n5368 VSS 1.05e-19 
C9318 VCC.n5369 VSS 4.53e-20 
C9319 VCC.n5370 VSS 2.68e-20 
C9320 VCC.n5371 VSS 2.68e-20 
C9321 VCC.n5372 VSS 6.59e-20 
C9322 VCC.n5373 VSS 9.26e-20 
C9323 VCC.n5374 VSS 6.59e-20 
C9324 VCC.n5375 VSS 2.47e-20 
C9325 VCC.n5376 VSS 2.47e-20 
C9326 VCC.n5377 VSS 2.88e-20 
C9327 VCC.n5378 VSS 3.5e-20 
C9328 VCC.n5379 VSS 3.5e-20 
C9329 VCC.n5380 VSS 4.53e-20 
C9330 VCC.n5381 VSS 1.2e-19 
C9331 VCC.n5382 VSS 5.2e-19 
C9332 VCC.n5383 VSS 1.3e-19 
C9333 VCC.n5384 VSS 4.13e-19 
C9334 VCC.n5385 VSS 9.53e-20 
C9335 VCC.n5386 VSS 5.97e-20 
C9336 VCC.n5387 VSS 7.41e-20 
C9337 VCC.n5388 VSS 5.35e-20 
C9338 VCC.n5389 VSS 5.15e-20 
C9339 VCC.n5390 VSS 3.09e-20 
C9340 VCC.n5391 VSS 3.09e-20 
C9341 VCC.n5392 VSS 3.91e-20 
C9342 VCC.n5393 VSS 2.47e-20 
C9343 VCC.n5394 VSS 3.7e-20 
C9344 VCC.n5395 VSS 1.17e-19 
C9345 VCC.n5396 VSS 1.38e-19 
C9346 VCC.n5397 VSS 7.2e-20 
C9347 VCC.n5398 VSS 4.73e-20 
C9348 VCC.n5399 VSS 3.5e-20 
C9349 VCC.n5400 VSS 3.5e-20 
C9350 VCC.n5401 VSS 4.53e-20 
C9351 VCC.n5402 VSS 5.97e-20 
C9352 VCC.n5403 VSS 3.5e-20 
C9353 VCC.n5404 VSS 3e-20 
C9354 VCC.n5405 VSS 1.3e-19 
C9355 VCC.n5406 VSS 1.53e-19 
C9356 VCC.t161 VSS 4.05e-19 
C9357 VCC.n5407 VSS 2.06e-19 
C9358 VCC.n5408 VSS 1.35e-19 
C9359 VCC.n5409 VSS 9.67e-20 
C9360 VCC.n5410 VSS 3.35e-20 
C9361 VCC.n5411 VSS 3.5e-20 
C9362 VCC.n5412 VSS 2.36e-19 
C9363 VCC.n5413 VSS 0.0023f 
C9364 VCC.t222 VSS 0.0031f 
C9365 VCC.t7 VSS 0.00366f 
C9366 VCC.t225 VSS 0.00365f 
C9367 VCC.t10 VSS 0.00386f 
C9368 VCC.n5414 VSS 0.00569f 
C9369 VCC.n5415 VSS 1.3e-19 
C9370 VCC.n5416 VSS 3.67e-19 
C9371 VCC.n5417 VSS 1.15e-19 
C9372 VCC.n5418 VSS 3.38e-19 
C9373 VCC.n5419 VSS 3.5e-20 
C9374 VCC.n5420 VSS 3.5e-20 
C9375 VCC.n5421 VSS 2.68e-20 
C9376 VCC.n5422 VSS 2.06e-20 
C9377 VCC.n5423 VSS 6.38e-20 
C9378 VCC.n5424 VSS 5.97e-20 
C9379 VCC.n5425 VSS 4.73e-20 
C9380 VCC.n5426 VSS 4.73e-20 
C9381 VCC.n5427 VSS 3.09e-20 
C9382 VCC.n5428 VSS 1.23e-20 
C9383 VCC.n5429 VSS 1.65e-20 
C9384 VCC.n5430 VSS 1.54e-19 
C9385 VCC.n5431 VSS 1.54e-19 
C9386 VCC.n5432 VSS 1.65e-20 
C9387 VCC.n5433 VSS 3.29e-20 
C9388 VCC.t162 VSS 1.67e-19 
C9389 VCC.n5434 VSS 0.00101f 
C9390 VCC.n5435 VSS 2.71e-19 
C9391 VCC.n5436 VSS 7.46e-19 
C9392 VCC.n5437 VSS 0.00333f 
C9393 VCC.n5438 VSS 2.46e-19 
C9394 VCC.n5439 VSS 3.02e-19 
C9395 VCC.n5440 VSS 3.7e-20 
C9396 VCC.n5441 VSS 5.15e-20 
C9397 VCC.n5442 VSS 6.38e-20 
C9398 VCC.n5443 VSS 4.73e-20 
C9399 VCC.n5444 VSS 4.73e-20 
C9400 VCC.n5445 VSS 2.68e-20 
C9401 VCC.n5446 VSS 3.29e-20 
C9402 VCC.n5447 VSS 1.65e-20 
C9403 VCC.n5448 VSS 1.54e-19 
C9404 VCC.n5449 VSS 1.54e-19 
C9405 VCC.n5450 VSS 5.56e-20 
C9406 VCC.n5451 VSS 2.88e-20 
C9407 VCC.n5452 VSS 1.65e-20 
C9408 VCC.n5453 VSS 3.09e-20 
C9409 VCC.n5454 VSS 4.73e-20 
C9410 VCC.n5455 VSS 4.73e-20 
C9411 VCC.n5456 VSS 4.32e-20 
C9412 VCC.n5457 VSS 1.17e-19 
C9413 VCC.n5458 VSS 3.33e-19 
C9414 VCC.n5459 VSS 1.35e-19 
C9415 VCC.n5460 VSS 4.37e-19 
C9416 VCC.n5461 VSS 5.24e-19 
C9417 VCC.n5462 VSS 1.36e-19 
C9418 VCC.n5463 VSS 1.01e-19 
C9419 VCC.n5464 VSS 1.05e-19 
C9420 VCC.n5465 VSS 2.06e-20 
C9421 VCC.n5466 VSS 2.26e-20 
C9422 VCC.n5467 VSS 3.7e-20 
C9423 VCC.n5468 VSS 5.15e-20 
C9424 VCC.n5469 VSS 1.38e-19 
C9425 VCC.n5470 VSS 3.91e-20 
C9426 VCC.n5471 VSS 2.88e-20 
C9427 VCC.n5472 VSS 4.32e-20 
C9428 VCC.n5473 VSS 1.17e-19 
C9429 VCC.n5474 VSS 3.7e-20 
C9430 VCC.n5475 VSS 3.91e-20 
C9431 VCC.n5476 VSS 3.5e-20 
C9432 VCC.n5477 VSS 1.65e-20 
C9433 VCC.n5478 VSS 8.23e-21 
C9434 VCC.n5479 VSS 3.5e-20 
C9435 VCC.n5480 VSS 3.5e-20 
C9436 VCC.n5481 VSS 1.4e-19 
C9437 VCC.n5482 VSS 5.4e-19 
C9438 VCC.n5483 VSS 8.42e-19 
C9439 VCC.n5484 VSS 5.4e-19 
C9440 VCC.n5485 VSS 1.4e-19 
C9441 VCC.n5486 VSS 1.4e-19 
C9442 VCC.n5487 VSS 2.18e-19 
C9443 VCC.n5488 VSS 7.82e-20 
C9444 VCC.n5489 VSS 4.32e-20 
C9445 VCC.n5490 VSS 4.32e-20 
C9446 VCC.n5491 VSS 1.05e-19 
C9447 VCC.n5492 VSS 1.05e-19 
C9448 VCC.n5493 VSS 4.32e-20 
C9449 VCC.n5494 VSS 3.7e-20 
C9450 VCC.n5495 VSS 2.68e-20 
C9451 VCC.n5496 VSS 5.76e-20 
C9452 VCC.n5497 VSS 6.38e-20 
C9453 VCC.n5498 VSS 3.5e-20 
C9454 VCC.n5499 VSS 3.5e-20 
C9455 VCC.n5500 VSS 1.17e-19 
C9456 VCC.n5501 VSS 1.38e-19 
C9457 VCC.n5502 VSS 5.15e-20 
C9458 VCC.n5503 VSS 1.05e-19 
C9459 VCC.n5504 VSS 2.26e-20 
C9460 VCC.n5505 VSS 5.76e-20 
C9461 VCC.n5506 VSS 3.7e-20 
C9462 VCC.n5507 VSS 3.7e-20 
C9463 VCC.n5508 VSS 3.09e-20 
C9464 VCC.n5509 VSS 1.85e-20 
C9465 VCC.n5510 VSS 1.65e-20 
C9466 VCC.n5511 VSS 8.23e-21 
C9467 VCC.n5512 VSS 1.13e-19 
C9468 VCC.n5513 VSS 3.33e-19 
C9469 VCC.t116 VSS 4.21e-19 
C9470 VCC.n5514 VSS 2.06e-19 
C9471 VCC.n5515 VSS 1.35e-19 
C9472 VCC.n5516 VSS 3.5e-20 
C9473 VCC.n5517 VSS 3.5e-20 
C9474 VCC.n5518 VSS 3.5e-20 
C9475 VCC.n5519 VSS 1.03e-20 
C9476 VCC.n5520 VSS 2.68e-20 
C9477 VCC.n5521 VSS 3.09e-20 
C9478 VCC.n5522 VSS 2.68e-20 
C9479 VCC.n5523 VSS 1.65e-20 
C9480 VCC.n5524 VSS 1.54e-19 
C9481 VCC.n5525 VSS 1.54e-19 
C9482 VCC.n5526 VSS 1.65e-20 
C9483 VCC.t117 VSS 1.56e-19 
C9484 VCC.n5527 VSS 7.62e-19 
C9485 VCC.n5528 VSS 1.23e-20 
C9486 VCC.n5529 VSS 2.47e-20 
C9487 VCC.n5530 VSS 4.73e-20 
C9488 VCC.n5531 VSS 6.59e-20 
C9489 VCC.n5532 VSS 5.15e-20 
C9490 VCC.n5533 VSS 2.47e-20 
C9491 VCC.n5534 VSS 7.41e-20 
C9492 VCC.n5535 VSS 9.47e-20 
C9493 VCC.n5536 VSS 1.32e-19 
C9494 VCC.n5537 VSS 7.71e-19 
C9495 VCC.n5538 VSS 9.83e-19 
C9496 VCC.n5539 VSS 2.36e-19 
C9497 VCC.n5540 VSS 3.21e-19 
C9498 VCC.n5541 VSS 2.61e-19 
C9499 VCC.n5542 VSS 0.00189f 
C9500 VCC.n5543 VSS 5.76e-20 
C9501 VCC.n5544 VSS 2.88e-20 
C9502 VCC.n5545 VSS 3.5e-20 
C9503 VCC.n5546 VSS 9.83e-19 
C9504 VCC.n5547 VSS 9.47e-20 
C9505 VCC.n5548 VSS 1.17e-19 
C9506 VCC.n5549 VSS 2.06e-19 
C9507 VCC.n5550 VSS 1.36e-19 
C9508 VCC.n5551 VSS 1.01e-19 
C9509 VCC.n5552 VSS 3.5e-20 
C9510 VCC.n5553 VSS 3.09e-20 
C9511 VCC.n5554 VSS 3.29e-20 
C9512 VCC.n5555 VSS 3.29e-20 
C9513 VCC.n5556 VSS 4.73e-20 
C9514 VCC.n5557 VSS 1.44e-20 
C9515 VCC.n5558 VSS 3.5e-20 
C9516 VCC.n5559 VSS 7.41e-20 
C9517 VCC.n5560 VSS 2.47e-20 
C9518 VCC.t9 VSS 1.56e-19 
C9519 VCC.n5561 VSS 5.76e-20 
C9520 VCC.n5562 VSS 2.06e-20 
C9521 VCC.n5563 VSS 5.76e-20 
C9522 VCC.n5564 VSS 3.7e-20 
C9523 VCC.n5565 VSS 4.32e-20 
C9524 VCC.n5566 VSS 2.68e-20 
C9525 VCC.n5567 VSS 3.91e-20 
C9526 VCC.n5568 VSS 6.38e-20 
C9527 VCC.n5569 VSS 1.85e-20 
C9528 VCC.n5570 VSS 3.5e-20 
C9529 VCC.n5571 VSS 3.09e-20 
C9530 VCC.n5572 VSS 3.7e-20 
C9531 VCC.n5573 VSS 3.09e-20 
C9532 VCC.n5574 VSS 2.26e-20 
C9533 VCC.n5575 VSS 1.05e-19 
C9534 VCC.n5576 VSS 3.5e-20 
C9535 VCC.n5577 VSS 3.5e-20 
C9536 VCC.n5578 VSS 8.42e-19 
C9537 VCC.n5579 VSS 2.18e-19 
C9538 VCC.n5580 VSS 1.4e-19 
C9539 VCC.n5581 VSS 4.32e-20 
C9540 VCC.n5582 VSS 7.82e-20 
C9541 VCC.n5583 VSS 5.76e-20 
C9542 VCC.n5584 VSS 2.68e-20 
C9543 VCC.n5585 VSS 4.32e-20 
C9544 VCC.n5586 VSS 3.91e-20 
C9545 VCC.n5587 VSS 3.7e-20 
C9546 VCC.n5588 VSS 3.7e-20 
C9547 VCC.n5589 VSS 5.76e-20 
C9548 VCC.n5590 VSS 4.73e-20 
C9549 VCC.n5591 VSS 3.5e-20 
C9550 VCC.t246 VSS 1.56e-19 
C9551 VCC.n5592 VSS 7.97e-19 
C9552 VCC.n5593 VSS 3.09e-20 
C9553 VCC.n5594 VSS 1.01e-19 
C9554 VCC.n5595 VSS 3.5e-20 
C9555 VCC.n5596 VSS 1.36e-19 
C9556 VCC.n5597 VSS 3.5e-20 
C9557 VCC.n5598 VSS 3.33e-19 
C9558 VCC.n5599 VSS 1.17e-19 
C9559 VCC.n5600 VSS 1.09e-19 
C9560 VCC.n5601 VSS 3.5e-20 
C9561 VCC.n5602 VSS 4.73e-20 
C9562 VCC.n5603 VSS 5.56e-20 
C9563 VCC.n5604 VSS 2.88e-20 
C9564 VCC.n5605 VSS 2.26e-20 
C9565 VCC.n5606 VSS 5.76e-20 
C9566 VCC.n5607 VSS 2.68e-20 
C9567 VCC.n5608 VSS 2.68e-20 
C9568 VCC.n5609 VSS 1.9e-19 
C9569 VCC.n5610 VSS 5.76e-20 
C9570 VCC.n5611 VSS 2.68e-20 
C9571 VCC.n5612 VSS 2.68e-20 
C9572 VCC.n5613 VSS 2.68e-20 
C9573 VCC.n5614 VSS 5.76e-20 
C9574 VCC.n5615 VSS 2.26e-20 
C9575 VCC.n5616 VSS 3.09e-20 
C9576 VCC.n5617 VSS 2.26e-20 
C9577 VCC.n5618 VSS 5.15e-20 
C9578 VCC.n5619 VSS 4.73e-20 
C9579 VCC.n5620 VSS 3.7e-20 
C9580 VCC.n5621 VSS 3.5e-20 
C9581 VCC.n5622 VSS 7.41e-20 
C9582 VCC.n5623 VSS 1.91e-19 
C9583 VCC.n5624 VSS 9.88e-20 
C9584 VCC.n5625 VSS 3e-20 
C9585 VCC.n5626 VSS 5.12e-19 
C9586 VCC.n5627 VSS 1.18e-19 
C9587 VCC.n5628 VSS 3.5e-20 
C9588 VCC.n5629 VSS 3.5e-20 
C9589 VCC.n5630 VSS 5.15e-20 
C9590 VCC.n5631 VSS 4.32e-20 
C9591 VCC.n5632 VSS 2.68e-20 
C9592 VCC.n5633 VSS 3.91e-20 
C9593 VCC.n5634 VSS 1.44e-20 
C9594 VCC.n5635 VSS 3.5e-20 
C9595 VCC.n5636 VSS 3e-20 
C9596 VCC.n5637 VSS 7.95e-19 
C9597 VCC.n5638 VSS 1.83e-19 
C9598 VCC.n5639 VSS 2.88e-20 
C9599 VCC.n5640 VSS 2.68e-20 
C9600 VCC.n5641 VSS 2.68e-20 
C9601 VCC.n5642 VSS 2.68e-20 
C9602 VCC.n5643 VSS 4.53e-20 
C9603 VCC.n5644 VSS 3.7e-20 
C9604 VCC.n5645 VSS 7.82e-20 
C9605 VCC.n5646 VSS 1.17e-19 
C9606 VCC.n5647 VSS 3.91e-20 
C9607 VCC.n5648 VSS 1.65e-20 
C9608 VCC.n5649 VSS 2.68e-20 
C9609 VCC.n5650 VSS 3.5e-20 
C9610 VCC.n5651 VSS 3e-20 
C9611 VCC.n5652 VSS 5.12e-19 
C9612 VCC.n5653 VSS 1.18e-19 
C9613 VCC.n5654 VSS 3.5e-20 
C9614 VCC.n5655 VSS 3.5e-20 
C9615 VCC.t192 VSS 1.55e-19 
C9616 VCC.n5656 VSS 7.57e-19 
C9617 VCC.n5657 VSS 4.73e-20 
C9618 VCC.n5658 VSS 1.54e-19 
C9619 VCC.n5659 VSS 2.88e-20 
C9620 VCC.n5660 VSS 2.88e-20 
C9621 VCC.n5661 VSS 3.5e-20 
C9622 VCC.n5662 VSS 5.76e-20 
C9623 VCC.n5663 VSS 9.88e-20 
C9624 VCC.n5664 VSS 1.3e-19 
C9625 VCC.n5665 VSS 3e-20 
C9626 VCC.t193 VSS 0.005f 
C9627 VCC.t164 VSS 0.00453f 
C9628 VCC.n5666 VSS 0.00229f 
C9629 VCC.n5667 VSS 1.91e-19 
C9630 VCC.n5668 VSS 3.5e-20 
C9631 VCC.n5669 VSS 3.14e-19 
C9632 VCC.n5670 VSS 3.5e-20 
C9633 VCC.n5671 VSS 2.47e-20 
C9634 VCC.n5672 VSS 5.76e-20 
C9635 VCC.n5673 VSS 2.47e-20 
C9636 VCC.n5674 VSS 8.23e-21 
C9637 VCC.n5675 VSS 2.88e-20 
C9638 VCC.n5676 VSS 5.76e-20 
C9639 VCC.n5677 VSS 2.47e-20 
C9640 VCC.n5678 VSS 2.88e-20 
C9641 VCC.n5679 VSS 2.47e-20 
C9642 VCC.n5680 VSS 5.15e-20 
C9643 VCC.n5681 VSS 4.73e-20 
C9644 VCC.n5682 VSS 3.7e-20 
C9645 VCC.n5683 VSS 3.5e-20 
C9646 VCC.n5684 VSS 7.41e-20 
C9647 VCC.t259 VSS 6.42e-19 
C9648 VCC.n5685 VSS 3e-20 
C9649 VCC.n5686 VSS 5.97e-20 
C9650 VCC.n5687 VSS 4.13e-19 
C9651 VCC.n5688 VSS 9.53e-20 
C9652 VCC.n5689 VSS 3.5e-20 
C9653 VCC.n5690 VSS 3.5e-20 
C9654 VCC.n5691 VSS 5.35e-20 
C9655 VCC.n5692 VSS 4.32e-20 
C9656 VCC.n5693 VSS 2.68e-20 
C9657 VCC.n5694 VSS 3.7e-20 
C9658 VCC.n5695 VSS 1.65e-20 
C9659 VCC.n5696 VSS 4.53e-20 
C9660 VCC.n5697 VSS 1.2e-19 
C9661 VCC.n5698 VSS 5.2e-19 
C9662 VCC.n5699 VSS 1.2e-19 
C9663 VCC.n5700 VSS 6.38e-20 
C9664 VCC.n5701 VSS 2.47e-20 
C9665 VCC.n5702 VSS 4.53e-20 
C9666 VCC.n5703 VSS 3.5e-20 
C9667 VCC.n5704 VSS 3.5e-20 
C9668 VCC.n5705 VSS 2.68e-20 
C9669 VCC.n5706 VSS 2.68e-20 
C9670 VCC.n5707 VSS 2.47e-20 
C9671 VCC.n5708 VSS 4.53e-20 
C9672 VCC.n5709 VSS 2.68e-20 
C9673 VCC.n5710 VSS 4.32e-20 
C9674 VCC.n5711 VSS 2.68e-20 
C9675 VCC.n5712 VSS 3.91e-20 
C9676 VCC.n5713 VSS 2.88e-20 
C9677 VCC.n5714 VSS 4.73e-20 
C9678 VCC.n5715 VSS 3.7e-20 
C9679 VCC.n5716 VSS 3.7e-20 
C9680 VCC.n5717 VSS 3.5e-20 
C9681 VCC.n5718 VSS 5.76e-20 
C9682 VCC.n5719 VSS 4.73e-20 
C9683 VCC.n5720 VSS 3.09e-20 
C9684 VCC.n5721 VSS 3.5e-20 
C9685 VCC.n5722 VSS 3.5e-20 
C9686 VCC.n5723 VSS 3.5e-20 
C9687 VCC.n5724 VSS 1.18e-19 
C9688 VCC.n5725 VSS 3e-20 
C9689 VCC.n5726 VSS 1.15e-19 
C9690 VCC.n5727 VSS 9.88e-20 
C9691 VCC.n5728 VSS 5.76e-20 
C9692 VCC.n5729 VSS 3.5e-20 
C9693 VCC.n5730 VSS 3.09e-20 
C9694 VCC.n5731 VSS 3.09e-20 
C9695 VCC.n5732 VSS 2.26e-20 
C9696 VCC.n5733 VSS 5.76e-20 
C9697 VCC.n5734 VSS 2.68e-20 
C9698 VCC.n5735 VSS 2.68e-20 
C9699 VCC.n5736 VSS 0.00185f 
C9700 VCC.n5737 VSS 2.72e-19 
C9701 VCC.n5738 VSS 2.26e-20 
C9702 VCC.n5739 VSS 1.87e-19 
C9703 VCC.n5740 VSS 3.5e-20 
C9704 VCC.n5741 VSS 2.68e-20 
C9705 VCC.n5742 VSS 5.97e-20 
C9706 VCC.n5743 VSS 4.73e-20 
C9707 VCC.n5744 VSS 4.73e-20 
C9708 VCC.n5745 VSS 5.15e-20 
C9709 VCC.n5746 VSS 7.41e-20 
C9710 VCC.n5747 VSS 3.7e-20 
C9711 VCC.n5748 VSS 2.26e-20 
C9712 VCC.n5749 VSS 6.38e-20 
C9713 VCC.n5750 VSS 4.73e-20 
C9714 VCC.n5751 VSS 3.29e-20 
C9715 VCC.n5752 VSS 3.5e-20 
C9716 VCC.n5753 VSS 3e-20 
C9717 VCC.t52 VSS 0.005f 
C9718 VCC.t81 VSS 0.00453f 
C9719 VCC.n5754 VSS 0.00228f 
C9720 VCC.n5755 VSS 1.3e-19 
C9721 VCC.t53 VSS 4.05e-19 
C9722 VCC.n5756 VSS 4.05e-19 
C9723 VCC.n5757 VSS 1.15e-19 
C9724 VCC.n5758 VSS 3.36e-19 
C9725 VCC.n5759 VSS 6.17e-21 
C9726 VCC.n5760 VSS 3.12e-19 
C9727 VCC.n5761 VSS 1.65e-20 
C9728 VCC.n5762 VSS 1.54e-19 
C9729 VCC.n5763 VSS 1.54e-19 
C9730 VCC.n5764 VSS 1.65e-20 
C9731 VCC.n5765 VSS 1.03e-20 
C9732 VCC.n5766 VSS 3.5e-20 
C9733 VCC.n5767 VSS 2.26e-20 
C9734 VCC.n5768 VSS 4.73e-20 
C9735 VCC.n5769 VSS 3.5e-20 
C9736 VCC.n5770 VSS 3e-20 
C9737 VCC.n5771 VSS 1.3e-19 
C9738 VCC.n5772 VSS 5.12e-19 
C9739 VCC.n5773 VSS 1.3e-19 
C9740 VCC.n5774 VSS 4.13e-19 
C9741 VCC.n5775 VSS 9.53e-20 
C9742 VCC.n5776 VSS 5.76e-20 
C9743 VCC.n5777 VSS 7.41e-20 
C9744 VCC.n5778 VSS 5.56e-20 
C9745 VCC.t54 VSS 1.55e-19 
C9746 VCC.n5779 VSS 3.91e-20 
C9747 VCC.n5780 VSS 3.91e-20 
C9748 VCC.n5781 VSS 1.85e-20 
C9749 VCC.n5782 VSS 7.55e-19 
C9750 VCC.n5783 VSS 4.94e-20 
C9751 VCC.n5784 VSS 5.15e-20 
C9752 VCC.n5785 VSS 7.2e-20 
C9753 VCC.n5786 VSS 1.38e-19 
C9754 VCC.n5787 VSS 1.17e-19 
C9755 VCC.n5788 VSS 4.32e-20 
C9756 VCC.n5789 VSS 2.88e-20 
C9757 VCC.n5790 VSS 2.68e-20 
C9758 VCC.n5791 VSS 3.5e-20 
C9759 VCC.n5792 VSS 3.5e-20 
C9760 VCC.n5793 VSS 2.88e-20 
C9761 VCC.n5794 VSS 2.68e-20 
C9762 VCC.n5795 VSS 2.68e-20 
C9763 VCC.n5796 VSS 2.68e-20 
C9764 VCC.n5797 VSS 4.12e-20 
C9765 VCC.n5798 VSS 4.12e-20 
C9766 VCC.n5799 VSS 3.91e-20 
C9767 VCC.n5800 VSS 4.53e-20 
C9768 VCC.n5801 VSS 4.53e-20 
C9769 VCC.n5802 VSS 1.05e-19 
C9770 VCC.n5803 VSS 1.05e-19 
C9771 VCC.n5804 VSS 4.32e-20 
C9772 VCC.n5805 VSS 3.7e-20 
C9773 VCC.n5806 VSS 2.68e-20 
C9774 VCC.n5807 VSS 2.68e-20 
C9775 VCC.n5808 VSS 6.79e-20 
C9776 VCC.n5809 VSS 9.26e-20 
C9777 VCC.n5810 VSS 1.83e-19 
C9778 VCC.n5811 VSS 7.95e-19 
C9779 VCC.n5812 VSS 5.2e-19 
C9780 VCC.n5813 VSS 1.3e-19 
C9781 VCC.n5814 VSS 3e-20 
C9782 VCC.n5815 VSS 3.5e-20 
C9783 VCC.n5816 VSS 5.97e-20 
C9784 VCC.n5817 VSS 7.41e-20 
C9785 VCC.n5818 VSS 5.15e-20 
C9786 VCC.n5819 VSS 5.15e-20 
C9787 VCC.n5820 VSS 3.09e-20 
C9788 VCC.n5821 VSS 3.09e-20 
C9789 VCC.n5822 VSS 3.7e-20 
C9790 VCC.n5823 VSS 2.68e-20 
C9791 VCC.n5824 VSS 3.91e-20 
C9792 VCC.n5825 VSS 1.17e-19 
C9793 VCC.n5826 VSS 1.38e-19 
C9794 VCC.n5827 VSS 7e-20 
C9795 VCC.n5828 VSS 4.73e-20 
C9796 VCC.n5829 VSS 3.5e-20 
C9797 VCC.n5830 VSS 3.5e-20 
C9798 VCC.n5831 VSS 3.5e-20 
C9799 VCC.n5832 VSS 4.53e-20 
C9800 VCC.n5833 VSS 1.18e-19 
C9801 VCC.n5834 VSS 5.12e-19 
C9802 VCC.n5835 VSS 1.3e-19 
C9803 VCC.n5836 VSS 1.61e-19 
C9804 VCC.n5837 VSS 9.9e-20 
C9805 VCC.n5838 VSS 0.00243f 
C9806 VCC.n5839 VSS 2.26e-20 
C9807 VCC.n5840 VSS 4.13e-19 
C9808 VCC.n5841 VSS 3.5e-20 
C9809 VCC.n5842 VSS 3.5e-20 
C9810 VCC.n5843 VSS 2.47e-20 
C9811 VCC.n5844 VSS 2.06e-20 
C9812 VCC.n5845 VSS 6.17e-20 
C9813 VCC.n5846 VSS 6.17e-20 
C9814 VCC.n5847 VSS 4.73e-20 
C9815 VCC.n5848 VSS 4.73e-20 
C9816 VCC.n5849 VSS 2.88e-20 
C9817 VCC.n5850 VSS 1.44e-20 
C9818 VCC.n5851 VSS 1.65e-20 
C9819 VCC.n5852 VSS 1.54e-19 
C9820 VCC.n5853 VSS 1.54e-19 
C9821 VCC.n5854 VSS 1.65e-20 
C9822 VCC.n5855 VSS 3.09e-20 
C9823 VCC.t260 VSS 1.55e-19 
C9824 VCC.n5856 VSS 0.00102f 
C9825 VCC.n5857 VSS 2.73e-19 
C9826 VCC.n5858 VSS 0.00136f 
C9827 VCC.n5859 VSS 2.73e-19 
C9828 VCC.n5860 VSS 0.00181f 
C9829 VCC.n5861 VSS 5.76e-20 
C9830 VCC.n5862 VSS 1.54e-19 
C9831 VCC.n5863 VSS 1.65e-20 
C9832 VCC.n5864 VSS 6.17e-20 
C9833 VCC.n5865 VSS 2.47e-20 
C9834 VCC.n5866 VSS 4.73e-20 
C9835 VCC.n5867 VSS 4.73e-20 
C9836 VCC.n5868 VSS 5.15e-20 
C9837 VCC.n5869 VSS 3.5e-20 
C9838 VCC.n5870 VSS 7.41e-20 
C9839 VCC.n5871 VSS 3.7e-20 
C9840 VCC.n5872 VSS 2.26e-20 
C9841 VCC.n5873 VSS 6.17e-20 
C9842 VCC.n5874 VSS 4.73e-20 
C9843 VCC.n5875 VSS 2.88e-20 
C9844 VCC.n5876 VSS 2.88e-20 
C9845 VCC.n5877 VSS 3.4e-19 
C9846 VCC.n5878 VSS 1.15e-19 
C9847 VCC.n5879 VSS 3.98e-19 
C9848 VCC.t191 VSS 4.05e-19 
C9849 VCC.n5880 VSS 1.22e-19 
C9850 VCC.n5881 VSS 1.3e-19 
C9851 VCC.n5882 VSS 3e-20 
C9852 VCC.n5883 VSS 3.5e-20 
C9853 VCC.n5884 VSS 3.5e-20 
C9854 VCC.n5885 VSS 4.73e-20 
C9855 VCC.n5886 VSS 2.47e-20 
C9856 VCC.n5887 VSS 1.23e-20 
C9857 VCC.n5888 VSS 1.65e-20 
C9858 VCC.n5889 VSS 2.47e-20 
C9859 VCC.n5890 VSS 5.76e-20 
C9860 VCC.n5891 VSS 1.38e-19 
C9861 VCC.n5892 VSS 7e-20 
C9862 VCC.n5893 VSS 3.7e-20 
C9863 VCC.n5894 VSS 2.47e-20 
C9864 VCC.n5895 VSS 3.7e-20 
C9865 VCC.n5896 VSS 1.85e-20 
C9866 VCC.n5897 VSS 3.09e-20 
C9867 VCC.n5898 VSS 5.35e-20 
C9868 VCC.n5899 VSS 4.73e-20 
C9869 VCC.n5900 VSS 5.35e-20 
C9870 VCC.n5901 VSS 7.41e-20 
C9871 VCC.n5902 VSS 5.76e-20 
C9872 VCC.n5903 VSS 9.53e-20 
C9873 VCC.n5904 VSS 4.13e-19 
C9874 VCC.n5905 VSS 1.3e-19 
C9875 VCC.n5906 VSS 5.2e-19 
C9876 VCC.n5907 VSS 1.2e-19 
C9877 VCC.n5908 VSS 4.73e-20 
C9878 VCC.n5909 VSS 2.68e-20 
C9879 VCC.n5910 VSS 3.5e-20 
C9880 VCC.n5911 VSS 3.5e-20 
C9881 VCC.n5912 VSS 2.68e-20 
C9882 VCC.n5913 VSS 2.68e-20 
C9883 VCC.n5914 VSS 4.32e-20 
C9884 VCC.n5915 VSS 4.32e-20 
C9885 VCC.n5916 VSS 4.32e-20 
C9886 VCC.n5917 VSS 2.88e-20 
C9887 VCC.n5918 VSS 3.5e-20 
C9888 VCC.n5919 VSS 2.68e-20 
C9889 VCC.n5920 VSS 7.82e-20 
C9890 VCC.n5921 VSS 4.73e-20 
C9891 VCC.n5922 VSS 4.73e-20 
C9892 VCC.n5923 VSS 1.05e-19 
C9893 VCC.n5924 VSS 1.05e-19 
C9894 VCC.n5925 VSS 4.53e-20 
C9895 VCC.n5926 VSS 2.68e-20 
C9896 VCC.n5927 VSS 2.68e-20 
C9897 VCC.n5928 VSS 6.59e-20 
C9898 VCC.n5929 VSS 9.26e-20 
C9899 VCC.n5930 VSS 6.59e-20 
C9900 VCC.n5931 VSS 2.47e-20 
C9901 VCC.n5932 VSS 2.47e-20 
C9902 VCC.n5933 VSS 2.88e-20 
C9903 VCC.n5934 VSS 3.5e-20 
C9904 VCC.n5935 VSS 3.5e-20 
C9905 VCC.n5936 VSS 4.53e-20 
C9906 VCC.n5937 VSS 1.2e-19 
C9907 VCC.n5938 VSS 5.2e-19 
C9908 VCC.n5939 VSS 1.3e-19 
C9909 VCC.n5940 VSS 4.13e-19 
C9910 VCC.n5941 VSS 9.53e-20 
C9911 VCC.n5942 VSS 5.97e-20 
C9912 VCC.n5943 VSS 7.41e-20 
C9913 VCC.n5944 VSS 5.35e-20 
C9914 VCC.n5945 VSS 5.15e-20 
C9915 VCC.n5946 VSS 3.09e-20 
C9916 VCC.n5947 VSS 3.09e-20 
C9917 VCC.n5948 VSS 3.91e-20 
C9918 VCC.n5949 VSS 2.47e-20 
C9919 VCC.n5950 VSS 3.7e-20 
C9920 VCC.n5951 VSS 1.17e-19 
C9921 VCC.n5952 VSS 1.38e-19 
C9922 VCC.n5953 VSS 7.2e-20 
C9923 VCC.n5954 VSS 4.73e-20 
C9924 VCC.n5955 VSS 3.5e-20 
C9925 VCC.n5956 VSS 3.5e-20 
C9926 VCC.n5957 VSS 4.53e-20 
C9927 VCC.n5958 VSS 5.97e-20 
C9928 VCC.n5959 VSS 3.5e-20 
C9929 VCC.n5960 VSS 3e-20 
C9930 VCC.n5961 VSS 1.3e-19 
C9931 VCC.n5962 VSS 1.53e-19 
C9932 VCC.t242 VSS 4.05e-19 
C9933 VCC.n5963 VSS 1.35e-19 
C9934 VCC.t245 VSS 4.21e-19 
C9935 VCC.n5964 VSS 2.06e-19 
C9936 VCC.n5965 VSS 1.32e-19 
C9937 VCC.n5966 VSS 9.67e-20 
C9938 VCC.n5967 VSS 3.35e-20 
C9939 VCC.n5968 VSS 3.5e-20 
C9940 VCC.n5969 VSS 2.36e-19 
C9941 VCC.n5970 VSS 0.0023f 
C9942 VCC.t244 VSS 0.0031f 
C9943 VCC.t240 VSS 0.00366f 
C9944 VCC.t247 VSS 0.00365f 
C9945 VCC.t239 VSS 0.00386f 
C9946 VCC.n5971 VSS 0.00569f 
C9947 VCC.n5972 VSS 1.3e-19 
C9948 VCC.n5973 VSS 3.67e-19 
C9949 VCC.n5974 VSS 1.15e-19 
C9950 VCC.n5975 VSS 3.38e-19 
C9951 VCC.n5976 VSS 3.5e-20 
C9952 VCC.n5977 VSS 3.5e-20 
C9953 VCC.n5978 VSS 2.68e-20 
C9954 VCC.n5979 VSS 2.06e-20 
C9955 VCC.n5980 VSS 6.38e-20 
C9956 VCC.n5981 VSS 5.97e-20 
C9957 VCC.n5982 VSS 4.73e-20 
C9958 VCC.n5983 VSS 4.73e-20 
C9959 VCC.n5984 VSS 3.09e-20 
C9960 VCC.n5985 VSS 1.23e-20 
C9961 VCC.n5986 VSS 1.65e-20 
C9962 VCC.n5987 VSS 1.54e-19 
C9963 VCC.n5988 VSS 1.54e-19 
C9964 VCC.n5989 VSS 1.65e-20 
C9965 VCC.n5990 VSS 3.29e-20 
C9966 VCC.t243 VSS 1.67e-19 
C9967 VCC.n5991 VSS 0.00101f 
C9968 VCC.n5992 VSS 2.71e-19 
C9969 VCC.n5993 VSS 7.46e-19 
C9970 VCC.n5994 VSS 0.00333f 
C9971 VCC.n5995 VSS 2.46e-19 
C9972 VCC.n5996 VSS 3.02e-19 
C9973 VCC.n5997 VSS 3.7e-20 
C9974 VCC.n5998 VSS 5.15e-20 
C9975 VCC.n5999 VSS 5.97e-20 
C9976 VCC.n6000 VSS 6.38e-20 
C9977 VCC.n6001 VSS 4.73e-20 
C9978 VCC.n6002 VSS 4.73e-20 
C9979 VCC.n6003 VSS 2.68e-20 
C9980 VCC.n6004 VSS 3.29e-20 
C9981 VCC.n6005 VSS 1.65e-20 
C9982 VCC.n6006 VSS 1.54e-19 
C9983 VCC.n6007 VSS 1.54e-19 
C9984 VCC.n6008 VSS 1.65e-20 
C9985 VCC.n6009 VSS 3.09e-20 
C9986 VCC.n6010 VSS 3.09e-20 
C9987 VCC.n6011 VSS 4.73e-20 
C9988 VCC.n6012 VSS 4.32e-20 
C9989 VCC.n6013 VSS 3.5e-20 
C9990 VCC.n6014 VSS 3.5e-20 
C9991 VCC.n6015 VSS 1.35e-19 
C9992 VCC.n6016 VSS 5.24e-19 
C9993 VCC.n6017 VSS 1.4e-19 
C9994 VCC.n6018 VSS 5.4e-19 
C9995 VCC.n6019 VSS 1.35e-19 
C9996 VCC.n6020 VSS 4.37e-19 
C9997 VCC.n6021 VSS 1.13e-19 
C9998 VCC.n6022 VSS 8.23e-21 
C9999 VCC.n6023 VSS 1.65e-20 
C10000 VCC.n6024 VSS 3.5e-20 
C10001 VCC.n6025 VSS 3.91e-20 
C10002 VCC.n6026 VSS 3.09e-20 
C10003 VCC.n6027 VSS 1.85e-20 
C10004 VCC.n6028 VSS 3.5e-20 
C10005 VCC.n6029 VSS 1.05e-19 
C10006 VCC.n6030 VSS 2.06e-20 
C10007 VCC.n6031 VSS 2.26e-20 
C10008 VCC.n6032 VSS 3.7e-20 
C10009 VCC.n6033 VSS 5.15e-20 
C10010 VCC.n6034 VSS 1.38e-19 
C10011 VCC.n6035 VSS 1.17e-19 
C10012 VCC.n6036 VSS 4.32e-20 
C10013 VCC.n6037 VSS 2.88e-20 
C10014 VCC.n6038 VSS 2.68e-20 
C10015 VCC.n6039 VSS 6.59e-20 
C10016 VCC.n6040 VSS 5.56e-20 
C10017 VCC.n6041 VSS 2.68e-20 
C10018 VCC.n6042 VSS 4.32e-20 
C10019 VCC.n6043 VSS 1.05e-19 
C10020 VCC.n6044 VSS 3.09e-20 
C10021 VCC.n6045 VSS 3.7e-20 
C10022 VCC.n6046 VSS 4.32e-20 
C10023 VCC.n6047 VSS 1.05e-19 
C10024 VCC.n6048 VSS 4.53e-20 
C10025 VCC.n6049 VSS 4.53e-20 
C10026 VCC.n6050 VSS 7.82e-20 
C10027 VCC.n6051 VSS 2.18e-19 
C10028 VCC.n6052 VSS 1.4e-19 
C10029 VCC.n6053 VSS 1.4e-19 
C10030 VCC.n6054 VSS 5.4e-19 
C10031 VCC.n6055 VSS 1.35e-19 
C10032 VCC.t8 VSS 4.21e-19 
C10033 VCC.n6056 VSS 3.33e-19 
C10034 VCC.n6057 VSS 1.13e-19 
C10035 VCC.n6058 VSS 8.23e-21 
C10036 VCC.n6059 VSS 1.65e-20 
C10037 VCC.n6060 VSS 3.5e-20 
C10038 VCC.n6061 VSS 3.5e-20 
C10039 VCC.n6062 VSS 3.5e-20 
C10040 VCC.n6063 VSS 1.17e-19 
C10041 VCC.n6064 VSS 1.38e-19 
C10042 VCC.n6065 VSS 5.15e-20 
C10043 VCC.n6066 VSS 4.73e-20 
C10044 VCC.n6067 VSS 7.2e-20 
C10045 VCC.n6068 VSS 2.68e-20 
C10046 VCC.n6069 VSS 1.65e-20 
C10047 VCC.n6070 VSS 1.54e-19 
C10048 VCC.n6071 VSS 1.54e-19 
C10049 VCC.n6072 VSS 1.65e-20 
C10050 VCC.n6073 VSS 2.47e-20 
C10051 VCC.n6074 VSS 1.23e-20 
C10052 VCC.n6075 VSS 7.62e-19 
C10053 VCC.n6076 VSS 4.12e-20 
C10054 VCC.n6077 VSS 5.15e-20 
C10055 VCC.n6078 VSS 6.59e-20 
C10056 VCC.n6079 VSS 5.76e-20 
C10057 VCC.n6080 VSS 4.73e-20 
C10058 VCC.n6081 VSS 2.26e-20 
C10059 VCC.n6082 VSS 2.68e-20 
C10060 VCC.n6083 VSS 1.03e-20 
C10061 VCC.n6084 VSS 3.5e-20 
C10062 VCC.n6085 VSS 3.5e-20 
C10063 VCC.n6086 VSS 1.35e-19 
C10064 VCC.n6087 VSS 4.53e-19 
C10065 VCC.n6088 VSS 7.71e-19 
C10066 VCC.n6089 VSS 1.32e-19 
C10067 VCC.n6090 VSS 3.5e-20 
C10068 VCC.n6091 VSS 3.42e-20 
C10069 VCC.n6092 VSS 2.36e-19 
C10070 VCC.n6093 VSS 3.21e-19 
C10071 VCC.n6094 VSS 2.61e-19 
C10072 VCC.n6095 VSS 0.00189f 
C10073 VCC.n6096 VSS 2.68e-19 
C10074 VCC.n6097 VSS 5.76e-20 
C10075 VCC.n6098 VSS 2.88e-20 
C10076 VCC.n6099 VSS 3.5e-20 
C10077 VCC.n6100 VSS 3.42e-20 
C10078 VCC.n6101 VSS 3.5e-20 
C10079 VCC.n6102 VSS 4.53e-19 
C10080 VCC.n6103 VSS 1.17e-19 
C10081 VCC.n6104 VSS 3.5e-20 
C10082 VCC.n6105 VSS 1.44e-20 
C10083 VCC.n6106 VSS 4.12e-20 
C10084 VCC.n6107 VSS 5.76e-20 
C10085 VCC.n6108 VSS 5.76e-20 
C10086 VCC.n6109 VSS 2.06e-20 
C10087 VCC.n6110 VSS 3.29e-20 
C10088 VCC.n6111 VSS 7.2e-20 
C10089 VCC.n6112 VSS 3.29e-20 
C10090 VCC.n6113 VSS 4.73e-20 
C10091 VCC.n6114 VSS 2.26e-20 
C10092 VCC.n6115 VSS 1.01e-19 
C10093 VCC.n6116 VSS 1.36e-19 
C10094 VCC.n6117 VSS 1.35e-19 
C10095 VCC.n6118 VSS 3.5e-20 
C10096 VCC.n6119 VSS 3.5e-20 
C10097 VCC.n6120 VSS 3.5e-20 
C10098 VCC.n6121 VSS 3.5e-20 
C10099 VCC.n6122 VSS 3.09e-20 
C10100 VCC.n6123 VSS 3.91e-20 
C10101 VCC.n6124 VSS 4.73e-20 
C10102 VCC.n6125 VSS 4.32e-20 
C10103 VCC.n6126 VSS 2.68e-20 
C10104 VCC.n6127 VSS 4.53e-20 
C10105 VCC.n6128 VSS 4.53e-20 
C10106 VCC.n6129 VSS 3.09e-20 
C10107 VCC.n6130 VSS 4.32e-20 
C10108 VCC.n6131 VSS 2.68e-20 
C10109 VCC.n6132 VSS 7.82e-20 
C10110 VCC.n6133 VSS 5.56e-20 
C10111 VCC.n6134 VSS 1.4e-19 
C10112 VCC.n6135 VSS 2.18e-19 
C10113 VCC.n6136 VSS 1.35e-19 
C10114 VCC.n6137 VSS 1.13e-19 
C10115 VCC.n6138 VSS 3.5e-20 
C10116 VCC.n6139 VSS 1.85e-20 
C10117 VCC.n6140 VSS 3.7e-20 
C10118 VCC.n6141 VSS 3.09e-20 
C10119 VCC.n6142 VSS 6.59e-20 
C10120 VCC.n6143 VSS 2.68e-20 
C10121 VCC.n6144 VSS 5.76e-20 
C10122 VCC.n6145 VSS 4.73e-20 
C10123 VCC.n6146 VSS 3.5e-20 
C10124 VCC.t170 VSS 1.56e-19 
C10125 VCC.n6147 VSS 7.97e-19 
C10126 VCC.n6148 VSS 3.09e-20 
C10127 VCC.n6149 VSS 3.5e-20 
C10128 VCC.n6150 VSS 3.5e-20 
C10129 VCC.t169 VSS 4.21e-19 
C10130 VCC.n6151 VSS 1.32e-19 
C10131 VCC.n6152 VSS 1.09e-19 
C10132 VCC.n6153 VSS 3.5e-20 
C10133 VCC.n6154 VSS 3.09e-20 
C10134 VCC.n6155 VSS 5.97e-20 
C10135 VCC.n6156 VSS 2.26e-20 
C10136 VCC.n6157 VSS 5.76e-20 
C10137 VCC.n6158 VSS 2.68e-20 
C10138 VCC.n6159 VSS 2.68e-20 
C10139 VCC.n6160 VSS 1.9e-19 
C10140 VCC.n6161 VSS 5.76e-20 
C10141 VCC.n6162 VSS 2.68e-20 
C10142 VCC.n6163 VSS 2.68e-20 
C10143 VCC.n6164 VSS 2.68e-20 
C10144 VCC.n6165 VSS 5.76e-20 
C10145 VCC.n6166 VSS 2.26e-20 
C10146 VCC.n6167 VSS 3.09e-20 
C10147 VCC.n6168 VSS 2.26e-20 
C10148 VCC.n6169 VSS 5.15e-20 
C10149 VCC.n6170 VSS 4.73e-20 
C10150 VCC.n6171 VSS 3.7e-20 
C10151 VCC.n6172 VSS 3.5e-20 
C10152 VCC.n6173 VSS 7.41e-20 
C10153 VCC.n6174 VSS 1.91e-19 
C10154 VCC.n6175 VSS 9.88e-20 
C10155 VCC.n6176 VSS 3e-20 
C10156 VCC.n6177 VSS 5.12e-19 
C10157 VCC.n6178 VSS 1.18e-19 
C10158 VCC.n6179 VSS 3.5e-20 
C10159 VCC.n6180 VSS 3.5e-20 
C10160 VCC.n6181 VSS 5.15e-20 
C10161 VCC.n6182 VSS 4.32e-20 
C10162 VCC.n6183 VSS 2.68e-20 
C10163 VCC.n6184 VSS 3.91e-20 
C10164 VCC.n6185 VSS 1.44e-20 
C10165 VCC.n6186 VSS 3.5e-20 
C10166 VCC.n6187 VSS 3e-20 
C10167 VCC.n6188 VSS 7.95e-19 
C10168 VCC.n6189 VSS 1.83e-19 
C10169 VCC.n6190 VSS 2.88e-20 
C10170 VCC.n6191 VSS 2.68e-20 
C10171 VCC.n6192 VSS 2.68e-20 
C10172 VCC.n6193 VSS 2.68e-20 
C10173 VCC.n6194 VSS 4.53e-20 
C10174 VCC.n6195 VSS 3.7e-20 
C10175 VCC.n6196 VSS 7.82e-20 
C10176 VCC.n6197 VSS 1.17e-19 
C10177 VCC.n6198 VSS 3.91e-20 
C10178 VCC.n6199 VSS 1.65e-20 
C10179 VCC.n6200 VSS 2.68e-20 
C10180 VCC.n6201 VSS 3.5e-20 
C10181 VCC.n6202 VSS 3e-20 
C10182 VCC.n6203 VSS 5.12e-19 
C10183 VCC.n6204 VSS 1.18e-19 
C10184 VCC.n6205 VSS 3.5e-20 
C10185 VCC.n6206 VSS 3.5e-20 
C10186 VCC.t16 VSS 1.55e-19 
C10187 VCC.n6207 VSS 7.57e-19 
C10188 VCC.n6208 VSS 4.73e-20 
C10189 VCC.n6209 VSS 1.54e-19 
C10190 VCC.n6210 VSS 2.88e-20 
C10191 VCC.n6211 VSS 2.88e-20 
C10192 VCC.n6212 VSS 3.5e-20 
C10193 VCC.n6213 VSS 5.76e-20 
C10194 VCC.n6214 VSS 9.88e-20 
C10195 VCC.n6215 VSS 1.3e-19 
C10196 VCC.n6216 VSS 3e-20 
C10197 VCC.t14 VSS 0.005f 
C10198 VCC.t132 VSS 0.00453f 
C10199 VCC.n6217 VSS 0.00229f 
C10200 VCC.n6218 VSS 1.91e-19 
C10201 VCC.n6219 VSS 3.5e-20 
C10202 VCC.n6220 VSS 3.14e-19 
C10203 VCC.n6221 VSS 2.47e-20 
C10204 VCC.n6222 VSS 5.76e-20 
C10205 VCC.n6223 VSS 2.47e-20 
C10206 VCC.n6224 VSS 8.23e-21 
C10207 VCC.n6225 VSS 2.88e-20 
C10208 VCC.n6226 VSS 5.76e-20 
C10209 VCC.n6227 VSS 2.47e-20 
C10210 VCC.n6228 VSS 2.88e-20 
C10211 VCC.n6229 VSS 2.47e-20 
C10212 VCC.n6230 VSS 5.15e-20 
C10213 VCC.n6231 VSS 4.73e-20 
C10214 VCC.n6232 VSS 3.7e-20 
C10215 VCC.n6233 VSS 3.5e-20 
C10216 VCC.n6234 VSS 7.41e-20 
C10217 VCC.t88 VSS 6.42e-19 
C10218 VCC.n6235 VSS 3e-20 
C10219 VCC.n6236 VSS 5.97e-20 
C10220 VCC.n6237 VSS 4.13e-19 
C10221 VCC.n6238 VSS 9.53e-20 
C10222 VCC.n6239 VSS 3.5e-20 
C10223 VCC.n6240 VSS 3.5e-20 
C10224 VCC.n6241 VSS 5.35e-20 
C10225 VCC.n6242 VSS 4.32e-20 
C10226 VCC.n6243 VSS 2.68e-20 
C10227 VCC.n6244 VSS 3.7e-20 
C10228 VCC.n6245 VSS 1.65e-20 
C10229 VCC.n6246 VSS 4.53e-20 
C10230 VCC.n6247 VSS 1.2e-19 
C10231 VCC.n6248 VSS 5.2e-19 
C10232 VCC.n6249 VSS 1.2e-19 
C10233 VCC.n6250 VSS 6.38e-20 
C10234 VCC.n6251 VSS 2.47e-20 
C10235 VCC.n6252 VSS 4.53e-20 
C10236 VCC.n6253 VSS 3.5e-20 
C10237 VCC.n6254 VSS 3.5e-20 
C10238 VCC.n6255 VSS 2.68e-20 
C10239 VCC.n6256 VSS 2.68e-20 
C10240 VCC.n6257 VSS 2.47e-20 
C10241 VCC.n6258 VSS 4.53e-20 
C10242 VCC.n6259 VSS 2.68e-20 
C10243 VCC.n6260 VSS 4.32e-20 
C10244 VCC.n6261 VSS 2.68e-20 
C10245 VCC.n6262 VSS 3.91e-20 
C10246 VCC.n6263 VSS 2.88e-20 
C10247 VCC.n6264 VSS 4.73e-20 
C10248 VCC.n6265 VSS 3.7e-20 
C10249 VCC.n6266 VSS 3.7e-20 
C10250 VCC.n6267 VSS 3.5e-20 
C10251 VCC.n6268 VSS 5.76e-20 
C10252 VCC.n6269 VSS 4.73e-20 
C10253 VCC.n6270 VSS 3.09e-20 
C10254 VCC.n6271 VSS 3.5e-20 
C10255 VCC.n6272 VSS 3.5e-20 
C10256 VCC.n6273 VSS 3.5e-20 
C10257 VCC.n6274 VSS 1.18e-19 
C10258 VCC.n6275 VSS 3e-20 
C10259 VCC.n6276 VSS 1.15e-19 
C10260 VCC.n6277 VSS 9.88e-20 
C10261 VCC.n6278 VSS 5.76e-20 
C10262 VCC.n6279 VSS 3.5e-20 
C10263 VCC.n6280 VSS 3.09e-20 
C10264 VCC.n6281 VSS 3.09e-20 
C10265 VCC.n6282 VSS 2.26e-20 
C10266 VCC.n6283 VSS 5.76e-20 
C10267 VCC.n6284 VSS 2.68e-20 
C10268 VCC.n6285 VSS 2.68e-20 
C10269 VCC.n6286 VSS 0.00185f 
C10270 VCC.n6287 VSS 2.72e-19 
C10271 VCC.n6288 VSS 2.26e-20 
C10272 VCC.n6289 VSS 1.87e-19 
C10273 VCC.n6290 VSS 3.5e-20 
C10274 VCC.n6291 VSS 2.68e-20 
C10275 VCC.n6292 VSS 5.97e-20 
C10276 VCC.n6293 VSS 4.73e-20 
C10277 VCC.n6294 VSS 4.73e-20 
C10278 VCC.n6295 VSS 5.15e-20 
C10279 VCC.n6296 VSS 7.41e-20 
C10280 VCC.n6297 VSS 3.7e-20 
C10281 VCC.n6298 VSS 2.26e-20 
C10282 VCC.n6299 VSS 6.38e-20 
C10283 VCC.n6300 VSS 4.73e-20 
C10284 VCC.n6301 VSS 3.29e-20 
C10285 VCC.n6302 VSS 3.5e-20 
C10286 VCC.n6303 VSS 3e-20 
C10287 VCC.t61 VSS 0.005f 
C10288 VCC.t221 VSS 0.00453f 
C10289 VCC.n6304 VSS 0.00228f 
C10290 VCC.n6305 VSS 1.3e-19 
C10291 VCC.t59 VSS 4.05e-19 
C10292 VCC.n6306 VSS 4.05e-19 
C10293 VCC.n6307 VSS 1.15e-19 
C10294 VCC.n6308 VSS 3.36e-19 
C10295 VCC.n6309 VSS 6.17e-21 
C10296 VCC.n6310 VSS 3.12e-19 
C10297 VCC.n6311 VSS 1.65e-20 
C10298 VCC.n6312 VSS 1.54e-19 
C10299 VCC.n6313 VSS 1.54e-19 
C10300 VCC.n6314 VSS 1.65e-20 
C10301 VCC.n6315 VSS 1.03e-20 
C10302 VCC.n6316 VSS 3.5e-20 
C10303 VCC.n6317 VSS 2.26e-20 
C10304 VCC.n6318 VSS 4.73e-20 
C10305 VCC.n6319 VSS 3.5e-20 
C10306 VCC.n6320 VSS 3e-20 
C10307 VCC.n6321 VSS 1.3e-19 
C10308 VCC.n6322 VSS 5.12e-19 
C10309 VCC.n6323 VSS 1.3e-19 
C10310 VCC.n6324 VSS 4.13e-19 
C10311 VCC.n6325 VSS 9.53e-20 
C10312 VCC.n6326 VSS 5.76e-20 
C10313 VCC.n6327 VSS 7.41e-20 
C10314 VCC.n6328 VSS 5.56e-20 
C10315 VCC.t60 VSS 1.55e-19 
C10316 VCC.n6329 VSS 3.91e-20 
C10317 VCC.n6330 VSS 3.91e-20 
C10318 VCC.n6331 VSS 1.85e-20 
C10319 VCC.n6332 VSS 7.55e-19 
C10320 VCC.n6333 VSS 4.94e-20 
C10321 VCC.n6334 VSS 5.15e-20 
C10322 VCC.n6335 VSS 7.2e-20 
C10323 VCC.n6336 VSS 1.38e-19 
C10324 VCC.n6337 VSS 1.17e-19 
C10325 VCC.n6338 VSS 4.32e-20 
C10326 VCC.n6339 VSS 2.88e-20 
C10327 VCC.n6340 VSS 2.68e-20 
C10328 VCC.n6341 VSS 3.5e-20 
C10329 VCC.n6342 VSS 3.5e-20 
C10330 VCC.n6343 VSS 2.88e-20 
C10331 VCC.n6344 VSS 2.68e-20 
C10332 VCC.n6345 VSS 2.68e-20 
C10333 VCC.n6346 VSS 2.68e-20 
C10334 VCC.n6347 VSS 4.12e-20 
C10335 VCC.n6348 VSS 4.12e-20 
C10336 VCC.n6349 VSS 3.91e-20 
C10337 VCC.n6350 VSS 4.53e-20 
C10338 VCC.n6351 VSS 4.53e-20 
C10339 VCC.n6352 VSS 1.05e-19 
C10340 VCC.n6353 VSS 1.05e-19 
C10341 VCC.n6354 VSS 4.32e-20 
C10342 VCC.n6355 VSS 3.7e-20 
C10343 VCC.n6356 VSS 2.68e-20 
C10344 VCC.n6357 VSS 2.68e-20 
C10345 VCC.n6358 VSS 6.79e-20 
C10346 VCC.n6359 VSS 9.26e-20 
C10347 VCC.n6360 VSS 1.83e-19 
C10348 VCC.n6361 VSS 7.95e-19 
C10349 VCC.n6362 VSS 5.2e-19 
C10350 VCC.n6363 VSS 1.3e-19 
C10351 VCC.n6364 VSS 3e-20 
C10352 VCC.n6365 VSS 3.5e-20 
C10353 VCC.n6366 VSS 5.97e-20 
C10354 VCC.n6367 VSS 7.41e-20 
C10355 VCC.n6368 VSS 5.15e-20 
C10356 VCC.n6369 VSS 5.15e-20 
C10357 VCC.n6370 VSS 3.09e-20 
C10358 VCC.n6371 VSS 3.09e-20 
C10359 VCC.n6372 VSS 3.7e-20 
C10360 VCC.n6373 VSS 2.68e-20 
C10361 VCC.n6374 VSS 3.91e-20 
C10362 VCC.n6375 VSS 1.17e-19 
C10363 VCC.n6376 VSS 1.38e-19 
C10364 VCC.n6377 VSS 7e-20 
C10365 VCC.n6378 VSS 4.73e-20 
C10366 VCC.n6379 VSS 3.5e-20 
C10367 VCC.n6380 VSS 3.5e-20 
C10368 VCC.n6381 VSS 3.5e-20 
C10369 VCC.n6382 VSS 4.53e-20 
C10370 VCC.n6383 VSS 1.18e-19 
C10371 VCC.n6384 VSS 5.12e-19 
C10372 VCC.n6385 VSS 1.3e-19 
C10373 VCC.n6386 VSS 1.61e-19 
C10374 VCC.n6387 VSS 9.9e-20 
C10375 VCC.n6388 VSS 0.00243f 
C10376 VCC.n6389 VSS 2.26e-20 
C10377 VCC.n6390 VSS 4.13e-19 
C10378 VCC.n6391 VSS 3.5e-20 
C10379 VCC.n6392 VSS 3.5e-20 
C10380 VCC.n6393 VSS 2.47e-20 
C10381 VCC.n6394 VSS 2.06e-20 
C10382 VCC.n6395 VSS 6.17e-20 
C10383 VCC.n6396 VSS 6.17e-20 
C10384 VCC.n6397 VSS 4.73e-20 
C10385 VCC.n6398 VSS 4.73e-20 
C10386 VCC.n6399 VSS 2.88e-20 
C10387 VCC.n6400 VSS 1.44e-20 
C10388 VCC.n6401 VSS 1.65e-20 
C10389 VCC.n6402 VSS 1.54e-19 
C10390 VCC.n6403 VSS 1.54e-19 
C10391 VCC.n6404 VSS 1.65e-20 
C10392 VCC.n6405 VSS 3.09e-20 
C10393 VCC.t89 VSS 1.55e-19 
C10394 VCC.n6406 VSS 0.00102f 
C10395 VCC.n6407 VSS 2.73e-19 
C10396 VCC.n6408 VSS 0.00136f 
C10397 VCC.n6409 VSS 2.73e-19 
C10398 VCC.n6410 VSS 0.00181f 
C10399 VCC.n6411 VSS 5.76e-20 
C10400 VCC.n6412 VSS 1.54e-19 
C10401 VCC.n6413 VSS 1.65e-20 
C10402 VCC.n6414 VSS 2.88e-20 
C10403 VCC.n6415 VSS 2.47e-20 
C10404 VCC.n6416 VSS 6.17e-20 
C10405 VCC.n6417 VSS 4.73e-20 
C10406 VCC.n6418 VSS 4.73e-20 
C10407 VCC.n6419 VSS 5.15e-20 
C10408 VCC.n6420 VSS 3.5e-20 
C10409 VCC.n6421 VSS 7.41e-20 
C10410 VCC.n6422 VSS 3.7e-20 
C10411 VCC.n6423 VSS 2.26e-20 
C10412 VCC.n6424 VSS 6.17e-20 
C10413 VCC.n6425 VSS 4.73e-20 
C10414 VCC.n6426 VSS 3.5e-20 
C10415 VCC.n6427 VSS 2.88e-20 
C10416 VCC.n6428 VSS 3.4e-19 
C10417 VCC.n6429 VSS 1.15e-19 
C10418 VCC.n6430 VSS 3.98e-19 
C10419 VCC.t15 VSS 4.05e-19 
C10420 VCC.n6431 VSS 1.22e-19 
C10421 VCC.n6432 VSS 1.3e-19 
C10422 VCC.n6433 VSS 3e-20 
C10423 VCC.n6434 VSS 3.5e-20 
C10424 VCC.n6435 VSS 3.5e-20 
C10425 VCC.n6436 VSS 4.73e-20 
C10426 VCC.n6437 VSS 2.47e-20 
C10427 VCC.n6438 VSS 1.23e-20 
C10428 VCC.n6439 VSS 1.65e-20 
C10429 VCC.n6440 VSS 2.47e-20 
C10430 VCC.n6441 VSS 5.76e-20 
C10431 VCC.n6442 VSS 1.38e-19 
C10432 VCC.n6443 VSS 7e-20 
C10433 VCC.n6444 VSS 3.7e-20 
C10434 VCC.n6445 VSS 2.47e-20 
C10435 VCC.n6446 VSS 3.7e-20 
C10436 VCC.n6447 VSS 1.85e-20 
C10437 VCC.n6448 VSS 3.09e-20 
C10438 VCC.n6449 VSS 5.35e-20 
C10439 VCC.n6450 VSS 4.73e-20 
C10440 VCC.n6451 VSS 5.35e-20 
C10441 VCC.n6452 VSS 7.41e-20 
C10442 VCC.n6453 VSS 5.76e-20 
C10443 VCC.n6454 VSS 9.53e-20 
C10444 VCC.n6455 VSS 4.13e-19 
C10445 VCC.n6456 VSS 1.3e-19 
C10446 VCC.n6457 VSS 5.2e-19 
C10447 VCC.n6458 VSS 1.2e-19 
C10448 VCC.n6459 VSS 4.73e-20 
C10449 VCC.n6460 VSS 2.68e-20 
C10450 VCC.n6461 VSS 3.5e-20 
C10451 VCC.n6462 VSS 3.5e-20 
C10452 VCC.n6463 VSS 2.68e-20 
C10453 VCC.n6464 VSS 2.68e-20 
C10454 VCC.n6465 VSS 4.32e-20 
C10455 VCC.n6466 VSS 4.32e-20 
C10456 VCC.n6467 VSS 4.32e-20 
C10457 VCC.n6468 VSS 2.88e-20 
C10458 VCC.n6469 VSS 3.5e-20 
C10459 VCC.n6470 VSS 2.68e-20 
C10460 VCC.n6471 VSS 7.82e-20 
C10461 VCC.n6472 VSS 4.73e-20 
C10462 VCC.n6473 VSS 4.73e-20 
C10463 VCC.n6474 VSS 1.05e-19 
C10464 VCC.n6475 VSS 1.05e-19 
C10465 VCC.n6476 VSS 4.53e-20 
C10466 VCC.n6477 VSS 2.68e-20 
C10467 VCC.n6478 VSS 2.68e-20 
C10468 VCC.n6479 VSS 6.59e-20 
C10469 VCC.n6480 VSS 9.26e-20 
C10470 VCC.n6481 VSS 6.59e-20 
C10471 VCC.n6482 VSS 2.47e-20 
C10472 VCC.n6483 VSS 2.47e-20 
C10473 VCC.n6484 VSS 2.88e-20 
C10474 VCC.n6485 VSS 3.5e-20 
C10475 VCC.n6486 VSS 3.5e-20 
C10476 VCC.n6487 VSS 4.53e-20 
C10477 VCC.n6488 VSS 1.2e-19 
C10478 VCC.n6489 VSS 5.2e-19 
C10479 VCC.n6490 VSS 1.3e-19 
C10480 VCC.n6491 VSS 4.13e-19 
C10481 VCC.n6492 VSS 9.53e-20 
C10482 VCC.n6493 VSS 5.97e-20 
C10483 VCC.n6494 VSS 7.41e-20 
C10484 VCC.n6495 VSS 5.35e-20 
C10485 VCC.n6496 VSS 5.15e-20 
C10486 VCC.n6497 VSS 3.09e-20 
C10487 VCC.n6498 VSS 3.09e-20 
C10488 VCC.n6499 VSS 3.91e-20 
C10489 VCC.n6500 VSS 2.47e-20 
C10490 VCC.n6501 VSS 3.7e-20 
C10491 VCC.n6502 VSS 1.17e-19 
C10492 VCC.n6503 VSS 1.38e-19 
C10493 VCC.n6504 VSS 7.2e-20 
C10494 VCC.n6505 VSS 4.73e-20 
C10495 VCC.n6506 VSS 3.5e-20 
C10496 VCC.n6507 VSS 3.5e-20 
C10497 VCC.n6508 VSS 4.53e-20 
C10498 VCC.n6509 VSS 5.97e-20 
C10499 VCC.n6510 VSS 3.5e-20 
C10500 VCC.n6511 VSS 3e-20 
C10501 VCC.n6512 VSS 1.3e-19 
C10502 VCC.n6513 VSS 1.53e-19 
C10503 VCC.t165 VSS 4.05e-19 
C10504 VCC.n6514 VSS 2.06e-19 
C10505 VCC.n6515 VSS 1.35e-19 
C10506 VCC.n6516 VSS 9.67e-20 
C10507 VCC.n6517 VSS 3.35e-20 
C10508 VCC.n6518 VSS 3.5e-20 
C10509 VCC.n6519 VSS 2.36e-19 
C10510 VCC.n6520 VSS 0.0023f 
C10511 VCC.t168 VSS 0.0031f 
C10512 VCC.t84 VSS 0.00366f 
C10513 VCC.t167 VSS 0.00365f 
C10514 VCC.t87 VSS 0.00386f 
C10515 VCC.n6521 VSS 0.00569f 
C10516 VCC.n6522 VSS 1.3e-19 
C10517 VCC.n6523 VSS 3.67e-19 
C10518 VCC.n6524 VSS 1.15e-19 
C10519 VCC.n6525 VSS 3.38e-19 
C10520 VCC.n6526 VSS 3.5e-20 
C10521 VCC.n6527 VSS 3.5e-20 
C10522 VCC.n6528 VSS 2.68e-20 
C10523 VCC.n6529 VSS 2.06e-20 
C10524 VCC.n6530 VSS 6.38e-20 
C10525 VCC.n6531 VSS 5.97e-20 
C10526 VCC.n6532 VSS 4.73e-20 
C10527 VCC.n6533 VSS 4.73e-20 
C10528 VCC.n6534 VSS 3.09e-20 
C10529 VCC.n6535 VSS 1.23e-20 
C10530 VCC.n6536 VSS 1.65e-20 
C10531 VCC.n6537 VSS 1.54e-19 
C10532 VCC.n6538 VSS 1.54e-19 
C10533 VCC.n6539 VSS 1.65e-20 
C10534 VCC.n6540 VSS 3.29e-20 
C10535 VCC.t166 VSS 1.67e-19 
C10536 VCC.n6541 VSS 0.00101f 
C10537 VCC.n6542 VSS 2.71e-19 
C10538 VCC.n6543 VSS 7.46e-19 
C10539 VCC.n6544 VSS 0.00333f 
C10540 VCC.n6545 VSS 2.46e-19 
C10541 VCC.n6546 VSS 3.02e-19 
C10542 VCC.n6547 VSS 3.7e-20 
C10543 VCC.n6548 VSS 5.15e-20 
C10544 VCC.n6549 VSS 6.38e-20 
C10545 VCC.n6550 VSS 4.73e-20 
C10546 VCC.n6551 VSS 4.73e-20 
C10547 VCC.n6552 VSS 2.68e-20 
C10548 VCC.n6553 VSS 3.29e-20 
C10549 VCC.n6554 VSS 1.65e-20 
C10550 VCC.n6555 VSS 1.54e-19 
C10551 VCC.n6556 VSS 1.54e-19 
C10552 VCC.n6557 VSS 5.56e-20 
C10553 VCC.n6558 VSS 2.88e-20 
C10554 VCC.n6559 VSS 1.65e-20 
C10555 VCC.n6560 VSS 3.09e-20 
C10556 VCC.n6561 VSS 4.73e-20 
C10557 VCC.n6562 VSS 4.73e-20 
C10558 VCC.n6563 VSS 4.32e-20 
C10559 VCC.n6564 VSS 1.17e-19 
C10560 VCC.n6565 VSS 3.33e-19 
C10561 VCC.n6566 VSS 1.35e-19 
C10562 VCC.n6567 VSS 4.37e-19 
C10563 VCC.n6568 VSS 5.24e-19 
C10564 VCC.n6569 VSS 1.36e-19 
C10565 VCC.n6570 VSS 1.01e-19 
C10566 VCC.n6571 VSS 1.05e-19 
C10567 VCC.n6572 VSS 2.06e-20 
C10568 VCC.n6573 VSS 2.26e-20 
C10569 VCC.n6574 VSS 3.7e-20 
C10570 VCC.n6575 VSS 5.15e-20 
C10571 VCC.n6576 VSS 1.38e-19 
C10572 VCC.n6577 VSS 3.91e-20 
C10573 VCC.n6578 VSS 2.88e-20 
C10574 VCC.n6579 VSS 4.32e-20 
C10575 VCC.n6580 VSS 1.17e-19 
C10576 VCC.n6581 VSS 3.7e-20 
C10577 VCC.n6582 VSS 3.91e-20 
C10578 VCC.n6583 VSS 3.5e-20 
C10579 VCC.n6584 VSS 1.65e-20 
C10580 VCC.n6585 VSS 8.23e-21 
C10581 VCC.n6586 VSS 3.5e-20 
C10582 VCC.n6587 VSS 3.5e-20 
C10583 VCC.n6588 VSS 1.4e-19 
C10584 VCC.n6589 VSS 5.4e-19 
C10585 VCC.n6590 VSS 8.42e-19 
C10586 VCC.n6591 VSS 5.4e-19 
C10587 VCC.n6592 VSS 1.4e-19 
C10588 VCC.n6593 VSS 1.4e-19 
C10589 VCC.n6594 VSS 2.18e-19 
C10590 VCC.n6595 VSS 7.82e-20 
C10591 VCC.n6596 VSS 4.32e-20 
C10592 VCC.n6597 VSS 4.32e-20 
C10593 VCC.n6598 VSS 1.05e-19 
C10594 VCC.n6599 VSS 1.05e-19 
C10595 VCC.n6600 VSS 4.32e-20 
C10596 VCC.n6601 VSS 3.7e-20 
C10597 VCC.n6602 VSS 2.68e-20 
C10598 VCC.n6603 VSS 5.76e-20 
C10599 VCC.n6604 VSS 6.38e-20 
C10600 VCC.n6605 VSS 3.5e-20 
C10601 VCC.n6606 VSS 3.5e-20 
C10602 VCC.n6607 VSS 1.17e-19 
C10603 VCC.n6608 VSS 1.38e-19 
C10604 VCC.n6609 VSS 5.15e-20 
C10605 VCC.n6610 VSS 1.05e-19 
C10606 VCC.n6611 VSS 2.26e-20 
C10607 VCC.n6612 VSS 5.76e-20 
C10608 VCC.n6613 VSS 3.7e-20 
C10609 VCC.n6614 VSS 3.7e-20 
C10610 VCC.n6615 VSS 3.09e-20 
C10611 VCC.n6616 VSS 1.85e-20 
C10612 VCC.n6617 VSS 1.65e-20 
C10613 VCC.n6618 VSS 8.23e-21 
C10614 VCC.n6619 VSS 1.13e-19 
C10615 VCC.n6620 VSS 3.33e-19 
C10616 VCC.t237 VSS 4.21e-19 
C10617 VCC.n6621 VSS 2.06e-19 
C10618 VCC.n6622 VSS 1.35e-19 
C10619 VCC.n6623 VSS 3.5e-20 
C10620 VCC.n6624 VSS 3.5e-20 
C10621 VCC.n6625 VSS 3.5e-20 
C10622 VCC.n6626 VSS 1.03e-20 
C10623 VCC.n6627 VSS 2.68e-20 
C10624 VCC.n6628 VSS 3.09e-20 
C10625 VCC.n6629 VSS 2.68e-20 
C10626 VCC.n6630 VSS 1.65e-20 
C10627 VCC.n6631 VSS 1.54e-19 
C10628 VCC.n6632 VSS 1.54e-19 
C10629 VCC.n6633 VSS 1.65e-20 
C10630 VCC.t238 VSS 1.56e-19 
C10631 VCC.n6634 VSS 7.62e-19 
C10632 VCC.n6635 VSS 1.23e-20 
C10633 VCC.n6636 VSS 2.47e-20 
C10634 VCC.n6637 VSS 4.73e-20 
C10635 VCC.n6638 VSS 6.59e-20 
C10636 VCC.n6639 VSS 5.15e-20 
C10637 VCC.n6640 VSS 2.47e-20 
C10638 VCC.n6641 VSS 7.41e-20 
C10639 VCC.n6642 VSS 9.47e-20 
C10640 VCC.n6643 VSS 1.32e-19 
C10641 VCC.n6644 VSS 7.71e-19 
C10642 VCC.n6645 VSS 9.83e-19 
C10643 VCC.n6646 VSS 2.36e-19 
C10644 VCC.n6647 VSS 3.21e-19 
C10645 VCC.n6648 VSS 2.61e-19 
C10646 VCC.n6649 VSS 0.00189f 
C10647 VCC.n6650 VSS 5.76e-20 
C10648 VCC.n6651 VSS 2.88e-20 
C10649 VCC.n6652 VSS 3.5e-20 
C10650 VCC.n6653 VSS 9.83e-19 
C10651 VCC.n6654 VSS 9.47e-20 
C10652 VCC.n6655 VSS 1.17e-19 
C10653 VCC.n6656 VSS 2.06e-19 
C10654 VCC.n6657 VSS 1.36e-19 
C10655 VCC.n6658 VSS 1.01e-19 
C10656 VCC.n6659 VSS 3.5e-20 
C10657 VCC.n6660 VSS 3.09e-20 
C10658 VCC.n6661 VSS 3.29e-20 
C10659 VCC.n6662 VSS 3.29e-20 
C10660 VCC.n6663 VSS 4.73e-20 
C10661 VCC.n6664 VSS 1.44e-20 
C10662 VCC.n6665 VSS 3.5e-20 
C10663 VCC.n6666 VSS 7.41e-20 
C10664 VCC.n6667 VSS 2.47e-20 
C10665 VCC.t86 VSS 1.56e-19 
C10666 VCC.n6668 VSS 5.76e-20 
C10667 VCC.n6669 VSS 2.06e-20 
C10668 VCC.n6670 VSS 5.76e-20 
C10669 VCC.n6671 VSS 3.7e-20 
C10670 VCC.n6672 VSS 4.32e-20 
C10671 VCC.n6673 VSS 2.68e-20 
C10672 VCC.n6674 VSS 3.91e-20 
C10673 VCC.n6675 VSS 6.38e-20 
C10674 VCC.n6676 VSS 1.85e-20 
C10675 VCC.n6677 VSS 3.5e-20 
C10676 VCC.n6678 VSS 3.09e-20 
C10677 VCC.n6679 VSS 3.7e-20 
C10678 VCC.n6680 VSS 3.09e-20 
C10679 VCC.n6681 VSS 2.26e-20 
C10680 VCC.n6682 VSS 1.05e-19 
C10681 VCC.n6683 VSS 3.5e-20 
C10682 VCC.n6684 VSS 3.5e-20 
C10683 VCC.n6685 VSS 8.42e-19 
C10684 VCC.n6686 VSS 2.18e-19 
C10685 VCC.n6687 VSS 1.4e-19 
C10686 VCC.n6688 VSS 4.32e-20 
C10687 VCC.n6689 VSS 7.82e-20 
C10688 VCC.n6690 VSS 5.76e-20 
C10689 VCC.n6691 VSS 2.68e-20 
C10690 VCC.n6692 VSS 4.32e-20 
C10691 VCC.n6693 VSS 3.91e-20 
C10692 VCC.n6694 VSS 3.7e-20 
C10693 VCC.n6695 VSS 3.7e-20 
C10694 VCC.n6696 VSS 5.76e-20 
C10695 VCC.n6697 VSS 4.73e-20 
C10696 VCC.n6698 VSS 3.5e-20 
C10697 VCC.t109 VSS 1.56e-19 
C10698 VCC.n6699 VSS 7.97e-19 
C10699 VCC.n6700 VSS 3.09e-20 
C10700 VCC.n6701 VSS 1.01e-19 
C10701 VCC.n6702 VSS 3.5e-20 
C10702 VCC.n6703 VSS 1.36e-19 
C10703 VCC.n6704 VSS 3.5e-20 
C10704 VCC.n6705 VSS 3.33e-19 
C10705 VCC.n6706 VSS 1.17e-19 
C10706 VCC.n6707 VSS 1.09e-19 
C10707 VCC.n6708 VSS 3.5e-20 
C10708 VCC.n6709 VSS 4.73e-20 
C10709 VCC.n6710 VSS 5.56e-20 
C10710 VCC.n6711 VSS 2.88e-20 
C10711 VCC.n6712 VSS 2.26e-20 
C10712 VCC.n6713 VSS 5.76e-20 
C10713 VCC.n6714 VSS 2.68e-20 
C10714 VCC.n6715 VSS 2.68e-20 
C10715 VCC.n6716 VSS 1.9e-19 
C10716 VCC.n6717 VSS 5.76e-20 
C10717 VCC.n6718 VSS 2.68e-20 
C10718 VCC.n6719 VSS 2.68e-20 
C10719 VCC.n6720 VSS 2.68e-20 
C10720 VCC.n6721 VSS 5.76e-20 
C10721 VCC.n6722 VSS 2.26e-20 
C10722 VCC.n6723 VSS 3.09e-20 
C10723 VCC.n6724 VSS 2.26e-20 
C10724 VCC.n6725 VSS 5.15e-20 
C10725 VCC.n6726 VSS 4.73e-20 
C10726 VCC.n6727 VSS 3.7e-20 
C10727 VCC.n6728 VSS 3.5e-20 
C10728 VCC.n6729 VSS 7.41e-20 
C10729 VCC.n6730 VSS 1.91e-19 
C10730 VCC.n6731 VSS 9.88e-20 
C10731 VCC.n6732 VSS 3e-20 
C10732 VCC.n6733 VSS 5.12e-19 
C10733 VCC.n6734 VSS 1.18e-19 
C10734 VCC.n6735 VSS 3.5e-20 
C10735 VCC.n6736 VSS 3.5e-20 
C10736 VCC.n6737 VSS 5.15e-20 
C10737 VCC.n6738 VSS 4.32e-20 
C10738 VCC.n6739 VSS 2.68e-20 
C10739 VCC.n6740 VSS 3.91e-20 
C10740 VCC.n6741 VSS 1.44e-20 
C10741 VCC.n6742 VSS 3.5e-20 
C10742 VCC.n6743 VSS 3e-20 
C10743 VCC.n6744 VSS 7.95e-19 
C10744 VCC.n6745 VSS 1.83e-19 
C10745 VCC.n6746 VSS 2.88e-20 
C10746 VCC.n6747 VSS 2.68e-20 
C10747 VCC.n6748 VSS 2.68e-20 
C10748 VCC.n6749 VSS 2.68e-20 
C10749 VCC.n6750 VSS 4.53e-20 
C10750 VCC.n6751 VSS 3.7e-20 
C10751 VCC.n6752 VSS 7.82e-20 
C10752 VCC.n6753 VSS 1.17e-19 
C10753 VCC.n6754 VSS 3.91e-20 
C10754 VCC.n6755 VSS 1.65e-20 
C10755 VCC.n6756 VSS 2.68e-20 
C10756 VCC.n6757 VSS 3.5e-20 
C10757 VCC.n6758 VSS 3e-20 
C10758 VCC.n6759 VSS 5.12e-19 
C10759 VCC.n6760 VSS 1.18e-19 
C10760 VCC.n6761 VSS 3.5e-20 
C10761 VCC.n6762 VSS 3.5e-20 
C10762 VCC.t157 VSS 1.55e-19 
C10763 VCC.n6763 VSS 7.57e-19 
C10764 VCC.n6764 VSS 4.73e-20 
C10765 VCC.n6765 VSS 1.54e-19 
C10766 VCC.n6766 VSS 2.88e-20 
C10767 VCC.n6767 VSS 2.88e-20 
C10768 VCC.n6768 VSS 3.5e-20 
C10769 VCC.n6769 VSS 5.76e-20 
C10770 VCC.n6770 VSS 9.88e-20 
C10771 VCC.n6771 VSS 1.3e-19 
C10772 VCC.n6772 VSS 3e-20 
C10773 VCC.t155 VSS 0.005f 
C10774 VCC.t62 VSS 0.00453f 
C10775 VCC.n6773 VSS 0.00229f 
C10776 VCC.n6774 VSS 1.91e-19 
C10777 VCC.n6775 VSS 3.5e-20 
C10778 VCC.n6776 VSS 3.14e-19 
C10779 VCC.n6777 VSS 3.5e-20 
C10780 VCC.n6778 VSS 2.47e-20 
C10781 VCC.n6779 VSS 5.76e-20 
C10782 VCC.n6780 VSS 2.47e-20 
C10783 VCC.n6781 VSS 8.23e-21 
C10784 VCC.n6782 VSS 2.88e-20 
C10785 VCC.n6783 VSS 5.76e-20 
C10786 VCC.n6784 VSS 2.47e-20 
C10787 VCC.n6785 VSS 2.88e-20 
C10788 VCC.n6786 VSS 2.47e-20 
C10789 VCC.n6787 VSS 5.15e-20 
C10790 VCC.n6788 VSS 4.73e-20 
C10791 VCC.n6789 VSS 3.7e-20 
C10792 VCC.n6790 VSS 3.5e-20 
C10793 VCC.n6791 VSS 7.41e-20 
C10794 VCC.t82 VSS 6.42e-19 
C10795 VCC.n6792 VSS 3e-20 
C10796 VCC.n6793 VSS 5.97e-20 
C10797 VCC.n6794 VSS 4.13e-19 
C10798 VCC.n6795 VSS 9.53e-20 
C10799 VCC.n6796 VSS 3.5e-20 
C10800 VCC.n6797 VSS 3.5e-20 
C10801 VCC.n6798 VSS 5.35e-20 
C10802 VCC.n6799 VSS 4.32e-20 
C10803 VCC.n6800 VSS 2.68e-20 
C10804 VCC.n6801 VSS 3.7e-20 
C10805 VCC.n6802 VSS 1.65e-20 
C10806 VCC.n6803 VSS 4.53e-20 
C10807 VCC.n6804 VSS 1.2e-19 
C10808 VCC.n6805 VSS 5.2e-19 
C10809 VCC.n6806 VSS 1.2e-19 
C10810 VCC.n6807 VSS 6.38e-20 
C10811 VCC.n6808 VSS 2.47e-20 
C10812 VCC.n6809 VSS 4.53e-20 
C10813 VCC.n6810 VSS 3.5e-20 
C10814 VCC.n6811 VSS 3.5e-20 
C10815 VCC.n6812 VSS 2.68e-20 
C10816 VCC.n6813 VSS 2.68e-20 
C10817 VCC.n6814 VSS 2.47e-20 
C10818 VCC.n6815 VSS 4.53e-20 
C10819 VCC.n6816 VSS 2.68e-20 
C10820 VCC.n6817 VSS 4.32e-20 
C10821 VCC.n6818 VSS 2.68e-20 
C10822 VCC.n6819 VSS 3.91e-20 
C10823 VCC.n6820 VSS 2.88e-20 
C10824 VCC.n6821 VSS 4.73e-20 
C10825 VCC.n6822 VSS 3.7e-20 
C10826 VCC.n6823 VSS 3.7e-20 
C10827 VCC.n6824 VSS 3.5e-20 
C10828 VCC.n6825 VSS 5.76e-20 
C10829 VCC.n6826 VSS 4.73e-20 
C10830 VCC.n6827 VSS 3.09e-20 
C10831 VCC.n6828 VSS 3.5e-20 
C10832 VCC.n6829 VSS 3.5e-20 
C10833 VCC.n6830 VSS 3.5e-20 
C10834 VCC.n6831 VSS 1.18e-19 
C10835 VCC.n6832 VSS 3e-20 
C10836 VCC.n6833 VSS 1.15e-19 
C10837 VCC.n6834 VSS 9.88e-20 
C10838 VCC.n6835 VSS 5.76e-20 
C10839 VCC.n6836 VSS 3.5e-20 
C10840 VCC.n6837 VSS 3.09e-20 
C10841 VCC.n6838 VSS 3.09e-20 
C10842 VCC.n6839 VSS 2.26e-20 
C10843 VCC.n6840 VSS 5.76e-20 
C10844 VCC.n6841 VSS 2.68e-20 
C10845 VCC.n6842 VSS 2.68e-20 
C10846 VCC.n6843 VSS 0.00185f 
C10847 VCC.n6844 VSS 2.72e-19 
C10848 VCC.n6845 VSS 2.26e-20 
C10849 VCC.n6846 VSS 1.87e-19 
C10850 VCC.n6847 VSS 3.5e-20 
C10851 VCC.n6848 VSS 2.68e-20 
C10852 VCC.n6849 VSS 5.97e-20 
C10853 VCC.n6850 VSS 4.73e-20 
C10854 VCC.n6851 VSS 4.73e-20 
C10855 VCC.n6852 VSS 5.15e-20 
C10856 VCC.n6853 VSS 7.41e-20 
C10857 VCC.n6854 VSS 3.7e-20 
C10858 VCC.n6855 VSS 2.26e-20 
C10859 VCC.n6856 VSS 6.38e-20 
C10860 VCC.n6857 VSS 4.73e-20 
C10861 VCC.n6858 VSS 3.29e-20 
C10862 VCC.n6859 VSS 3.5e-20 
C10863 VCC.n6860 VSS 3e-20 
C10864 VCC.t43 VSS 0.005f 
C10865 VCC.t205 VSS 0.00453f 
C10866 VCC.n6861 VSS 0.00228f 
C10867 VCC.n6862 VSS 1.3e-19 
C10868 VCC.t41 VSS 4.05e-19 
C10869 VCC.n6863 VSS 4.05e-19 
C10870 VCC.n6864 VSS 1.15e-19 
C10871 VCC.n6865 VSS 3.36e-19 
C10872 VCC.n6866 VSS 6.17e-21 
C10873 VCC.n6867 VSS 3.12e-19 
C10874 VCC.n6868 VSS 1.65e-20 
C10875 VCC.n6869 VSS 1.54e-19 
C10876 VCC.n6870 VSS 1.54e-19 
C10877 VCC.n6871 VSS 1.65e-20 
C10878 VCC.n6872 VSS 1.03e-20 
C10879 VCC.n6873 VSS 3.5e-20 
C10880 VCC.n6874 VSS 2.26e-20 
C10881 VCC.n6875 VSS 4.73e-20 
C10882 VCC.n6876 VSS 3.5e-20 
C10883 VCC.n6877 VSS 3e-20 
C10884 VCC.n6878 VSS 1.3e-19 
C10885 VCC.n6879 VSS 5.12e-19 
C10886 VCC.n6880 VSS 1.3e-19 
C10887 VCC.n6881 VSS 4.13e-19 
C10888 VCC.n6882 VSS 9.53e-20 
C10889 VCC.n6883 VSS 5.76e-20 
C10890 VCC.n6884 VSS 7.41e-20 
C10891 VCC.n6885 VSS 5.56e-20 
C10892 VCC.t42 VSS 1.55e-19 
C10893 VCC.n6886 VSS 3.91e-20 
C10894 VCC.n6887 VSS 3.91e-20 
C10895 VCC.n6888 VSS 1.85e-20 
C10896 VCC.n6889 VSS 7.55e-19 
C10897 VCC.n6890 VSS 4.94e-20 
C10898 VCC.n6891 VSS 5.15e-20 
C10899 VCC.n6892 VSS 7.2e-20 
C10900 VCC.n6893 VSS 1.38e-19 
C10901 VCC.n6894 VSS 1.17e-19 
C10902 VCC.n6895 VSS 4.32e-20 
C10903 VCC.n6896 VSS 2.88e-20 
C10904 VCC.n6897 VSS 2.68e-20 
C10905 VCC.n6898 VSS 3.5e-20 
C10906 VCC.n6899 VSS 3.5e-20 
C10907 VCC.n6900 VSS 2.88e-20 
C10908 VCC.n6901 VSS 2.68e-20 
C10909 VCC.n6902 VSS 2.68e-20 
C10910 VCC.n6903 VSS 2.68e-20 
C10911 VCC.n6904 VSS 4.12e-20 
C10912 VCC.n6905 VSS 4.12e-20 
C10913 VCC.n6906 VSS 3.91e-20 
C10914 VCC.n6907 VSS 4.53e-20 
C10915 VCC.n6908 VSS 4.53e-20 
C10916 VCC.n6909 VSS 1.05e-19 
C10917 VCC.n6910 VSS 1.05e-19 
C10918 VCC.n6911 VSS 4.32e-20 
C10919 VCC.n6912 VSS 3.7e-20 
C10920 VCC.n6913 VSS 2.68e-20 
C10921 VCC.n6914 VSS 2.68e-20 
C10922 VCC.n6915 VSS 6.79e-20 
C10923 VCC.n6916 VSS 9.26e-20 
C10924 VCC.n6917 VSS 1.83e-19 
C10925 VCC.n6918 VSS 7.95e-19 
C10926 VCC.n6919 VSS 5.2e-19 
C10927 VCC.n6920 VSS 1.3e-19 
C10928 VCC.n6921 VSS 3e-20 
C10929 VCC.n6922 VSS 3.5e-20 
C10930 VCC.n6923 VSS 5.97e-20 
C10931 VCC.n6924 VSS 7.41e-20 
C10932 VCC.n6925 VSS 5.15e-20 
C10933 VCC.n6926 VSS 5.15e-20 
C10934 VCC.n6927 VSS 3.09e-20 
C10935 VCC.n6928 VSS 3.09e-20 
C10936 VCC.n6929 VSS 3.7e-20 
C10937 VCC.n6930 VSS 2.68e-20 
C10938 VCC.n6931 VSS 3.91e-20 
C10939 VCC.n6932 VSS 1.17e-19 
C10940 VCC.n6933 VSS 1.38e-19 
C10941 VCC.n6934 VSS 7e-20 
C10942 VCC.n6935 VSS 4.73e-20 
C10943 VCC.n6936 VSS 3.5e-20 
C10944 VCC.n6937 VSS 3.5e-20 
C10945 VCC.n6938 VSS 3.5e-20 
C10946 VCC.n6939 VSS 4.53e-20 
C10947 VCC.n6940 VSS 1.18e-19 
C10948 VCC.n6941 VSS 5.12e-19 
C10949 VCC.n6942 VSS 1.3e-19 
C10950 VCC.n6943 VSS 1.61e-19 
C10951 VCC.n6944 VSS 9.9e-20 
C10952 VCC.n6945 VSS 0.00243f 
C10953 VCC.n6946 VSS 2.26e-20 
C10954 VCC.n6947 VSS 4.13e-19 
C10955 VCC.n6948 VSS 3.5e-20 
C10956 VCC.n6949 VSS 3.5e-20 
C10957 VCC.n6950 VSS 2.47e-20 
C10958 VCC.n6951 VSS 2.06e-20 
C10959 VCC.n6952 VSS 6.17e-20 
C10960 VCC.n6953 VSS 6.17e-20 
C10961 VCC.n6954 VSS 4.73e-20 
C10962 VCC.n6955 VSS 4.73e-20 
C10963 VCC.n6956 VSS 2.88e-20 
C10964 VCC.n6957 VSS 1.44e-20 
C10965 VCC.n6958 VSS 1.65e-20 
C10966 VCC.n6959 VSS 1.54e-19 
C10967 VCC.n6960 VSS 1.54e-19 
C10968 VCC.n6961 VSS 1.65e-20 
C10969 VCC.n6962 VSS 3.09e-20 
C10970 VCC.t83 VSS 1.55e-19 
C10971 VCC.n6963 VSS 0.00102f 
C10972 VCC.n6964 VSS 2.73e-19 
C10973 VCC.n6965 VSS 0.00136f 
C10974 VCC.n6966 VSS 2.73e-19 
C10975 VCC.n6967 VSS 0.00181f 
C10976 VCC.n6968 VSS 5.76e-20 
C10977 VCC.n6969 VSS 1.54e-19 
C10978 VCC.n6970 VSS 1.65e-20 
C10979 VCC.n6971 VSS 6.17e-20 
C10980 VCC.n6972 VSS 2.47e-20 
C10981 VCC.n6973 VSS 4.73e-20 
C10982 VCC.n6974 VSS 4.73e-20 
C10983 VCC.n6975 VSS 5.15e-20 
C10984 VCC.n6976 VSS 3.5e-20 
C10985 VCC.n6977 VSS 7.41e-20 
C10986 VCC.n6978 VSS 3.7e-20 
C10987 VCC.n6979 VSS 2.26e-20 
C10988 VCC.n6980 VSS 6.17e-20 
C10989 VCC.n6981 VSS 4.73e-20 
C10990 VCC.n6982 VSS 2.88e-20 
C10991 VCC.n6983 VSS 2.88e-20 
C10992 VCC.n6984 VSS 3.4e-19 
C10993 VCC.n6985 VSS 1.15e-19 
C10994 VCC.n6986 VSS 3.98e-19 
C10995 VCC.t156 VSS 4.05e-19 
C10996 VCC.n6987 VSS 1.22e-19 
C10997 VCC.n6988 VSS 1.3e-19 
C10998 VCC.n6989 VSS 3e-20 
C10999 VCC.n6990 VSS 3.5e-20 
C11000 VCC.n6991 VSS 3.5e-20 
C11001 VCC.n6992 VSS 4.73e-20 
C11002 VCC.n6993 VSS 2.47e-20 
C11003 VCC.n6994 VSS 1.23e-20 
C11004 VCC.n6995 VSS 1.65e-20 
C11005 VCC.n6996 VSS 2.47e-20 
C11006 VCC.n6997 VSS 5.76e-20 
C11007 VCC.n6998 VSS 1.38e-19 
C11008 VCC.n6999 VSS 7e-20 
C11009 VCC.n7000 VSS 3.7e-20 
C11010 VCC.n7001 VSS 2.47e-20 
C11011 VCC.n7002 VSS 3.7e-20 
C11012 VCC.n7003 VSS 1.85e-20 
C11013 VCC.n7004 VSS 3.09e-20 
C11014 VCC.n7005 VSS 5.35e-20 
C11015 VCC.n7006 VSS 4.73e-20 
C11016 VCC.n7007 VSS 5.35e-20 
C11017 VCC.n7008 VSS 7.41e-20 
C11018 VCC.n7009 VSS 5.76e-20 
C11019 VCC.n7010 VSS 9.53e-20 
C11020 VCC.n7011 VSS 4.13e-19 
C11021 VCC.n7012 VSS 1.3e-19 
C11022 VCC.n7013 VSS 5.2e-19 
C11023 VCC.n7014 VSS 1.2e-19 
C11024 VCC.n7015 VSS 4.73e-20 
C11025 VCC.n7016 VSS 2.68e-20 
C11026 VCC.n7017 VSS 3.5e-20 
C11027 VCC.n7018 VSS 3.5e-20 
C11028 VCC.n7019 VSS 2.68e-20 
C11029 VCC.n7020 VSS 2.68e-20 
C11030 VCC.n7021 VSS 4.32e-20 
C11031 VCC.n7022 VSS 4.32e-20 
C11032 VCC.n7023 VSS 4.32e-20 
C11033 VCC.n7024 VSS 2.88e-20 
C11034 VCC.n7025 VSS 3.5e-20 
C11035 VCC.n7026 VSS 2.68e-20 
C11036 VCC.n7027 VSS 7.82e-20 
C11037 VCC.n7028 VSS 4.73e-20 
C11038 VCC.n7029 VSS 4.73e-20 
C11039 VCC.n7030 VSS 1.05e-19 
C11040 VCC.n7031 VSS 1.05e-19 
C11041 VCC.n7032 VSS 4.53e-20 
C11042 VCC.n7033 VSS 2.68e-20 
C11043 VCC.n7034 VSS 2.68e-20 
C11044 VCC.n7035 VSS 6.59e-20 
C11045 VCC.n7036 VSS 9.26e-20 
C11046 VCC.n7037 VSS 6.59e-20 
C11047 VCC.n7038 VSS 2.47e-20 
C11048 VCC.n7039 VSS 2.47e-20 
C11049 VCC.n7040 VSS 2.88e-20 
C11050 VCC.n7041 VSS 3.5e-20 
C11051 VCC.n7042 VSS 3.5e-20 
C11052 VCC.n7043 VSS 4.53e-20 
C11053 VCC.n7044 VSS 1.2e-19 
C11054 VCC.n7045 VSS 5.2e-19 
C11055 VCC.n7046 VSS 1.3e-19 
C11056 VCC.n7047 VSS 4.13e-19 
C11057 VCC.n7048 VSS 9.53e-20 
C11058 VCC.n7049 VSS 5.97e-20 
C11059 VCC.n7050 VSS 7.41e-20 
C11060 VCC.n7051 VSS 5.35e-20 
C11061 VCC.n7052 VSS 5.15e-20 
C11062 VCC.n7053 VSS 3.09e-20 
C11063 VCC.n7054 VSS 3.09e-20 
C11064 VCC.n7055 VSS 3.91e-20 
C11065 VCC.n7056 VSS 2.47e-20 
C11066 VCC.n7057 VSS 3.7e-20 
C11067 VCC.n7058 VSS 1.17e-19 
C11068 VCC.n7059 VSS 1.38e-19 
C11069 VCC.n7060 VSS 7.2e-20 
C11070 VCC.n7061 VSS 4.73e-20 
C11071 VCC.n7062 VSS 3.5e-20 
C11072 VCC.n7063 VSS 3.5e-20 
C11073 VCC.n7064 VSS 4.53e-20 
C11074 VCC.n7065 VSS 5.97e-20 
C11075 VCC.n7066 VSS 3.5e-20 
C11076 VCC.n7067 VSS 3e-20 
C11077 VCC.n7068 VSS 1.3e-19 
C11078 VCC.n7069 VSS 1.53e-19 
C11079 VCC.t130 VSS 4.05e-19 
C11080 VCC.n7070 VSS 1.35e-19 
C11081 VCC.t108 VSS 4.21e-19 
C11082 VCC.n7071 VSS 2.06e-19 
C11083 VCC.n7072 VSS 1.32e-19 
C11084 VCC.n7073 VSS 9.67e-20 
C11085 VCC.n7074 VSS 3.35e-20 
C11086 VCC.n7075 VSS 3.5e-20 
C11087 VCC.n7076 VSS 2.36e-19 
C11088 VCC.n7077 VSS 0.0023f 
C11089 VCC.t107 VSS 0.0031f 
C11090 VCC.t307 VSS 0.00366f 
C11091 VCC.t110 VSS 0.00365f 
C11092 VCC.t310 VSS 0.00386f 
C11093 VCC.n7078 VSS 0.00569f 
C11094 VCC.n7079 VSS 1.3e-19 
C11095 VCC.n7080 VSS 3.67e-19 
C11096 VCC.n7081 VSS 1.15e-19 
C11097 VCC.n7082 VSS 3.38e-19 
C11098 VCC.n7083 VSS 3.5e-20 
C11099 VCC.n7084 VSS 3.5e-20 
C11100 VCC.n7085 VSS 2.68e-20 
C11101 VCC.n7086 VSS 2.06e-20 
C11102 VCC.n7087 VSS 6.38e-20 
C11103 VCC.n7088 VSS 5.97e-20 
C11104 VCC.n7089 VSS 4.73e-20 
C11105 VCC.n7090 VSS 4.73e-20 
C11106 VCC.n7091 VSS 3.09e-20 
C11107 VCC.n7092 VSS 1.23e-20 
C11108 VCC.n7093 VSS 1.65e-20 
C11109 VCC.n7094 VSS 1.54e-19 
C11110 VCC.n7095 VSS 1.54e-19 
C11111 VCC.n7096 VSS 1.65e-20 
C11112 VCC.n7097 VSS 3.29e-20 
C11113 VCC.t131 VSS 1.67e-19 
C11114 VCC.n7098 VSS 0.00101f 
C11115 VCC.n7099 VSS 2.71e-19 
C11116 VCC.n7100 VSS 7.46e-19 
C11117 VCC.n7101 VSS 0.00333f 
C11118 VCC.n7102 VSS 2.46e-19 
C11119 VCC.n7103 VSS 3.02e-19 
C11120 VCC.n7104 VSS 3.7e-20 
C11121 VCC.n7105 VSS 5.15e-20 
C11122 VCC.n7106 VSS 5.97e-20 
C11123 VCC.n7107 VSS 6.38e-20 
C11124 VCC.n7108 VSS 4.73e-20 
C11125 VCC.n7109 VSS 4.73e-20 
C11126 VCC.n7110 VSS 2.68e-20 
C11127 VCC.n7111 VSS 3.29e-20 
C11128 VCC.n7112 VSS 1.65e-20 
C11129 VCC.n7113 VSS 1.54e-19 
C11130 VCC.n7114 VSS 1.54e-19 
C11131 VCC.n7115 VSS 1.65e-20 
C11132 VCC.n7116 VSS 3.09e-20 
C11133 VCC.n7117 VSS 3.09e-20 
C11134 VCC.n7118 VSS 4.73e-20 
C11135 VCC.n7119 VSS 4.32e-20 
C11136 VCC.n7120 VSS 3.5e-20 
C11137 VCC.n7121 VSS 3.5e-20 
C11138 VCC.n7122 VSS 1.35e-19 
C11139 VCC.n7123 VSS 5.24e-19 
C11140 VCC.n7124 VSS 1.4e-19 
C11141 VCC.n7125 VSS 5.4e-19 
C11142 VCC.n7126 VSS 1.35e-19 
C11143 VCC.n7127 VSS 4.37e-19 
C11144 VCC.n7128 VSS 1.13e-19 
C11145 VCC.n7129 VSS 8.23e-21 
C11146 VCC.n7130 VSS 1.65e-20 
C11147 VCC.n7131 VSS 3.5e-20 
C11148 VCC.n7132 VSS 3.91e-20 
C11149 VCC.n7133 VSS 3.09e-20 
C11150 VCC.n7134 VSS 1.85e-20 
C11151 VCC.n7135 VSS 3.5e-20 
C11152 VCC.n7136 VSS 1.05e-19 
C11153 VCC.n7137 VSS 2.06e-20 
C11154 VCC.n7138 VSS 2.26e-20 
C11155 VCC.n7139 VSS 3.7e-20 
C11156 VCC.n7140 VSS 5.15e-20 
C11157 VCC.n7141 VSS 1.38e-19 
C11158 VCC.n7142 VSS 1.17e-19 
C11159 VCC.n7143 VSS 4.32e-20 
C11160 VCC.n7144 VSS 2.88e-20 
C11161 VCC.n7145 VSS 2.68e-20 
C11162 VCC.n7146 VSS 6.59e-20 
C11163 VCC.n7147 VSS 5.56e-20 
C11164 VCC.n7148 VSS 2.68e-20 
C11165 VCC.n7149 VSS 4.32e-20 
C11166 VCC.n7150 VSS 1.05e-19 
C11167 VCC.n7151 VSS 3.09e-20 
C11168 VCC.n7152 VSS 3.7e-20 
C11169 VCC.n7153 VSS 4.32e-20 
C11170 VCC.n7154 VSS 1.05e-19 
C11171 VCC.n7155 VSS 4.53e-20 
C11172 VCC.n7156 VSS 4.53e-20 
C11173 VCC.n7157 VSS 7.82e-20 
C11174 VCC.n7158 VSS 2.18e-19 
C11175 VCC.n7159 VSS 1.4e-19 
C11176 VCC.n7160 VSS 1.4e-19 
C11177 VCC.n7161 VSS 5.4e-19 
C11178 VCC.n7162 VSS 1.35e-19 
C11179 VCC.t85 VSS 4.21e-19 
C11180 VCC.n7163 VSS 3.33e-19 
C11181 VCC.n7164 VSS 1.13e-19 
C11182 VCC.n7165 VSS 8.23e-21 
C11183 VCC.n7166 VSS 1.65e-20 
C11184 VCC.n7167 VSS 3.5e-20 
C11185 VCC.n7168 VSS 3.5e-20 
C11186 VCC.n7169 VSS 3.5e-20 
C11187 VCC.n7170 VSS 1.17e-19 
C11188 VCC.n7171 VSS 1.38e-19 
C11189 VCC.n7172 VSS 5.15e-20 
C11190 VCC.n7173 VSS 4.73e-20 
C11191 VCC.n7174 VSS 7.2e-20 
C11192 VCC.n7175 VSS 2.68e-20 
C11193 VCC.n7176 VSS 1.65e-20 
C11194 VCC.n7177 VSS 1.54e-19 
C11195 VCC.n7178 VSS 1.54e-19 
C11196 VCC.n7179 VSS 1.65e-20 
C11197 VCC.n7180 VSS 2.47e-20 
C11198 VCC.n7181 VSS 1.23e-20 
C11199 VCC.n7182 VSS 7.62e-19 
C11200 VCC.n7183 VSS 4.12e-20 
C11201 VCC.n7184 VSS 5.15e-20 
C11202 VCC.n7185 VSS 6.59e-20 
C11203 VCC.n7186 VSS 5.76e-20 
C11204 VCC.n7187 VSS 4.73e-20 
C11205 VCC.n7188 VSS 2.26e-20 
C11206 VCC.n7189 VSS 2.68e-20 
C11207 VCC.n7190 VSS 1.03e-20 
C11208 VCC.n7191 VSS 3.5e-20 
C11209 VCC.n7192 VSS 3.5e-20 
C11210 VCC.n7193 VSS 1.35e-19 
C11211 VCC.n7194 VSS 4.53e-19 
C11212 VCC.n7195 VSS 7.71e-19 
C11213 VCC.n7196 VSS 1.32e-19 
C11214 VCC.n7197 VSS 3.5e-20 
C11215 VCC.n7198 VSS 3.42e-20 
C11216 VCC.n7199 VSS 2.36e-19 
C11217 VCC.n7200 VSS 3.21e-19 
C11218 VCC.n7201 VSS 2.61e-19 
C11219 VCC.n7202 VSS 0.00189f 
C11220 VCC.n7203 VSS 2.68e-19 
C11221 VCC.n7204 VSS 5.76e-20 
C11222 VCC.n7205 VSS 2.88e-20 
C11223 VCC.n7206 VSS 3.5e-20 
C11224 VCC.n7207 VSS 3.42e-20 
C11225 VCC.n7208 VSS 3.5e-20 
C11226 VCC.n7209 VSS 4.53e-19 
C11227 VCC.n7210 VSS 1.17e-19 
C11228 VCC.n7211 VSS 3.5e-20 
C11229 VCC.n7212 VSS 1.44e-20 
C11230 VCC.n7213 VSS 4.12e-20 
C11231 VCC.n7214 VSS 5.76e-20 
C11232 VCC.n7215 VSS 5.76e-20 
C11233 VCC.n7216 VSS 2.06e-20 
C11234 VCC.n7217 VSS 3.29e-20 
C11235 VCC.n7218 VSS 7.2e-20 
C11236 VCC.n7219 VSS 3.29e-20 
C11237 VCC.n7220 VSS 4.73e-20 
C11238 VCC.n7221 VSS 2.26e-20 
C11239 VCC.n7222 VSS 1.01e-19 
C11240 VCC.n7223 VSS 1.36e-19 
C11241 VCC.n7224 VSS 1.35e-19 
C11242 VCC.n7225 VSS 3.5e-20 
C11243 VCC.n7226 VSS 3.5e-20 
C11244 VCC.n7227 VSS 3.5e-20 
C11245 VCC.n7228 VSS 3.5e-20 
C11246 VCC.n7229 VSS 3.09e-20 
C11247 VCC.n7230 VSS 3.91e-20 
C11248 VCC.n7231 VSS 4.73e-20 
C11249 VCC.n7232 VSS 4.32e-20 
C11250 VCC.n7233 VSS 2.68e-20 
C11251 VCC.n7234 VSS 4.53e-20 
C11252 VCC.n7235 VSS 4.53e-20 
C11253 VCC.n7236 VSS 3.09e-20 
C11254 VCC.n7237 VSS 4.32e-20 
C11255 VCC.n7238 VSS 2.68e-20 
C11256 VCC.n7239 VSS 7.82e-20 
C11257 VCC.n7240 VSS 5.56e-20 
C11258 VCC.n7241 VSS 1.4e-19 
C11259 VCC.n7242 VSS 2.18e-19 
C11260 VCC.n7243 VSS 1.35e-19 
C11261 VCC.n7244 VSS 1.13e-19 
C11262 VCC.n7245 VSS 3.5e-20 
C11263 VCC.n7246 VSS 1.85e-20 
C11264 VCC.n7247 VSS 3.7e-20 
C11265 VCC.n7248 VSS 3.09e-20 
C11266 VCC.n7249 VSS 6.59e-20 
C11267 VCC.n7250 VSS 2.68e-20 
C11268 VCC.n7251 VSS 5.76e-20 
C11269 VCC.n7252 VSS 4.73e-20 
C11270 VCC.n7253 VSS 3.5e-20 
C11271 VCC.t70 VSS 1.56e-19 
C11272 VCC.n7254 VSS 7.97e-19 
C11273 VCC.n7255 VSS 3.09e-20 
C11274 VCC.n7256 VSS 3.5e-20 
C11275 VCC.n7257 VSS 3.5e-20 
C11276 VCC.t69 VSS 4.21e-19 
C11277 VCC.n7258 VSS 1.32e-19 
C11278 VCC.n7259 VSS 1.09e-19 
C11279 VCC.n7260 VSS 3.5e-20 
C11280 VCC.n7261 VSS 3.09e-20 
C11281 VCC.n7262 VSS 5.97e-20 
C11282 VCC.n7263 VSS 2.26e-20 
C11283 VCC.n7264 VSS 5.76e-20 
C11284 VCC.n7265 VSS 2.68e-20 
C11285 VCC.n7266 VSS 2.68e-20 
C11286 VCC.n7267 VSS 1.9e-19 
C11287 VCC.n7268 VSS 5.76e-20 
C11288 VCC.n7269 VSS 2.68e-20 
C11289 VCC.n7270 VSS 2.68e-20 
C11290 VCC.n7271 VSS 2.68e-20 
C11291 VCC.n7272 VSS 5.76e-20 
C11292 VCC.n7273 VSS 2.26e-20 
C11293 VCC.n7274 VSS 3.09e-20 
C11294 VCC.n7275 VSS 2.26e-20 
C11295 VCC.n7276 VSS 5.15e-20 
C11296 VCC.n7277 VSS 4.73e-20 
C11297 VCC.n7278 VSS 3.7e-20 
C11298 VCC.n7279 VSS 3.5e-20 
C11299 VCC.n7280 VSS 7.41e-20 
C11300 VCC.n7281 VSS 1.91e-19 
C11301 VCC.n7282 VSS 9.88e-20 
C11302 VCC.n7283 VSS 3e-20 
C11303 VCC.n7284 VSS 5.12e-19 
C11304 VCC.n7285 VSS 1.18e-19 
C11305 VCC.n7286 VSS 3.5e-20 
C11306 VCC.n7287 VSS 3.5e-20 
C11307 VCC.n7288 VSS 5.15e-20 
C11308 VCC.n7289 VSS 4.32e-20 
C11309 VCC.n7290 VSS 2.68e-20 
C11310 VCC.n7291 VSS 3.91e-20 
C11311 VCC.n7292 VSS 1.44e-20 
C11312 VCC.n7293 VSS 3.5e-20 
C11313 VCC.n7294 VSS 3e-20 
C11314 VCC.n7295 VSS 7.95e-19 
C11315 VCC.n7296 VSS 1.83e-19 
C11316 VCC.n7297 VSS 2.88e-20 
C11317 VCC.n7298 VSS 2.68e-20 
C11318 VCC.n7299 VSS 2.68e-20 
C11319 VCC.n7300 VSS 2.68e-20 
C11320 VCC.n7301 VSS 4.53e-20 
C11321 VCC.n7302 VSS 3.7e-20 
C11322 VCC.n7303 VSS 7.82e-20 
C11323 VCC.n7304 VSS 1.17e-19 
C11324 VCC.n7305 VSS 3.91e-20 
C11325 VCC.n7306 VSS 1.65e-20 
C11326 VCC.n7307 VSS 2.68e-20 
C11327 VCC.n7308 VSS 3.5e-20 
C11328 VCC.n7309 VSS 3e-20 
C11329 VCC.n7310 VSS 5.12e-19 
C11330 VCC.n7311 VSS 1.18e-19 
C11331 VCC.n7312 VSS 3.5e-20 
C11332 VCC.n7313 VSS 3.5e-20 
C11333 VCC.t280 VSS 1.55e-19 
C11334 VCC.n7314 VSS 7.57e-19 
C11335 VCC.n7315 VSS 4.73e-20 
C11336 VCC.n7316 VSS 1.54e-19 
C11337 VCC.n7317 VSS 2.88e-20 
C11338 VCC.n7318 VSS 2.88e-20 
C11339 VCC.n7319 VSS 3.5e-20 
C11340 VCC.n7320 VSS 5.76e-20 
C11341 VCC.n7321 VSS 9.88e-20 
C11342 VCC.n7322 VSS 1.3e-19 
C11343 VCC.n7323 VSS 3e-20 
C11344 VCC.t281 VSS 0.005f 
C11345 VCC.t119 VSS 0.00453f 
C11346 VCC.n7324 VSS 0.00229f 
C11347 VCC.n7325 VSS 1.91e-19 
C11348 VCC.n7326 VSS 3.5e-20 
C11349 VCC.n7327 VSS 3.14e-19 
C11350 VCC.n7328 VSS 2.47e-20 
C11351 VCC.n7329 VSS 5.76e-20 
C11352 VCC.n7330 VSS 2.47e-20 
C11353 VCC.n7331 VSS 8.23e-21 
C11354 VCC.n7332 VSS 2.88e-20 
C11355 VCC.n7333 VSS 5.76e-20 
C11356 VCC.n7334 VSS 2.47e-20 
C11357 VCC.n7335 VSS 2.88e-20 
C11358 VCC.n7336 VSS 2.47e-20 
C11359 VCC.n7337 VSS 5.15e-20 
C11360 VCC.n7338 VSS 4.73e-20 
C11361 VCC.n7339 VSS 3.7e-20 
C11362 VCC.n7340 VSS 3.5e-20 
C11363 VCC.n7341 VSS 7.41e-20 
C11364 VCC.t172 VSS 6.42e-19 
C11365 VCC.n7342 VSS 3e-20 
C11366 VCC.n7343 VSS 5.97e-20 
C11367 VCC.n7344 VSS 4.13e-19 
C11368 VCC.n7345 VSS 9.53e-20 
C11369 VCC.n7346 VSS 3.5e-20 
C11370 VCC.n7347 VSS 3.5e-20 
C11371 VCC.n7348 VSS 5.35e-20 
C11372 VCC.n7349 VSS 4.32e-20 
C11373 VCC.n7350 VSS 2.68e-20 
C11374 VCC.n7351 VSS 3.7e-20 
C11375 VCC.n7352 VSS 1.65e-20 
C11376 VCC.n7353 VSS 4.53e-20 
C11377 VCC.n7354 VSS 1.2e-19 
C11378 VCC.n7355 VSS 5.2e-19 
C11379 VCC.n7356 VSS 1.2e-19 
C11380 VCC.n7357 VSS 6.38e-20 
C11381 VCC.n7358 VSS 2.47e-20 
C11382 VCC.n7359 VSS 4.53e-20 
C11383 VCC.n7360 VSS 3.5e-20 
C11384 VCC.n7361 VSS 3.5e-20 
C11385 VCC.n7362 VSS 2.68e-20 
C11386 VCC.n7363 VSS 2.68e-20 
C11387 VCC.n7364 VSS 2.47e-20 
C11388 VCC.n7365 VSS 4.53e-20 
C11389 VCC.n7366 VSS 2.68e-20 
C11390 VCC.n7367 VSS 4.32e-20 
C11391 VCC.n7368 VSS 2.68e-20 
C11392 VCC.n7369 VSS 3.91e-20 
C11393 VCC.n7370 VSS 2.88e-20 
C11394 VCC.n7371 VSS 4.73e-20 
C11395 VCC.n7372 VSS 3.7e-20 
C11396 VCC.n7373 VSS 3.7e-20 
C11397 VCC.n7374 VSS 3.5e-20 
C11398 VCC.n7375 VSS 5.76e-20 
C11399 VCC.n7376 VSS 4.73e-20 
C11400 VCC.n7377 VSS 3.09e-20 
C11401 VCC.n7378 VSS 3.5e-20 
C11402 VCC.n7379 VSS 3.5e-20 
C11403 VCC.n7380 VSS 3.5e-20 
C11404 VCC.n7381 VSS 1.18e-19 
C11405 VCC.n7382 VSS 3e-20 
C11406 VCC.n7383 VSS 1.15e-19 
C11407 VCC.n7384 VSS 9.88e-20 
C11408 VCC.n7385 VSS 5.76e-20 
C11409 VCC.n7386 VSS 3.5e-20 
C11410 VCC.n7387 VSS 3.09e-20 
C11411 VCC.n7388 VSS 3.09e-20 
C11412 VCC.n7389 VSS 2.26e-20 
C11413 VCC.n7390 VSS 5.76e-20 
C11414 VCC.n7391 VSS 2.68e-20 
C11415 VCC.n7392 VSS 2.68e-20 
C11416 VCC.n7393 VSS 0.00185f 
C11417 VCC.n7394 VSS 2.72e-19 
C11418 VCC.n7395 VSS 2.26e-20 
C11419 VCC.n7396 VSS 1.87e-19 
C11420 VCC.n7397 VSS 3.5e-20 
C11421 VCC.n7398 VSS 2.68e-20 
C11422 VCC.n7399 VSS 5.97e-20 
C11423 VCC.n7400 VSS 4.73e-20 
C11424 VCC.n7401 VSS 4.73e-20 
C11425 VCC.n7402 VSS 5.15e-20 
C11426 VCC.n7403 VSS 7.41e-20 
C11427 VCC.n7404 VSS 3.7e-20 
C11428 VCC.n7405 VSS 2.26e-20 
C11429 VCC.n7406 VSS 6.38e-20 
C11430 VCC.n7407 VSS 4.73e-20 
C11431 VCC.n7408 VSS 3.29e-20 
C11432 VCC.n7409 VSS 3.5e-20 
C11433 VCC.n7410 VSS 3e-20 
C11434 VCC.t11 VSS 0.005f 
C11435 VCC.t48 VSS 0.00453f 
C11436 VCC.n7411 VSS 0.00228f 
C11437 VCC.n7412 VSS 1.3e-19 
C11438 VCC.t12 VSS 4.05e-19 
C11439 VCC.n7413 VSS 4.05e-19 
C11440 VCC.n7414 VSS 1.15e-19 
C11441 VCC.n7415 VSS 3.36e-19 
C11442 VCC.n7416 VSS 6.17e-21 
C11443 VCC.n7417 VSS 3.12e-19 
C11444 VCC.n7418 VSS 1.65e-20 
C11445 VCC.n7419 VSS 1.54e-19 
C11446 VCC.n7420 VSS 1.54e-19 
C11447 VCC.n7421 VSS 1.65e-20 
C11448 VCC.n7422 VSS 1.03e-20 
C11449 VCC.n7423 VSS 3.5e-20 
C11450 VCC.n7424 VSS 2.26e-20 
C11451 VCC.n7425 VSS 4.73e-20 
C11452 VCC.n7426 VSS 3.5e-20 
C11453 VCC.n7427 VSS 3e-20 
C11454 VCC.n7428 VSS 1.3e-19 
C11455 VCC.n7429 VSS 5.12e-19 
C11456 VCC.n7430 VSS 1.3e-19 
C11457 VCC.n7431 VSS 4.13e-19 
C11458 VCC.n7432 VSS 9.53e-20 
C11459 VCC.n7433 VSS 5.76e-20 
C11460 VCC.n7434 VSS 7.41e-20 
C11461 VCC.n7435 VSS 5.56e-20 
C11462 VCC.t13 VSS 1.55e-19 
C11463 VCC.n7436 VSS 3.91e-20 
C11464 VCC.n7437 VSS 3.91e-20 
C11465 VCC.n7438 VSS 1.85e-20 
C11466 VCC.n7439 VSS 7.55e-19 
C11467 VCC.n7440 VSS 4.94e-20 
C11468 VCC.n7441 VSS 5.15e-20 
C11469 VCC.n7442 VSS 7.2e-20 
C11470 VCC.n7443 VSS 1.38e-19 
C11471 VCC.n7444 VSS 1.17e-19 
C11472 VCC.n7445 VSS 4.32e-20 
C11473 VCC.n7446 VSS 2.88e-20 
C11474 VCC.n7447 VSS 2.68e-20 
C11475 VCC.n7448 VSS 3.5e-20 
C11476 VCC.n7449 VSS 3.5e-20 
C11477 VCC.n7450 VSS 2.88e-20 
C11478 VCC.n7451 VSS 2.68e-20 
C11479 VCC.n7452 VSS 2.68e-20 
C11480 VCC.n7453 VSS 2.68e-20 
C11481 VCC.n7454 VSS 4.12e-20 
C11482 VCC.n7455 VSS 4.12e-20 
C11483 VCC.n7456 VSS 3.91e-20 
C11484 VCC.n7457 VSS 4.53e-20 
C11485 VCC.n7458 VSS 4.53e-20 
C11486 VCC.n7459 VSS 1.05e-19 
C11487 VCC.n7460 VSS 1.05e-19 
C11488 VCC.n7461 VSS 4.32e-20 
C11489 VCC.n7462 VSS 3.7e-20 
C11490 VCC.n7463 VSS 2.68e-20 
C11491 VCC.n7464 VSS 2.68e-20 
C11492 VCC.n7465 VSS 6.79e-20 
C11493 VCC.n7466 VSS 9.26e-20 
C11494 VCC.n7467 VSS 1.83e-19 
C11495 VCC.n7468 VSS 7.95e-19 
C11496 VCC.n7469 VSS 5.2e-19 
C11497 VCC.n7470 VSS 1.3e-19 
C11498 VCC.n7471 VSS 3e-20 
C11499 VCC.n7472 VSS 3.5e-20 
C11500 VCC.n7473 VSS 5.97e-20 
C11501 VCC.n7474 VSS 7.41e-20 
C11502 VCC.n7475 VSS 5.15e-20 
C11503 VCC.n7476 VSS 5.15e-20 
C11504 VCC.n7477 VSS 3.09e-20 
C11505 VCC.n7478 VSS 3.09e-20 
C11506 VCC.n7479 VSS 3.7e-20 
C11507 VCC.n7480 VSS 2.68e-20 
C11508 VCC.n7481 VSS 3.91e-20 
C11509 VCC.n7482 VSS 1.17e-19 
C11510 VCC.n7483 VSS 1.38e-19 
C11511 VCC.n7484 VSS 7e-20 
C11512 VCC.n7485 VSS 4.73e-20 
C11513 VCC.n7486 VSS 3.5e-20 
C11514 VCC.n7487 VSS 3.5e-20 
C11515 VCC.n7488 VSS 3.5e-20 
C11516 VCC.n7489 VSS 4.53e-20 
C11517 VCC.n7490 VSS 1.18e-19 
C11518 VCC.n7491 VSS 5.12e-19 
C11519 VCC.n7492 VSS 1.3e-19 
C11520 VCC.n7493 VSS 1.61e-19 
C11521 VCC.n7494 VSS 9.9e-20 
C11522 VCC.n7495 VSS 0.00243f 
C11523 VCC.n7496 VSS 2.26e-20 
C11524 VCC.n7497 VSS 4.13e-19 
C11525 VCC.n7498 VSS 3.5e-20 
C11526 VCC.n7499 VSS 3.5e-20 
C11527 VCC.n7500 VSS 2.47e-20 
C11528 VCC.n7501 VSS 2.06e-20 
C11529 VCC.n7502 VSS 6.17e-20 
C11530 VCC.n7503 VSS 6.17e-20 
C11531 VCC.n7504 VSS 4.73e-20 
C11532 VCC.n7505 VSS 4.73e-20 
C11533 VCC.n7506 VSS 2.88e-20 
C11534 VCC.n7507 VSS 1.44e-20 
C11535 VCC.n7508 VSS 1.65e-20 
C11536 VCC.n7509 VSS 1.54e-19 
C11537 VCC.n7510 VSS 1.54e-19 
C11538 VCC.n7511 VSS 1.65e-20 
C11539 VCC.n7512 VSS 3.09e-20 
C11540 VCC.t173 VSS 1.55e-19 
C11541 VCC.n7513 VSS 0.00102f 
C11542 VCC.n7514 VSS 2.73e-19 
C11543 VCC.n7515 VSS 0.00136f 
C11544 VCC.n7516 VSS 2.73e-19 
C11545 VCC.n7517 VSS 0.00181f 
C11546 VCC.n7518 VSS 5.76e-20 
C11547 VCC.n7519 VSS 1.54e-19 
C11548 VCC.n7520 VSS 1.65e-20 
C11549 VCC.n7521 VSS 2.88e-20 
C11550 VCC.n7522 VSS 2.47e-20 
C11551 VCC.n7523 VSS 6.17e-20 
C11552 VCC.n7524 VSS 4.73e-20 
C11553 VCC.n7525 VSS 4.73e-20 
C11554 VCC.n7526 VSS 5.15e-20 
C11555 VCC.n7527 VSS 3.5e-20 
C11556 VCC.n7528 VSS 7.41e-20 
C11557 VCC.n7529 VSS 3.7e-20 
C11558 VCC.n7530 VSS 2.26e-20 
C11559 VCC.n7531 VSS 6.17e-20 
C11560 VCC.n7532 VSS 4.73e-20 
C11561 VCC.n7533 VSS 3.5e-20 
C11562 VCC.n7534 VSS 2.88e-20 
C11563 VCC.n7535 VSS 3.4e-19 
C11564 VCC.n7536 VSS 1.15e-19 
C11565 VCC.n7537 VSS 3.98e-19 
C11566 VCC.t279 VSS 4.05e-19 
C11567 VCC.n7538 VSS 1.22e-19 
C11568 VCC.n7539 VSS 1.3e-19 
C11569 VCC.n7540 VSS 3e-20 
C11570 VCC.n7541 VSS 3.5e-20 
C11571 VCC.n7542 VSS 3.5e-20 
C11572 VCC.n7543 VSS 4.73e-20 
C11573 VCC.n7544 VSS 2.47e-20 
C11574 VCC.n7545 VSS 1.23e-20 
C11575 VCC.n7546 VSS 1.65e-20 
C11576 VCC.n7547 VSS 2.47e-20 
C11577 VCC.n7548 VSS 5.76e-20 
C11578 VCC.n7549 VSS 1.38e-19 
C11579 VCC.n7550 VSS 7e-20 
C11580 VCC.n7551 VSS 3.7e-20 
C11581 VCC.n7552 VSS 2.47e-20 
C11582 VCC.n7553 VSS 3.7e-20 
C11583 VCC.n7554 VSS 1.85e-20 
C11584 VCC.n7555 VSS 3.09e-20 
C11585 VCC.n7556 VSS 5.35e-20 
C11586 VCC.n7557 VSS 4.73e-20 
C11587 VCC.n7558 VSS 5.35e-20 
C11588 VCC.n7559 VSS 7.41e-20 
C11589 VCC.n7560 VSS 5.76e-20 
C11590 VCC.n7561 VSS 9.53e-20 
C11591 VCC.n7562 VSS 4.13e-19 
C11592 VCC.n7563 VSS 1.3e-19 
C11593 VCC.n7564 VSS 5.2e-19 
C11594 VCC.n7565 VSS 1.2e-19 
C11595 VCC.n7566 VSS 4.73e-20 
C11596 VCC.n7567 VSS 2.68e-20 
C11597 VCC.n7568 VSS 3.5e-20 
C11598 VCC.n7569 VSS 3.5e-20 
C11599 VCC.n7570 VSS 2.68e-20 
C11600 VCC.n7571 VSS 2.68e-20 
C11601 VCC.n7572 VSS 4.32e-20 
C11602 VCC.n7573 VSS 4.32e-20 
C11603 VCC.n7574 VSS 4.32e-20 
C11604 VCC.n7575 VSS 2.88e-20 
C11605 VCC.n7576 VSS 3.5e-20 
C11606 VCC.n7577 VSS 2.68e-20 
C11607 VCC.n7578 VSS 7.82e-20 
C11608 VCC.n7579 VSS 4.73e-20 
C11609 VCC.n7580 VSS 4.73e-20 
C11610 VCC.n7581 VSS 1.05e-19 
C11611 VCC.n7582 VSS 1.05e-19 
C11612 VCC.n7583 VSS 4.53e-20 
C11613 VCC.n7584 VSS 2.68e-20 
C11614 VCC.n7585 VSS 2.68e-20 
C11615 VCC.n7586 VSS 6.59e-20 
C11616 VCC.n7587 VSS 9.26e-20 
C11617 VCC.n7588 VSS 6.59e-20 
C11618 VCC.n7589 VSS 2.47e-20 
C11619 VCC.n7590 VSS 2.47e-20 
C11620 VCC.n7591 VSS 2.88e-20 
C11621 VCC.n7592 VSS 3.5e-20 
C11622 VCC.n7593 VSS 3.5e-20 
C11623 VCC.n7594 VSS 4.53e-20 
C11624 VCC.n7595 VSS 1.2e-19 
C11625 VCC.n7596 VSS 5.2e-19 
C11626 VCC.n7597 VSS 1.3e-19 
C11627 VCC.n7598 VSS 4.13e-19 
C11628 VCC.n7599 VSS 9.53e-20 
C11629 VCC.n7600 VSS 5.97e-20 
C11630 VCC.n7601 VSS 7.41e-20 
C11631 VCC.n7602 VSS 5.35e-20 
C11632 VCC.n7603 VSS 5.15e-20 
C11633 VCC.n7604 VSS 3.09e-20 
C11634 VCC.n7605 VSS 3.09e-20 
C11635 VCC.n7606 VSS 3.91e-20 
C11636 VCC.n7607 VSS 2.47e-20 
C11637 VCC.n7608 VSS 3.7e-20 
C11638 VCC.n7609 VSS 1.17e-19 
C11639 VCC.n7610 VSS 1.38e-19 
C11640 VCC.n7611 VSS 7.2e-20 
C11641 VCC.n7612 VSS 4.73e-20 
C11642 VCC.n7613 VSS 3.5e-20 
C11643 VCC.n7614 VSS 3.5e-20 
C11644 VCC.n7615 VSS 4.53e-20 
C11645 VCC.n7616 VSS 5.97e-20 
C11646 VCC.n7617 VSS 3.5e-20 
C11647 VCC.n7618 VSS 3e-20 
C11648 VCC.n7619 VSS 1.3e-19 
C11649 VCC.n7620 VSS 1.53e-19 
C11650 VCC.t63 VSS 4.05e-19 
C11651 VCC.n7621 VSS 2.06e-19 
C11652 VCC.n7622 VSS 1.35e-19 
C11653 VCC.n7623 VSS 9.67e-20 
C11654 VCC.n7624 VSS 3.35e-20 
C11655 VCC.n7625 VSS 3.5e-20 
C11656 VCC.n7626 VSS 2.36e-19 
C11657 VCC.n7627 VSS 0.0023f 
C11658 VCC.t72 VSS 0.0031f 
C11659 VCC.t38 VSS 0.00366f 
C11660 VCC.t71 VSS 0.00365f 
C11661 VCC.t37 VSS 0.00386f 
C11662 VCC.n7628 VSS 0.00569f 
C11663 VCC.n7629 VSS 1.3e-19 
C11664 VCC.n7630 VSS 3.67e-19 
C11665 VCC.n7631 VSS 1.15e-19 
C11666 VCC.n7632 VSS 3.38e-19 
C11667 VCC.n7633 VSS 3.5e-20 
C11668 VCC.n7634 VSS 3.5e-20 
C11669 VCC.n7635 VSS 2.68e-20 
C11670 VCC.n7636 VSS 2.06e-20 
C11671 VCC.n7637 VSS 6.38e-20 
C11672 VCC.n7638 VSS 5.97e-20 
C11673 VCC.n7639 VSS 4.73e-20 
C11674 VCC.n7640 VSS 4.73e-20 
C11675 VCC.n7641 VSS 3.09e-20 
C11676 VCC.n7642 VSS 1.23e-20 
C11677 VCC.n7643 VSS 1.65e-20 
C11678 VCC.n7644 VSS 1.54e-19 
C11679 VCC.n7645 VSS 1.54e-19 
C11680 VCC.n7646 VSS 1.65e-20 
C11681 VCC.n7647 VSS 3.29e-20 
C11682 VCC.t64 VSS 1.67e-19 
C11683 VCC.n7648 VSS 0.00101f 
C11684 VCC.n7649 VSS 2.71e-19 
C11685 VCC.n7650 VSS 7.46e-19 
C11686 VCC.n7651 VSS 0.00333f 
C11687 VCC.n7652 VSS 2.46e-19 
C11688 VCC.n7653 VSS 3.02e-19 
C11689 VCC.n7654 VSS 3.7e-20 
C11690 VCC.n7655 VSS 5.15e-20 
C11691 VCC.n7656 VSS 6.38e-20 
C11692 VCC.n7657 VSS 4.73e-20 
C11693 VCC.n7658 VSS 4.73e-20 
C11694 VCC.n7659 VSS 2.68e-20 
C11695 VCC.n7660 VSS 3.29e-20 
C11696 VCC.n7661 VSS 1.65e-20 
C11697 VCC.n7662 VSS 1.54e-19 
C11698 VCC.n7663 VSS 1.54e-19 
C11699 VCC.n7664 VSS 5.56e-20 
C11700 VCC.n7665 VSS 2.88e-20 
C11701 VCC.n7666 VSS 1.65e-20 
C11702 VCC.n7667 VSS 3.09e-20 
C11703 VCC.n7668 VSS 4.73e-20 
C11704 VCC.n7669 VSS 4.73e-20 
C11705 VCC.n7670 VSS 4.32e-20 
C11706 VCC.n7671 VSS 1.17e-19 
C11707 VCC.n7672 VSS 3.33e-19 
C11708 VCC.n7673 VSS 1.35e-19 
C11709 VCC.n7674 VSS 4.37e-19 
C11710 VCC.n7675 VSS 5.24e-19 
C11711 VCC.n7676 VSS 1.36e-19 
C11712 VCC.n7677 VSS 1.01e-19 
C11713 VCC.n7678 VSS 1.05e-19 
C11714 VCC.n7679 VSS 2.06e-20 
C11715 VCC.n7680 VSS 2.26e-20 
C11716 VCC.n7681 VSS 3.7e-20 
C11717 VCC.n7682 VSS 5.15e-20 
C11718 VCC.n7683 VSS 1.38e-19 
C11719 VCC.n7684 VSS 3.91e-20 
C11720 VCC.n7685 VSS 2.88e-20 
C11721 VCC.n7686 VSS 4.32e-20 
C11722 VCC.n7687 VSS 1.17e-19 
C11723 VCC.n7688 VSS 3.7e-20 
C11724 VCC.n7689 VSS 3.91e-20 
C11725 VCC.n7690 VSS 3.5e-20 
C11726 VCC.n7691 VSS 1.65e-20 
C11727 VCC.n7692 VSS 8.23e-21 
C11728 VCC.n7693 VSS 3.5e-20 
C11729 VCC.n7694 VSS 3.5e-20 
C11730 VCC.n7695 VSS 1.4e-19 
C11731 VCC.n7696 VSS 5.4e-19 
C11732 VCC.n7697 VSS 8.42e-19 
C11733 VCC.n7698 VSS 5.4e-19 
C11734 VCC.n7699 VSS 1.4e-19 
C11735 VCC.n7700 VSS 1.4e-19 
C11736 VCC.n7701 VSS 2.18e-19 
C11737 VCC.n7702 VSS 7.82e-20 
C11738 VCC.n7703 VSS 4.32e-20 
C11739 VCC.n7704 VSS 4.32e-20 
C11740 VCC.n7705 VSS 1.05e-19 
C11741 VCC.n7706 VSS 1.05e-19 
C11742 VCC.n7707 VSS 4.32e-20 
C11743 VCC.n7708 VSS 3.7e-20 
C11744 VCC.n7709 VSS 2.68e-20 
C11745 VCC.n7710 VSS 5.76e-20 
C11746 VCC.n7711 VSS 6.38e-20 
C11747 VCC.n7712 VSS 3.5e-20 
C11748 VCC.n7713 VSS 3.5e-20 
C11749 VCC.n7714 VSS 1.17e-19 
C11750 VCC.n7715 VSS 1.38e-19 
C11751 VCC.n7716 VSS 5.15e-20 
C11752 VCC.n7717 VSS 1.05e-19 
C11753 VCC.n7718 VSS 2.26e-20 
C11754 VCC.n7719 VSS 5.76e-20 
C11755 VCC.n7720 VSS 3.7e-20 
C11756 VCC.n7721 VSS 3.7e-20 
C11757 VCC.n7722 VSS 3.09e-20 
C11758 VCC.n7723 VSS 1.85e-20 
C11759 VCC.n7724 VSS 1.65e-20 
C11760 VCC.n7725 VSS 8.23e-21 
C11761 VCC.n7726 VSS 1.13e-19 
C11762 VCC.n7727 VSS 3.33e-19 
C11763 VCC.t308 VSS 4.21e-19 
C11764 VCC.n7728 VSS 2.06e-19 
C11765 VCC.n7729 VSS 1.35e-19 
C11766 VCC.n7730 VSS 3.5e-20 
C11767 VCC.n7731 VSS 3.5e-20 
C11768 VCC.n7732 VSS 3.5e-20 
C11769 VCC.n7733 VSS 1.03e-20 
C11770 VCC.n7734 VSS 2.68e-20 
C11771 VCC.n7735 VSS 3.09e-20 
C11772 VCC.n7736 VSS 2.68e-20 
C11773 VCC.n7737 VSS 1.65e-20 
C11774 VCC.n7738 VSS 1.54e-19 
C11775 VCC.n7739 VSS 1.54e-19 
C11776 VCC.n7740 VSS 1.65e-20 
C11777 VCC.t309 VSS 1.56e-19 
C11778 VCC.n7741 VSS 7.62e-19 
C11779 VCC.n7742 VSS 1.23e-20 
C11780 VCC.n7743 VSS 2.47e-20 
C11781 VCC.n7744 VSS 4.73e-20 
C11782 VCC.n7745 VSS 6.59e-20 
C11783 VCC.n7746 VSS 5.15e-20 
C11784 VCC.n7747 VSS 2.47e-20 
C11785 VCC.n7748 VSS 7.41e-20 
C11786 VCC.n7749 VSS 9.47e-20 
C11787 VCC.n7750 VSS 1.32e-19 
C11788 VCC.n7751 VSS 7.71e-19 
C11789 VCC.n7752 VSS 9.83e-19 
C11790 VCC.n7753 VSS 2.36e-19 
C11791 VCC.n7754 VSS 3.21e-19 
C11792 VCC.n7755 VSS 2.61e-19 
C11793 VCC.n7756 VSS 0.00189f 
C11794 VCC.n7757 VSS 5.76e-20 
C11795 VCC.n7758 VSS 2.88e-20 
C11796 VCC.n7759 VSS 3.5e-20 
C11797 VCC.n7760 VSS 9.83e-19 
C11798 VCC.n7761 VSS 9.47e-20 
C11799 VCC.n7762 VSS 1.17e-19 
C11800 VCC.n7763 VSS 2.06e-19 
C11801 VCC.n7764 VSS 1.36e-19 
C11802 VCC.n7765 VSS 1.01e-19 
C11803 VCC.n7766 VSS 3.5e-20 
C11804 VCC.n7767 VSS 3.09e-20 
C11805 VCC.n7768 VSS 3.29e-20 
C11806 VCC.n7769 VSS 3.29e-20 
C11807 VCC.n7770 VSS 4.73e-20 
C11808 VCC.n7771 VSS 1.44e-20 
C11809 VCC.n7772 VSS 3.5e-20 
C11810 VCC.n7773 VSS 7.41e-20 
C11811 VCC.n7774 VSS 2.47e-20 
C11812 VCC.t40 VSS 1.56e-19 
C11813 VCC.n7775 VSS 5.76e-20 
C11814 VCC.n7776 VSS 2.06e-20 
C11815 VCC.n7777 VSS 5.76e-20 
C11816 VCC.n7778 VSS 3.7e-20 
C11817 VCC.n7779 VSS 4.32e-20 
C11818 VCC.n7780 VSS 2.68e-20 
C11819 VCC.n7781 VSS 3.91e-20 
C11820 VCC.n7782 VSS 6.38e-20 
C11821 VCC.n7783 VSS 1.85e-20 
C11822 VCC.n7784 VSS 3.5e-20 
C11823 VCC.n7785 VSS 3.09e-20 
C11824 VCC.n7786 VSS 3.7e-20 
C11825 VCC.n7787 VSS 3.09e-20 
C11826 VCC.n7788 VSS 2.26e-20 
C11827 VCC.n7789 VSS 1.05e-19 
C11828 VCC.n7790 VSS 3.5e-20 
C11829 VCC.n7791 VSS 3.5e-20 
C11830 VCC.n7792 VSS 8.42e-19 
C11831 VCC.n7793 VSS 2.18e-19 
C11832 VCC.n7794 VSS 1.4e-19 
C11833 VCC.n7795 VSS 4.32e-20 
C11834 VCC.n7796 VSS 7.82e-20 
C11835 VCC.n7797 VSS 5.76e-20 
C11836 VCC.n7798 VSS 2.68e-20 
C11837 VCC.n7799 VSS 4.32e-20 
C11838 VCC.n7800 VSS 3.91e-20 
C11839 VCC.n7801 VSS 3.7e-20 
C11840 VCC.n7802 VSS 3.7e-20 
C11841 VCC.n7803 VSS 5.76e-20 
C11842 VCC.n7804 VSS 4.73e-20 
C11843 VCC.n7805 VSS 3.5e-20 
C11844 VCC.t219 VSS 1.56e-19 
C11845 VCC.n7806 VSS 7.97e-19 
C11846 VCC.n7807 VSS 3.09e-20 
C11847 VCC.n7808 VSS 1.01e-19 
C11848 VCC.n7809 VSS 3.5e-20 
C11849 VCC.n7810 VSS 1.36e-19 
C11850 VCC.n7811 VSS 3.5e-20 
C11851 VCC.n7812 VSS 3.33e-19 
C11852 VCC.n7813 VSS 1.17e-19 
C11853 VCC.n7814 VSS 1.09e-19 
C11854 VCC.n7815 VSS 3.5e-20 
C11855 VCC.n7816 VSS 4.73e-20 
C11856 VCC.n7817 VSS 5.56e-20 
C11857 VCC.n7818 VSS 2.88e-20 
C11858 VCC.n7819 VSS 2.26e-20 
C11859 VCC.n7820 VSS 5.76e-20 
C11860 VCC.n7821 VSS 2.68e-20 
C11861 VCC.n7822 VSS 2.68e-20 
C11862 VCC.n7823 VSS 1.9e-19 
C11863 VCC.n7824 VSS 5.76e-20 
C11864 VCC.n7825 VSS 2.68e-20 
C11865 VCC.n7826 VSS 2.68e-20 
C11866 VCC.n7827 VSS 2.68e-20 
C11867 VCC.n7828 VSS 5.76e-20 
C11868 VCC.n7829 VSS 2.26e-20 
C11869 VCC.n7830 VSS 3.09e-20 
C11870 VCC.n7831 VSS 2.26e-20 
C11871 VCC.n7832 VSS 5.15e-20 
C11872 VCC.n7833 VSS 4.73e-20 
C11873 VCC.n7834 VSS 3.7e-20 
C11874 VCC.n7835 VSS 3.5e-20 
C11875 VCC.n7836 VSS 7.41e-20 
C11876 VCC.n7837 VSS 1.91e-19 
C11877 VCC.n7838 VSS 9.88e-20 
C11878 VCC.n7839 VSS 3e-20 
C11879 VCC.n7840 VSS 5.12e-19 
C11880 VCC.n7841 VSS 1.18e-19 
C11881 VCC.n7842 VSS 3.5e-20 
C11882 VCC.n7843 VSS 3.5e-20 
C11883 VCC.n7844 VSS 5.15e-20 
C11884 VCC.n7845 VSS 4.32e-20 
C11885 VCC.n7846 VSS 2.68e-20 
C11886 VCC.n7847 VSS 3.91e-20 
C11887 VCC.n7848 VSS 1.44e-20 
C11888 VCC.n7849 VSS 3.5e-20 
C11889 VCC.n7850 VSS 3e-20 
C11890 VCC.n7851 VSS 7.95e-19 
C11891 VCC.n7852 VSS 1.83e-19 
C11892 VCC.n7853 VSS 2.88e-20 
C11893 VCC.n7854 VSS 2.68e-20 
C11894 VCC.n7855 VSS 2.68e-20 
C11895 VCC.n7856 VSS 2.68e-20 
C11896 VCC.n7857 VSS 4.53e-20 
C11897 VCC.n7858 VSS 3.7e-20 
C11898 VCC.n7859 VSS 7.82e-20 
C11899 VCC.n7860 VSS 1.17e-19 
C11900 VCC.n7861 VSS 3.91e-20 
C11901 VCC.n7862 VSS 1.65e-20 
C11902 VCC.n7863 VSS 2.68e-20 
C11903 VCC.n7864 VSS 3.5e-20 
C11904 VCC.n7865 VSS 3e-20 
C11905 VCC.n7866 VSS 5.12e-19 
C11906 VCC.n7867 VSS 1.18e-19 
C11907 VCC.n7868 VSS 3.5e-20 
C11908 VCC.n7869 VSS 3.5e-20 
C11909 VCC.t216 VSS 1.55e-19 
C11910 VCC.n7870 VSS 7.57e-19 
C11911 VCC.n7871 VSS 4.73e-20 
C11912 VCC.n7872 VSS 1.54e-19 
C11913 VCC.n7873 VSS 2.88e-20 
C11914 VCC.n7874 VSS 2.88e-20 
C11915 VCC.n7875 VSS 3.5e-20 
C11916 VCC.n7876 VSS 5.76e-20 
C11917 VCC.n7877 VSS 9.88e-20 
C11918 VCC.n7878 VSS 1.3e-19 
C11919 VCC.n7879 VSS 3e-20 
C11920 VCC.t214 VSS 0.005f 
C11921 VCC.t278 VSS 0.00453f 
C11922 VCC.n7880 VSS 0.00229f 
C11923 VCC.n7881 VSS 1.91e-19 
C11924 VCC.n7882 VSS 3.5e-20 
C11925 VCC.n7883 VSS 3.14e-19 
C11926 VCC.n7884 VSS 3.5e-20 
C11927 VCC.n7885 VSS 2.47e-20 
C11928 VCC.n7886 VSS 5.76e-20 
C11929 VCC.n7887 VSS 2.47e-20 
C11930 VCC.n7888 VSS 8.23e-21 
C11931 VCC.n7889 VSS 2.88e-20 
C11932 VCC.n7890 VSS 5.76e-20 
C11933 VCC.n7891 VSS 2.47e-20 
C11934 VCC.n7892 VSS 2.88e-20 
C11935 VCC.n7893 VSS 2.47e-20 
C11936 VCC.n7894 VSS 5.15e-20 
C11937 VCC.n7895 VSS 4.73e-20 
C11938 VCC.n7896 VSS 3.7e-20 
C11939 VCC.n7897 VSS 3.5e-20 
C11940 VCC.n7898 VSS 7.41e-20 
C11941 VCC.t206 VSS 6.42e-19 
C11942 VCC.n7899 VSS 3e-20 
C11943 VCC.n7900 VSS 5.97e-20 
C11944 VCC.n7901 VSS 4.13e-19 
C11945 VCC.n7902 VSS 9.53e-20 
C11946 VCC.n7903 VSS 3.5e-20 
C11947 VCC.n7904 VSS 3.5e-20 
C11948 VCC.n7905 VSS 5.35e-20 
C11949 VCC.n7906 VSS 4.32e-20 
C11950 VCC.n7907 VSS 2.68e-20 
C11951 VCC.n7908 VSS 3.7e-20 
C11952 VCC.n7909 VSS 1.65e-20 
C11953 VCC.n7910 VSS 4.53e-20 
C11954 VCC.n7911 VSS 1.2e-19 
C11955 VCC.n7912 VSS 5.2e-19 
C11956 VCC.n7913 VSS 1.2e-19 
C11957 VCC.n7914 VSS 6.38e-20 
C11958 VCC.n7915 VSS 2.47e-20 
C11959 VCC.n7916 VSS 4.53e-20 
C11960 VCC.n7917 VSS 3.5e-20 
C11961 VCC.n7918 VSS 3.5e-20 
C11962 VCC.n7919 VSS 2.68e-20 
C11963 VCC.n7920 VSS 2.68e-20 
C11964 VCC.n7921 VSS 2.47e-20 
C11965 VCC.n7922 VSS 4.53e-20 
C11966 VCC.n7923 VSS 2.68e-20 
C11967 VCC.n7924 VSS 4.32e-20 
C11968 VCC.n7925 VSS 2.68e-20 
C11969 VCC.n7926 VSS 3.91e-20 
C11970 VCC.n7927 VSS 2.88e-20 
C11971 VCC.n7928 VSS 4.73e-20 
C11972 VCC.n7929 VSS 3.7e-20 
C11973 VCC.n7930 VSS 3.7e-20 
C11974 VCC.n7931 VSS 3.5e-20 
C11975 VCC.n7932 VSS 5.76e-20 
C11976 VCC.n7933 VSS 4.73e-20 
C11977 VCC.n7934 VSS 3.09e-20 
C11978 VCC.n7935 VSS 3.5e-20 
C11979 VCC.n7936 VSS 3.5e-20 
C11980 VCC.n7937 VSS 3.5e-20 
C11981 VCC.n7938 VSS 1.18e-19 
C11982 VCC.n7939 VSS 3e-20 
C11983 VCC.n7940 VSS 1.15e-19 
C11984 VCC.n7941 VSS 9.88e-20 
C11985 VCC.n7942 VSS 5.76e-20 
C11986 VCC.n7943 VSS 3.5e-20 
C11987 VCC.n7944 VSS 3.09e-20 
C11988 VCC.n7945 VSS 3.09e-20 
C11989 VCC.n7946 VSS 2.26e-20 
C11990 VCC.n7947 VSS 5.76e-20 
C11991 VCC.n7948 VSS 2.68e-20 
C11992 VCC.n7949 VSS 2.68e-20 
C11993 VCC.n7950 VSS 0.00185f 
C11994 VCC.n7951 VSS 2.72e-19 
C11995 VCC.n7952 VSS 2.26e-20 
C11996 VCC.n7953 VSS 1.87e-19 
C11997 VCC.n7954 VSS 3.5e-20 
C11998 VCC.n7955 VSS 2.68e-20 
C11999 VCC.n7956 VSS 5.97e-20 
C12000 VCC.n7957 VSS 4.73e-20 
C12001 VCC.n7958 VSS 4.73e-20 
C12002 VCC.n7959 VSS 5.15e-20 
C12003 VCC.n7960 VSS 7.41e-20 
C12004 VCC.n7961 VSS 3.7e-20 
C12005 VCC.n7962 VSS 2.26e-20 
C12006 VCC.n7963 VSS 6.38e-20 
C12007 VCC.n7964 VSS 4.73e-20 
C12008 VCC.n7965 VSS 3.29e-20 
C12009 VCC.n7966 VSS 3.5e-20 
C12010 VCC.n7967 VSS 3e-20 
C12011 VCC.t80 VSS 0.005f 
C12012 VCC.t174 VSS 0.00453f 
C12013 VCC.n7968 VSS 0.00228f 
C12014 VCC.n7969 VSS 1.3e-19 
C12015 VCC.t78 VSS 4.05e-19 
C12016 VCC.n7970 VSS 4.05e-19 
C12017 VCC.n7971 VSS 1.15e-19 
C12018 VCC.n7972 VSS 3.36e-19 
C12019 VCC.n7973 VSS 6.17e-21 
C12020 VCC.n7974 VSS 3.12e-19 
C12021 VCC.n7975 VSS 1.65e-20 
C12022 VCC.n7976 VSS 1.54e-19 
C12023 VCC.n7977 VSS 1.54e-19 
C12024 VCC.n7978 VSS 1.65e-20 
C12025 VCC.n7979 VSS 1.03e-20 
C12026 VCC.n7980 VSS 3.5e-20 
C12027 VCC.n7981 VSS 2.26e-20 
C12028 VCC.n7982 VSS 4.73e-20 
C12029 VCC.n7983 VSS 3.5e-20 
C12030 VCC.n7984 VSS 3e-20 
C12031 VCC.n7985 VSS 1.3e-19 
C12032 VCC.n7986 VSS 5.12e-19 
C12033 VCC.n7987 VSS 1.3e-19 
C12034 VCC.n7988 VSS 4.13e-19 
C12035 VCC.n7989 VSS 9.53e-20 
C12036 VCC.n7990 VSS 5.76e-20 
C12037 VCC.n7991 VSS 7.41e-20 
C12038 VCC.n7992 VSS 5.56e-20 
C12039 VCC.t79 VSS 1.55e-19 
C12040 VCC.n7993 VSS 3.91e-20 
C12041 VCC.n7994 VSS 3.91e-20 
C12042 VCC.n7995 VSS 1.85e-20 
C12043 VCC.n7996 VSS 7.55e-19 
C12044 VCC.n7997 VSS 4.94e-20 
C12045 VCC.n7998 VSS 5.15e-20 
C12046 VCC.n7999 VSS 7.2e-20 
C12047 VCC.n8000 VSS 1.38e-19 
C12048 VCC.n8001 VSS 1.17e-19 
C12049 VCC.n8002 VSS 4.32e-20 
C12050 VCC.n8003 VSS 2.88e-20 
C12051 VCC.n8004 VSS 2.68e-20 
C12052 VCC.n8005 VSS 3.5e-20 
C12053 VCC.n8006 VSS 3.5e-20 
C12054 VCC.n8007 VSS 2.88e-20 
C12055 VCC.n8008 VSS 2.68e-20 
C12056 VCC.n8009 VSS 2.68e-20 
C12057 VCC.n8010 VSS 2.68e-20 
C12058 VCC.n8011 VSS 4.12e-20 
C12059 VCC.n8012 VSS 4.12e-20 
C12060 VCC.n8013 VSS 3.91e-20 
C12061 VCC.n8014 VSS 4.53e-20 
C12062 VCC.n8015 VSS 4.53e-20 
C12063 VCC.n8016 VSS 1.05e-19 
C12064 VCC.n8017 VSS 1.05e-19 
C12065 VCC.n8018 VSS 4.32e-20 
C12066 VCC.n8019 VSS 3.7e-20 
C12067 VCC.n8020 VSS 2.68e-20 
C12068 VCC.n8021 VSS 2.68e-20 
C12069 VCC.n8022 VSS 6.79e-20 
C12070 VCC.n8023 VSS 9.26e-20 
C12071 VCC.n8024 VSS 1.83e-19 
C12072 VCC.n8025 VSS 7.95e-19 
C12073 VCC.n8026 VSS 5.2e-19 
C12074 VCC.n8027 VSS 1.3e-19 
C12075 VCC.n8028 VSS 3e-20 
C12076 VCC.n8029 VSS 3.5e-20 
C12077 VCC.n8030 VSS 5.97e-20 
C12078 VCC.n8031 VSS 7.41e-20 
C12079 VCC.n8032 VSS 5.15e-20 
C12080 VCC.n8033 VSS 5.15e-20 
C12081 VCC.n8034 VSS 3.09e-20 
C12082 VCC.n8035 VSS 3.09e-20 
C12083 VCC.n8036 VSS 3.7e-20 
C12084 VCC.n8037 VSS 2.68e-20 
C12085 VCC.n8038 VSS 3.91e-20 
C12086 VCC.n8039 VSS 1.17e-19 
C12087 VCC.n8040 VSS 1.38e-19 
C12088 VCC.n8041 VSS 7e-20 
C12089 VCC.n8042 VSS 4.73e-20 
C12090 VCC.n8043 VSS 3.5e-20 
C12091 VCC.n8044 VSS 3.5e-20 
C12092 VCC.n8045 VSS 3.5e-20 
C12093 VCC.n8046 VSS 4.53e-20 
C12094 VCC.n8047 VSS 1.18e-19 
C12095 VCC.n8048 VSS 5.12e-19 
C12096 VCC.n8049 VSS 1.3e-19 
C12097 VCC.n8050 VSS 1.61e-19 
C12098 VCC.n8051 VSS 9.9e-20 
C12099 VCC.n8052 VSS 0.00243f 
C12100 VCC.n8053 VSS 2.26e-20 
C12101 VCC.n8054 VSS 4.13e-19 
C12102 VCC.n8055 VSS 3.5e-20 
C12103 VCC.n8056 VSS 3.5e-20 
C12104 VCC.n8057 VSS 2.47e-20 
C12105 VCC.n8058 VSS 2.06e-20 
C12106 VCC.n8059 VSS 6.17e-20 
C12107 VCC.n8060 VSS 6.17e-20 
C12108 VCC.n8061 VSS 4.73e-20 
C12109 VCC.n8062 VSS 4.73e-20 
C12110 VCC.n8063 VSS 2.88e-20 
C12111 VCC.n8064 VSS 1.44e-20 
C12112 VCC.n8065 VSS 1.65e-20 
C12113 VCC.n8066 VSS 1.54e-19 
C12114 VCC.n8067 VSS 1.54e-19 
C12115 VCC.n8068 VSS 1.65e-20 
C12116 VCC.n8069 VSS 3.09e-20 
C12117 VCC.t207 VSS 1.55e-19 
C12118 VCC.n8070 VSS 0.00102f 
C12119 VCC.n8071 VSS 2.73e-19 
C12120 VCC.n8072 VSS 0.00136f 
C12121 VCC.n8073 VSS 2.73e-19 
C12122 VCC.n8074 VSS 0.00181f 
C12123 VCC.n8075 VSS 5.76e-20 
C12124 VCC.n8076 VSS 1.54e-19 
C12125 VCC.n8077 VSS 1.65e-20 
C12126 VCC.n8078 VSS 6.17e-20 
C12127 VCC.n8079 VSS 2.47e-20 
C12128 VCC.n8080 VSS 4.73e-20 
C12129 VCC.n8081 VSS 4.73e-20 
C12130 VCC.n8082 VSS 5.15e-20 
C12131 VCC.n8083 VSS 3.5e-20 
C12132 VCC.n8084 VSS 7.41e-20 
C12133 VCC.n8085 VSS 3.7e-20 
C12134 VCC.n8086 VSS 2.26e-20 
C12135 VCC.n8087 VSS 6.17e-20 
C12136 VCC.n8088 VSS 4.73e-20 
C12137 VCC.n8089 VSS 2.88e-20 
C12138 VCC.n8090 VSS 2.88e-20 
C12139 VCC.n8091 VSS 3.4e-19 
C12140 VCC.n8092 VSS 1.15e-19 
C12141 VCC.n8093 VSS 3.98e-19 
C12142 VCC.t215 VSS 4.05e-19 
C12143 VCC.n8094 VSS 1.22e-19 
C12144 VCC.n8095 VSS 1.3e-19 
C12145 VCC.n8096 VSS 3e-20 
C12146 VCC.n8097 VSS 3.5e-20 
C12147 VCC.n8098 VSS 3.5e-20 
C12148 VCC.n8099 VSS 4.73e-20 
C12149 VCC.n8100 VSS 2.47e-20 
C12150 VCC.n8101 VSS 1.23e-20 
C12151 VCC.n8102 VSS 1.65e-20 
C12152 VCC.n8103 VSS 2.47e-20 
C12153 VCC.n8104 VSS 5.76e-20 
C12154 VCC.n8105 VSS 1.38e-19 
C12155 VCC.n8106 VSS 7e-20 
C12156 VCC.n8107 VSS 3.7e-20 
C12157 VCC.n8108 VSS 2.47e-20 
C12158 VCC.n8109 VSS 3.7e-20 
C12159 VCC.n8110 VSS 1.85e-20 
C12160 VCC.n8111 VSS 3.09e-20 
C12161 VCC.n8112 VSS 5.35e-20 
C12162 VCC.n8113 VSS 4.73e-20 
C12163 VCC.n8114 VSS 5.35e-20 
C12164 VCC.n8115 VSS 7.41e-20 
C12165 VCC.n8116 VSS 5.76e-20 
C12166 VCC.n8117 VSS 9.53e-20 
C12167 VCC.n8118 VSS 4.13e-19 
C12168 VCC.n8119 VSS 1.3e-19 
C12169 VCC.n8120 VSS 5.2e-19 
C12170 VCC.n8121 VSS 1.2e-19 
C12171 VCC.n8122 VSS 4.73e-20 
C12172 VCC.n8123 VSS 2.68e-20 
C12173 VCC.n8124 VSS 3.5e-20 
C12174 VCC.n8125 VSS 3.5e-20 
C12175 VCC.n8126 VSS 2.68e-20 
C12176 VCC.n8127 VSS 2.68e-20 
C12177 VCC.n8128 VSS 4.32e-20 
C12178 VCC.n8129 VSS 4.32e-20 
C12179 VCC.n8130 VSS 4.32e-20 
C12180 VCC.n8131 VSS 2.88e-20 
C12181 VCC.n8132 VSS 3.5e-20 
C12182 VCC.n8133 VSS 2.68e-20 
C12183 VCC.n8134 VSS 7.82e-20 
C12184 VCC.n8135 VSS 4.73e-20 
C12185 VCC.n8136 VSS 4.73e-20 
C12186 VCC.n8137 VSS 1.05e-19 
C12187 VCC.n8138 VSS 1.05e-19 
C12188 VCC.n8139 VSS 4.53e-20 
C12189 VCC.n8140 VSS 2.68e-20 
C12190 VCC.n8141 VSS 2.68e-20 
C12191 VCC.n8142 VSS 6.59e-20 
C12192 VCC.n8143 VSS 9.26e-20 
C12193 VCC.n8144 VSS 6.59e-20 
C12194 VCC.n8145 VSS 2.47e-20 
C12195 VCC.n8146 VSS 2.47e-20 
C12196 VCC.n8147 VSS 2.88e-20 
C12197 VCC.n8148 VSS 3.5e-20 
C12198 VCC.n8149 VSS 3.5e-20 
C12199 VCC.n8150 VSS 4.53e-20 
C12200 VCC.n8151 VSS 1.2e-19 
C12201 VCC.n8152 VSS 5.2e-19 
C12202 VCC.n8153 VSS 1.3e-19 
C12203 VCC.n8154 VSS 4.13e-19 
C12204 VCC.n8155 VSS 9.53e-20 
C12205 VCC.n8156 VSS 5.97e-20 
C12206 VCC.n8157 VSS 7.41e-20 
C12207 VCC.n8158 VSS 5.35e-20 
C12208 VCC.n8159 VSS 5.15e-20 
C12209 VCC.n8160 VSS 3.09e-20 
C12210 VCC.n8161 VSS 3.09e-20 
C12211 VCC.n8162 VSS 3.91e-20 
C12212 VCC.n8163 VSS 2.47e-20 
C12213 VCC.n8164 VSS 3.7e-20 
C12214 VCC.n8165 VSS 1.17e-19 
C12215 VCC.n8166 VSS 1.38e-19 
C12216 VCC.n8167 VSS 7.2e-20 
C12217 VCC.n8168 VSS 4.73e-20 
C12218 VCC.n8169 VSS 3.5e-20 
C12219 VCC.n8170 VSS 3.5e-20 
C12220 VCC.n8171 VSS 4.53e-20 
C12221 VCC.n8172 VSS 5.97e-20 
C12222 VCC.n8173 VSS 3.5e-20 
C12223 VCC.n8174 VSS 3e-20 
C12224 VCC.n8175 VSS 1.3e-19 
C12225 VCC.n8176 VSS 1.53e-19 
C12226 VCC.t120 VSS 4.05e-19 
C12227 VCC.n8177 VSS 1.35e-19 
C12228 VCC.t218 VSS 4.21e-19 
C12229 VCC.n8178 VSS 2.06e-19 
C12230 VCC.n8179 VSS 1.32e-19 
C12231 VCC.n8180 VSS 9.67e-20 
C12232 VCC.n8181 VSS 3.35e-20 
C12233 VCC.n8182 VSS 3.5e-20 
C12234 VCC.n8183 VSS 2.36e-19 
C12235 VCC.n8184 VSS 0.0023f 
C12236 VCC.t217 VSS 0.0031f 
C12237 VCC.t296 VSS 0.00366f 
C12238 VCC.t220 VSS 0.00365f 
C12239 VCC.t297 VSS 0.00386f 
C12240 VCC.n8185 VSS 0.00569f 
C12241 VCC.n8186 VSS 1.3e-19 
C12242 VCC.n8187 VSS 3.67e-19 
C12243 VCC.n8188 VSS 1.15e-19 
C12244 VCC.n8189 VSS 3.38e-19 
C12245 VCC.n8190 VSS 3.5e-20 
C12246 VCC.n8191 VSS 3.5e-20 
C12247 VCC.n8192 VSS 2.68e-20 
C12248 VCC.n8193 VSS 2.06e-20 
C12249 VCC.n8194 VSS 6.38e-20 
C12250 VCC.n8195 VSS 5.97e-20 
C12251 VCC.n8196 VSS 4.73e-20 
C12252 VCC.n8197 VSS 4.73e-20 
C12253 VCC.n8198 VSS 3.09e-20 
C12254 VCC.n8199 VSS 1.23e-20 
C12255 VCC.n8200 VSS 1.65e-20 
C12256 VCC.n8201 VSS 1.54e-19 
C12257 VCC.n8202 VSS 1.54e-19 
C12258 VCC.n8203 VSS 1.65e-20 
C12259 VCC.n8204 VSS 3.29e-20 
C12260 VCC.t121 VSS 1.67e-19 
C12261 VCC.n8205 VSS 0.00101f 
C12262 VCC.n8206 VSS 2.71e-19 
C12263 VCC.n8207 VSS 7.46e-19 
C12264 VCC.n8208 VSS 0.00333f 
C12265 VCC.n8209 VSS 2.46e-19 
C12266 VCC.n8210 VSS 3.02e-19 
C12267 VCC.n8211 VSS 3.7e-20 
C12268 VCC.n8212 VSS 5.15e-20 
C12269 VCC.n8213 VSS 5.97e-20 
C12270 VCC.n8214 VSS 6.38e-20 
C12271 VCC.n8215 VSS 4.73e-20 
C12272 VCC.n8216 VSS 4.73e-20 
C12273 VCC.n8217 VSS 2.68e-20 
C12274 VCC.n8218 VSS 3.29e-20 
C12275 VCC.n8219 VSS 1.65e-20 
C12276 VCC.n8220 VSS 1.54e-19 
C12277 VCC.n8221 VSS 1.54e-19 
C12278 VCC.n8222 VSS 1.65e-20 
C12279 VCC.n8223 VSS 3.09e-20 
C12280 VCC.n8224 VSS 3.09e-20 
C12281 VCC.n8225 VSS 4.73e-20 
C12282 VCC.n8226 VSS 4.32e-20 
C12283 VCC.n8227 VSS 3.5e-20 
C12284 VCC.n8228 VSS 3.5e-20 
C12285 VCC.n8229 VSS 1.35e-19 
C12286 VCC.n8230 VSS 5.24e-19 
C12287 VCC.n8231 VSS 1.4e-19 
C12288 VCC.n8232 VSS 5.4e-19 
C12289 VCC.n8233 VSS 1.35e-19 
C12290 VCC.n8234 VSS 4.37e-19 
C12291 VCC.n8235 VSS 1.13e-19 
C12292 VCC.n8236 VSS 8.23e-21 
C12293 VCC.n8237 VSS 1.65e-20 
C12294 VCC.n8238 VSS 3.5e-20 
C12295 VCC.n8239 VSS 3.91e-20 
C12296 VCC.n8240 VSS 3.09e-20 
C12297 VCC.n8241 VSS 1.85e-20 
C12298 VCC.n8242 VSS 3.5e-20 
C12299 VCC.n8243 VSS 1.05e-19 
C12300 VCC.n8244 VSS 2.06e-20 
C12301 VCC.n8245 VSS 2.26e-20 
C12302 VCC.n8246 VSS 3.7e-20 
C12303 VCC.n8247 VSS 5.15e-20 
C12304 VCC.n8248 VSS 1.38e-19 
C12305 VCC.n8249 VSS 1.17e-19 
C12306 VCC.n8250 VSS 4.32e-20 
C12307 VCC.n8251 VSS 2.88e-20 
C12308 VCC.n8252 VSS 2.68e-20 
C12309 VCC.n8253 VSS 6.59e-20 
C12310 VCC.n8254 VSS 5.56e-20 
C12311 VCC.n8255 VSS 2.68e-20 
C12312 VCC.n8256 VSS 4.32e-20 
C12313 VCC.n8257 VSS 1.05e-19 
C12314 VCC.n8258 VSS 3.09e-20 
C12315 VCC.n8259 VSS 3.7e-20 
C12316 VCC.n8260 VSS 4.32e-20 
C12317 VCC.n8261 VSS 1.05e-19 
C12318 VCC.n8262 VSS 4.53e-20 
C12319 VCC.n8263 VSS 4.53e-20 
C12320 VCC.n8264 VSS 7.82e-20 
C12321 VCC.n8265 VSS 2.18e-19 
C12322 VCC.n8266 VSS 1.4e-19 
C12323 VCC.n8267 VSS 1.4e-19 
C12324 VCC.n8268 VSS 5.4e-19 
C12325 VCC.n8269 VSS 1.35e-19 
C12326 VCC.t39 VSS 4.21e-19 
C12327 VCC.n8270 VSS 3.33e-19 
C12328 VCC.n8271 VSS 1.13e-19 
C12329 VCC.n8272 VSS 8.23e-21 
C12330 VCC.n8273 VSS 1.65e-20 
C12331 VCC.n8274 VSS 3.5e-20 
C12332 VCC.n8275 VSS 3.5e-20 
C12333 VCC.n8276 VSS 3.5e-20 
C12334 VCC.n8277 VSS 1.17e-19 
C12335 VCC.n8278 VSS 1.38e-19 
C12336 VCC.n8279 VSS 5.15e-20 
C12337 VCC.n8280 VSS 4.73e-20 
C12338 VCC.n8281 VSS 7.2e-20 
C12339 VCC.n8282 VSS 2.68e-20 
C12340 VCC.n8283 VSS 1.65e-20 
C12341 VCC.n8284 VSS 1.54e-19 
C12342 VCC.n8285 VSS 1.54e-19 
C12343 VCC.n8286 VSS 1.65e-20 
C12344 VCC.n8287 VSS 2.47e-20 
C12345 VCC.n8288 VSS 1.23e-20 
C12346 VCC.n8289 VSS 7.62e-19 
C12347 VCC.n8290 VSS 4.12e-20 
C12348 VCC.n8291 VSS 5.15e-20 
C12349 VCC.n8292 VSS 6.59e-20 
C12350 VCC.n8293 VSS 5.76e-20 
C12351 VCC.n8294 VSS 4.73e-20 
C12352 VCC.n8295 VSS 2.26e-20 
C12353 VCC.n8296 VSS 2.68e-20 
C12354 VCC.n8297 VSS 1.03e-20 
C12355 VCC.n8298 VSS 3.5e-20 
C12356 VCC.n8299 VSS 3.5e-20 
C12357 VCC.n8300 VSS 1.35e-19 
C12358 VCC.n8301 VSS 4.53e-19 
C12359 VCC.n8302 VSS 7.71e-19 
C12360 VCC.n8303 VSS 1.32e-19 
C12361 VCC.n8304 VSS 3.5e-20 
C12362 VCC.n8305 VSS 3.42e-20 
C12363 VCC.n8306 VSS 2.36e-19 
C12364 VCC.n8307 VSS 3.21e-19 
C12365 VCC.n8308 VSS 2.61e-19 
C12366 VCC.n8309 VSS 0.00189f 
C12367 VCC.n8310 VSS 2.68e-19 
C12368 VCC.n8311 VSS 5.76e-20 
C12369 VCC.n8312 VSS 2.88e-20 
C12370 VCC.n8313 VSS 3.5e-20 
C12371 VCC.n8314 VSS 3.42e-20 
C12372 VCC.n8315 VSS 3.5e-20 
C12373 VCC.n8316 VSS 4.53e-19 
C12374 VCC.n8317 VSS 1.17e-19 
C12375 VCC.n8318 VSS 3.5e-20 
C12376 VCC.n8319 VSS 1.44e-20 
C12377 VCC.n8320 VSS 4.12e-20 
C12378 VCC.n8321 VSS 5.76e-20 
C12379 VCC.n8322 VSS 5.76e-20 
C12380 VCC.n8323 VSS 2.06e-20 
C12381 VCC.n8324 VSS 3.29e-20 
C12382 VCC.n8325 VSS 7.2e-20 
C12383 VCC.n8326 VSS 3.29e-20 
C12384 VCC.n8327 VSS 4.73e-20 
C12385 VCC.n8328 VSS 2.26e-20 
C12386 VCC.n8329 VSS 1.01e-19 
C12387 VCC.n8330 VSS 1.36e-19 
C12388 VCC.n8331 VSS 1.35e-19 
C12389 VCC.n8332 VSS 3.5e-20 
C12390 VCC.n8333 VSS 3.5e-20 
C12391 VCC.n8334 VSS 3.5e-20 
C12392 VCC.n8335 VSS 3.5e-20 
C12393 VCC.n8336 VSS 3.09e-20 
C12394 VCC.n8337 VSS 3.91e-20 
C12395 VCC.n8338 VSS 4.73e-20 
C12396 VCC.n8339 VSS 4.32e-20 
C12397 VCC.n8340 VSS 2.68e-20 
C12398 VCC.n8341 VSS 4.53e-20 
C12399 VCC.n8342 VSS 4.53e-20 
C12400 VCC.n8343 VSS 3.09e-20 
C12401 VCC.n8344 VSS 4.32e-20 
C12402 VCC.n8345 VSS 2.68e-20 
C12403 VCC.n8346 VSS 7.82e-20 
C12404 VCC.n8347 VSS 5.56e-20 
C12405 VCC.n8348 VSS 1.4e-19 
C12406 VCC.n8349 VSS 2.18e-19 
C12407 VCC.n8350 VSS 1.35e-19 
C12408 VCC.n8351 VSS 1.13e-19 
C12409 VCC.n8352 VSS 3.5e-20 
C12410 VCC.n8353 VSS 1.85e-20 
C12411 VCC.n8354 VSS 3.7e-20 
C12412 VCC.n8355 VSS 3.09e-20 
C12413 VCC.n8356 VSS 6.59e-20 
C12414 VCC.n8357 VSS 2.68e-20 
C12415 VCC.n8358 VSS 5.76e-20 
C12416 VCC.n8359 VSS 4.73e-20 
C12417 VCC.n8360 VSS 3.5e-20 
C12418 VCC.t66 VSS 1.56e-19 
C12419 VCC.n8361 VSS 7.97e-19 
C12420 VCC.n8362 VSS 3.09e-20 
C12421 VCC.n8363 VSS 3.5e-20 
C12422 VCC.n8364 VSS 3.5e-20 
C12423 VCC.t65 VSS 4.21e-19 
C12424 VCC.n8365 VSS 1.32e-19 
C12425 VCC.n8366 VSS 1.09e-19 
C12426 VCC.n8367 VSS 3.5e-20 
C12427 VCC.n8368 VSS 3.09e-20 
C12428 VCC.n8369 VSS 5.97e-20 
C12429 VCC.n8370 VSS 2.26e-20 
C12430 VCC.n8371 VSS 5.76e-20 
C12431 VCC.n8372 VSS 2.68e-20 
C12432 VCC.n8373 VSS 2.68e-20 
C12433 VCC.n8374 VSS 1.9e-19 
C12434 VCC.n8375 VSS 5.76e-20 
C12435 VCC.n8376 VSS 2.68e-20 
C12436 VCC.n8377 VSS 2.68e-20 
C12437 VCC.n8378 VSS 2.68e-20 
C12438 VCC.n8379 VSS 5.76e-20 
C12439 VCC.n8380 VSS 2.26e-20 
C12440 VCC.n8381 VSS 3.09e-20 
C12441 VCC.n8382 VSS 2.26e-20 
C12442 VCC.n8383 VSS 5.15e-20 
C12443 VCC.n8384 VSS 4.73e-20 
C12444 VCC.n8385 VSS 3.7e-20 
C12445 VCC.n8386 VSS 3.5e-20 
C12446 VCC.n8387 VSS 7.41e-20 
C12447 VCC.n8388 VSS 1.91e-19 
C12448 VCC.n8389 VSS 9.88e-20 
C12449 VCC.n8390 VSS 3e-20 
C12450 VCC.n8391 VSS 5.12e-19 
C12451 VCC.n8392 VSS 1.18e-19 
C12452 VCC.n8393 VSS 3.5e-20 
C12453 VCC.n8394 VSS 3.5e-20 
C12454 VCC.n8395 VSS 5.15e-20 
C12455 VCC.n8396 VSS 4.32e-20 
C12456 VCC.n8397 VSS 2.68e-20 
C12457 VCC.n8398 VSS 3.91e-20 
C12458 VCC.n8399 VSS 1.44e-20 
C12459 VCC.n8400 VSS 3.5e-20 
C12460 VCC.n8401 VSS 3e-20 
C12461 VCC.n8402 VSS 7.95e-19 
C12462 VCC.n8403 VSS 1.83e-19 
C12463 VCC.n8404 VSS 2.88e-20 
C12464 VCC.n8405 VSS 2.68e-20 
C12465 VCC.n8406 VSS 2.68e-20 
C12466 VCC.n8407 VSS 2.68e-20 
C12467 VCC.n8408 VSS 4.53e-20 
C12468 VCC.n8409 VSS 3.7e-20 
C12469 VCC.n8410 VSS 7.82e-20 
C12470 VCC.n8411 VSS 1.17e-19 
C12471 VCC.n8412 VSS 3.91e-20 
C12472 VCC.n8413 VSS 1.65e-20 
C12473 VCC.n8414 VSS 2.68e-20 
C12474 VCC.n8415 VSS 3.5e-20 
C12475 VCC.n8416 VSS 3e-20 
C12476 VCC.n8417 VSS 5.12e-19 
C12477 VCC.n8418 VSS 1.18e-19 
C12478 VCC.n8419 VSS 3.5e-20 
C12479 VCC.n8420 VSS 3.5e-20 
C12480 VCC.t153 VSS 1.55e-19 
C12481 VCC.n8421 VSS 7.57e-19 
C12482 VCC.n8422 VSS 4.73e-20 
C12483 VCC.n8423 VSS 1.54e-19 
C12484 VCC.n8424 VSS 2.88e-20 
C12485 VCC.n8425 VSS 2.88e-20 
C12486 VCC.n8426 VSS 3.5e-20 
C12487 VCC.n8427 VSS 5.76e-20 
C12488 VCC.n8428 VSS 9.88e-20 
C12489 VCC.n8429 VSS 1.3e-19 
C12490 VCC.n8430 VSS 3e-20 
C12491 VCC.t154 VSS 0.005f 
C12492 VCC.t55 VSS 0.00453f 
C12493 VCC.n8431 VSS 0.00229f 
C12494 VCC.n8432 VSS 1.91e-19 
C12495 VCC.n8433 VSS 3.5e-20 
C12496 VCC.n8434 VSS 3.14e-19 
C12497 VCC.n8435 VSS 2.47e-20 
C12498 VCC.n8436 VSS 2.73e-19 
C12499 VCC.n8437 VSS 0.00185f 
C12500 VCC.n8438 VSS 5.76e-20 
C12501 VCC.n8439 VSS 1.54e-19 
C12502 VCC.n8440 VSS 1.65e-20 
C12503 VCC.n8441 VSS 2.88e-20 
C12504 VCC.n8442 VSS 2.47e-20 
C12505 VCC.n8443 VSS 6.17e-20 
C12506 VCC.n8444 VSS 4.73e-20 
C12507 VCC.n8445 VSS 4.73e-20 
C12508 VCC.n8446 VSS 5.15e-20 
C12509 VCC.n8447 VSS 3.5e-20 
C12510 VCC.n8448 VSS 7.41e-20 
C12511 VCC.n8449 VSS 3.7e-20 
C12512 VCC.n8450 VSS 2.26e-20 
C12513 VCC.n8451 VSS 6.17e-20 
C12514 VCC.n8452 VSS 4.73e-20 
C12515 VCC.n8453 VSS 3.5e-20 
C12516 VCC.n8454 VSS 2.88e-20 
C12517 VCC.n8455 VSS 3.4e-19 
C12518 VCC.n8456 VSS 1.15e-19 
C12519 VCC.n8457 VSS 3.98e-19 
C12520 VCC.t152 VSS 4.05e-19 
C12521 VCC.n8458 VSS 1.22e-19 
C12522 VCC.n8459 VSS 1.3e-19 
C12523 VCC.n8460 VSS 3e-20 
C12524 VCC.n8461 VSS 3.5e-20 
C12525 VCC.n8462 VSS 3.5e-20 
C12526 VCC.n8463 VSS 4.73e-20 
C12527 VCC.n8464 VSS 2.47e-20 
C12528 VCC.n8465 VSS 1.23e-20 
C12529 VCC.n8466 VSS 1.65e-20 
C12530 VCC.n8467 VSS 2.47e-20 
C12531 VCC.n8468 VSS 5.76e-20 
C12532 VCC.n8469 VSS 1.38e-19 
C12533 VCC.n8470 VSS 7e-20 
C12534 VCC.n8471 VSS 3.7e-20 
C12535 VCC.n8472 VSS 2.47e-20 
C12536 VCC.n8473 VSS 3.7e-20 
C12537 VCC.n8474 VSS 1.85e-20 
C12538 VCC.n8475 VSS 3.09e-20 
C12539 VCC.n8476 VSS 5.35e-20 
C12540 VCC.n8477 VSS 4.73e-20 
C12541 VCC.n8478 VSS 5.35e-20 
C12542 VCC.n8479 VSS 7.41e-20 
C12543 VCC.n8480 VSS 5.76e-20 
C12544 VCC.n8481 VSS 9.53e-20 
C12545 VCC.n8482 VSS 4.13e-19 
C12546 VCC.n8483 VSS 1.3e-19 
C12547 VCC.n8484 VSS 5.2e-19 
C12548 VCC.n8485 VSS 1.2e-19 
C12549 VCC.n8486 VSS 4.73e-20 
C12550 VCC.n8487 VSS 2.68e-20 
C12551 VCC.n8488 VSS 3.5e-20 
C12552 VCC.n8489 VSS 3.5e-20 
C12553 VCC.n8490 VSS 2.68e-20 
C12554 VCC.n8491 VSS 2.68e-20 
C12555 VCC.n8492 VSS 4.32e-20 
C12556 VCC.n8493 VSS 4.32e-20 
C12557 VCC.n8494 VSS 4.32e-20 
C12558 VCC.n8495 VSS 2.88e-20 
C12559 VCC.n8496 VSS 3.5e-20 
C12560 VCC.n8497 VSS 2.68e-20 
C12561 VCC.n8498 VSS 7.82e-20 
C12562 VCC.n8499 VSS 4.73e-20 
C12563 VCC.n8500 VSS 4.73e-20 
C12564 VCC.n8501 VSS 1.05e-19 
C12565 VCC.n8502 VSS 1.05e-19 
C12566 VCC.n8503 VSS 4.53e-20 
C12567 VCC.n8504 VSS 2.68e-20 
C12568 VCC.n8505 VSS 2.68e-20 
C12569 VCC.n8506 VSS 6.59e-20 
C12570 VCC.n8507 VSS 9.26e-20 
C12571 VCC.n8508 VSS 6.59e-20 
C12572 VCC.n8509 VSS 2.47e-20 
C12573 VCC.n8510 VSS 2.47e-20 
C12574 VCC.n8511 VSS 2.88e-20 
C12575 VCC.n8512 VSS 3.5e-20 
C12576 VCC.n8513 VSS 3.5e-20 
C12577 VCC.n8514 VSS 4.53e-20 
C12578 VCC.n8515 VSS 1.2e-19 
C12579 VCC.n8516 VSS 5.2e-19 
C12580 VCC.n8517 VSS 1.3e-19 
C12581 VCC.n8518 VSS 4.13e-19 
C12582 VCC.n8519 VSS 9.53e-20 
C12583 VCC.n8520 VSS 5.97e-20 
C12584 VCC.n8521 VSS 7.41e-20 
C12585 VCC.n8522 VSS 5.35e-20 
C12586 VCC.n8523 VSS 5.15e-20 
C12587 VCC.n8524 VSS 3.09e-20 
C12588 VCC.n8525 VSS 3.09e-20 
C12589 VCC.n8526 VSS 3.91e-20 
C12590 VCC.n8527 VSS 2.47e-20 
C12591 VCC.n8528 VSS 3.7e-20 
C12592 VCC.n8529 VSS 1.17e-19 
C12593 VCC.n8530 VSS 1.38e-19 
C12594 VCC.n8531 VSS 7.2e-20 
C12595 VCC.n8532 VSS 4.73e-20 
C12596 VCC.n8533 VSS 3.5e-20 
C12597 VCC.n8534 VSS 3.5e-20 
C12598 VCC.n8535 VSS 4.53e-20 
C12599 VCC.n8536 VSS 5.97e-20 
C12600 VCC.n8537 VSS 3.5e-20 
C12601 VCC.n8538 VSS 3e-20 
C12602 VCC.n8539 VSS 1.3e-19 
C12603 VCC.n8540 VSS 1.53e-19 
C12604 VCC.t276 VSS 4.05e-19 
C12605 VCC.n8541 VSS 2.06e-19 
C12606 VCC.n8542 VSS 1.35e-19 
C12607 VCC.n8543 VSS 9.67e-20 
C12608 VCC.n8544 VSS 3.35e-20 
C12609 VCC.n8545 VSS 3.5e-20 
C12610 VCC.n8546 VSS 2.36e-19 
C12611 VCC.n8547 VSS 0.0023f 
C12612 VCC.t68 VSS 0.0031f 
C12613 VCC.t128 VSS 0.00366f 
C12614 VCC.t67 VSS 0.00365f 
C12615 VCC.t129 VSS 0.00386f 
C12616 VCC.n8548 VSS 0.00569f 
C12617 VCC.n8549 VSS 1.3e-19 
C12618 VCC.n8550 VSS 3.67e-19 
C12619 VCC.n8551 VSS 1.15e-19 
C12620 VCC.n8552 VSS 3.38e-19 
C12621 VCC.n8553 VSS 3.5e-20 
C12622 VCC.n8554 VSS 3.5e-20 
C12623 VCC.n8555 VSS 2.68e-20 
C12624 VCC.n8556 VSS 2.06e-20 
C12625 VCC.n8557 VSS 6.38e-20 
C12626 VCC.n8558 VSS 5.97e-20 
C12627 VCC.n8559 VSS 4.73e-20 
C12628 VCC.n8560 VSS 4.73e-20 
C12629 VCC.n8561 VSS 3.09e-20 
C12630 VCC.n8562 VSS 1.23e-20 
C12631 VCC.n8563 VSS 1.65e-20 
C12632 VCC.n8564 VSS 1.54e-19 
C12633 VCC.n8565 VSS 1.54e-19 
C12634 VCC.n8566 VSS 1.65e-20 
C12635 VCC.n8567 VSS 3.29e-20 
C12636 VCC.t277 VSS 1.67e-19 
C12637 VCC.n8568 VSS 0.00101f 
C12638 VCC.n8569 VSS 2.71e-19 
C12639 VCC.n8570 VSS 7.46e-19 
C12640 VCC.n8571 VSS 0.00333f 
C12641 VCC.n8572 VSS 2.46e-19 
C12642 VCC.n8573 VSS 3.02e-19 
C12643 VCC.n8574 VSS 3.7e-20 
C12644 VCC.n8575 VSS 5.15e-20 
C12645 VCC.n8576 VSS 6.38e-20 
C12646 VCC.n8577 VSS 4.73e-20 
C12647 VCC.n8578 VSS 4.73e-20 
C12648 VCC.n8579 VSS 2.68e-20 
C12649 VCC.n8580 VSS 3.29e-20 
C12650 VCC.n8581 VSS 1.65e-20 
C12651 VCC.n8582 VSS 1.54e-19 
C12652 VCC.n8583 VSS 1.54e-19 
C12653 VCC.n8584 VSS 5.56e-20 
C12654 VCC.n8585 VSS 2.88e-20 
C12655 VCC.n8586 VSS 1.65e-20 
C12656 VCC.n8587 VSS 3.09e-20 
C12657 VCC.n8588 VSS 4.73e-20 
C12658 VCC.n8589 VSS 4.73e-20 
C12659 VCC.n8590 VSS 4.32e-20 
C12660 VCC.n8591 VSS 1.17e-19 
C12661 VCC.n8592 VSS 3.33e-19 
C12662 VCC.n8593 VSS 1.35e-19 
C12663 VCC.n8594 VSS 4.37e-19 
C12664 VCC.n8595 VSS 5.24e-19 
C12665 VCC.n8596 VSS 1.36e-19 
C12666 VCC.n8597 VSS 1.01e-19 
C12667 VCC.n8598 VSS 1.05e-19 
C12668 VCC.n8599 VSS 2.06e-20 
C12669 VCC.n8600 VSS 2.26e-20 
C12670 VCC.n8601 VSS 3.7e-20 
C12671 VCC.n8602 VSS 5.15e-20 
C12672 VCC.n8603 VSS 1.38e-19 
C12673 VCC.n8604 VSS 3.91e-20 
C12674 VCC.n8605 VSS 2.88e-20 
C12675 VCC.n8606 VSS 4.32e-20 
C12676 VCC.n8607 VSS 1.17e-19 
C12677 VCC.n8608 VSS 3.7e-20 
C12678 VCC.n8609 VSS 3.91e-20 
C12679 VCC.n8610 VSS 3.5e-20 
C12680 VCC.n8611 VSS 1.65e-20 
C12681 VCC.n8612 VSS 8.23e-21 
C12682 VCC.n8613 VSS 3.5e-20 
C12683 VCC.n8614 VSS 3.5e-20 
C12684 VCC.n8615 VSS 1.4e-19 
C12685 VCC.n8616 VSS 5.4e-19 
C12686 VCC.n8617 VSS 8.42e-19 
C12687 VCC.n8618 VSS 5.4e-19 
C12688 VCC.n8619 VSS 1.4e-19 
C12689 VCC.n8620 VSS 1.4e-19 
C12690 VCC.n8621 VSS 2.18e-19 
C12691 VCC.n8622 VSS 7.82e-20 
C12692 VCC.n8623 VSS 4.32e-20 
C12693 VCC.n8624 VSS 4.32e-20 
C12694 VCC.n8625 VSS 1.05e-19 
C12695 VCC.n8626 VSS 1.05e-19 
C12696 VCC.n8627 VSS 4.32e-20 
C12697 VCC.n8628 VSS 3.7e-20 
C12698 VCC.n8629 VSS 2.68e-20 
C12699 VCC.n8630 VSS 5.76e-20 
C12700 VCC.n8631 VSS 6.38e-20 
C12701 VCC.n8632 VSS 3.5e-20 
C12702 VCC.n8633 VSS 3.5e-20 
C12703 VCC.n8634 VSS 1.17e-19 
C12704 VCC.n8635 VSS 1.38e-19 
C12705 VCC.n8636 VSS 5.15e-20 
C12706 VCC.n8637 VSS 1.05e-19 
C12707 VCC.n8638 VSS 2.26e-20 
C12708 VCC.n8639 VSS 5.76e-20 
C12709 VCC.n8640 VSS 3.7e-20 
C12710 VCC.n8641 VSS 3.7e-20 
C12711 VCC.n8642 VSS 3.09e-20 
C12712 VCC.n8643 VSS 1.85e-20 
C12713 VCC.n8644 VSS 1.65e-20 
C12714 VCC.n8645 VSS 8.23e-21 
C12715 VCC.n8646 VSS 1.13e-19 
C12716 VCC.n8647 VSS 3.33e-19 
C12717 VCC.t294 VSS 4.21e-19 
C12718 VCC.n8648 VSS 2.06e-19 
C12719 VCC.n8649 VSS 1.35e-19 
C12720 VCC.n8650 VSS 3.5e-20 
C12721 VCC.n8651 VSS 3.5e-20 
C12722 VCC.n8652 VSS 3.5e-20 
C12723 VCC.n8653 VSS 1.03e-20 
C12724 VCC.n8654 VSS 2.68e-20 
C12725 VCC.n8655 VSS 3.09e-20 
C12726 VCC.n8656 VSS 2.68e-20 
C12727 VCC.n8657 VSS 1.65e-20 
C12728 VCC.n8658 VSS 1.54e-19 
C12729 VCC.n8659 VSS 1.54e-19 
C12730 VCC.n8660 VSS 1.65e-20 
C12731 VCC.t295 VSS 1.56e-19 
C12732 VCC.n8661 VSS 7.62e-19 
C12733 VCC.n8662 VSS 1.23e-20 
C12734 VCC.n8663 VSS 2.47e-20 
C12735 VCC.n8664 VSS 4.73e-20 
C12736 VCC.n8665 VSS 6.59e-20 
C12737 VCC.n8666 VSS 5.15e-20 
C12738 VCC.n8667 VSS 2.47e-20 
C12739 VCC.n8668 VSS 7.41e-20 
C12740 VCC.n8669 VSS 9.47e-20 
C12741 VCC.n8670 VSS 1.32e-19 
C12742 VCC.n8671 VSS 7.71e-19 
C12743 VCC.n8672 VSS 9.83e-19 
C12744 VCC.n8673 VSS 2.36e-19 
C12745 VCC.n8674 VSS 3.21e-19 
C12746 VCC.n8675 VSS 2.61e-19 
C12747 VCC.n8676 VSS 0.00189f 
C12748 VCC.n8677 VSS 0.00247f 
C12749 VCC.n8678 VSS 0.00274f 
C12750 VCC.n8679 VSS 3.52e-19 
C12751 VCC.n8680 VSS 0.00276f 
C12752 VCC.n8681 VSS 0.00246f 
C12753 VCC.n8682 VSS 0.00274f 
.ends

X1 D0 VREFL D1 D2 D3 D4 D5 D0_BUF VREFH D1_BUF D2_BUF D3_BUF D4_BUF
+ D5_BUF VOUT VCC VSS x6_bit_dac


.param mc_mm_switch=0
.param mc_pr_switch=0
.lib "/foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice.tt.red" tt

V1 VSS 0 dc 0
V2 VCC 0 dc 3.3

V3 VREFL 0 dc 0
V4 VREFH 0 dc 3.3

V5  D0 0 PULSE(0 1.8 4n 1p 1p 4n 8n)
V6  D1 0 PULSE(0 1.8 8n 1p 1p 8n 16n)
V7  D2 0 PULSE(0 1.8 16n 1p 1p 16n 32n)
V8  D3 0 PULSE(0 1.8 32n 1p 1p 32n 64n)
V9  D4 0 PULSE(0 1.8 64n 1p 1p 64n 128n)
V10 D5 0 PULSE(0 1.8 128n 1p 1p 128n 256n)

.tran 1n 256n uic


.control
run

set xbrushwidth=3
set hcopydevtype = svg

plot D3 D4 D5 VOUT

hardcopy 4_bit_dac_RCX.svg D0 D1 D2 D3 VOUT

.endc
.end
